// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 3 2025 14:09:01

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    rgb_g,
    T01,
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    clock_output,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T45,
    T12,
    s4_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output rgb_g;
    output T01;
    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output clock_output;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T45;
    output T12;
    output s4_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__50564;
    wire N__50563;
    wire N__50562;
    wire N__50553;
    wire N__50552;
    wire N__50551;
    wire N__50544;
    wire N__50543;
    wire N__50542;
    wire N__50535;
    wire N__50534;
    wire N__50533;
    wire N__50526;
    wire N__50525;
    wire N__50524;
    wire N__50517;
    wire N__50516;
    wire N__50515;
    wire N__50508;
    wire N__50507;
    wire N__50506;
    wire N__50499;
    wire N__50498;
    wire N__50497;
    wire N__50490;
    wire N__50489;
    wire N__50488;
    wire N__50481;
    wire N__50480;
    wire N__50479;
    wire N__50472;
    wire N__50471;
    wire N__50470;
    wire N__50463;
    wire N__50462;
    wire N__50461;
    wire N__50454;
    wire N__50453;
    wire N__50452;
    wire N__50445;
    wire N__50444;
    wire N__50443;
    wire N__50436;
    wire N__50435;
    wire N__50434;
    wire N__50427;
    wire N__50426;
    wire N__50425;
    wire N__50418;
    wire N__50417;
    wire N__50416;
    wire N__50409;
    wire N__50408;
    wire N__50407;
    wire N__50390;
    wire N__50387;
    wire N__50386;
    wire N__50385;
    wire N__50382;
    wire N__50379;
    wire N__50376;
    wire N__50371;
    wire N__50366;
    wire N__50363;
    wire N__50362;
    wire N__50359;
    wire N__50356;
    wire N__50355;
    wire N__50354;
    wire N__50349;
    wire N__50346;
    wire N__50343;
    wire N__50338;
    wire N__50335;
    wire N__50332;
    wire N__50329;
    wire N__50324;
    wire N__50321;
    wire N__50320;
    wire N__50319;
    wire N__50318;
    wire N__50317;
    wire N__50316;
    wire N__50315;
    wire N__50314;
    wire N__50313;
    wire N__50312;
    wire N__50311;
    wire N__50310;
    wire N__50309;
    wire N__50308;
    wire N__50307;
    wire N__50306;
    wire N__50305;
    wire N__50304;
    wire N__50303;
    wire N__50302;
    wire N__50301;
    wire N__50300;
    wire N__50299;
    wire N__50298;
    wire N__50297;
    wire N__50296;
    wire N__50295;
    wire N__50294;
    wire N__50293;
    wire N__50292;
    wire N__50291;
    wire N__50290;
    wire N__50289;
    wire N__50288;
    wire N__50287;
    wire N__50286;
    wire N__50285;
    wire N__50284;
    wire N__50283;
    wire N__50282;
    wire N__50281;
    wire N__50280;
    wire N__50279;
    wire N__50278;
    wire N__50277;
    wire N__50276;
    wire N__50275;
    wire N__50274;
    wire N__50273;
    wire N__50272;
    wire N__50271;
    wire N__50270;
    wire N__50269;
    wire N__50268;
    wire N__50267;
    wire N__50266;
    wire N__50265;
    wire N__50264;
    wire N__50263;
    wire N__50262;
    wire N__50261;
    wire N__50260;
    wire N__50259;
    wire N__50258;
    wire N__50257;
    wire N__50256;
    wire N__50255;
    wire N__50254;
    wire N__50253;
    wire N__50252;
    wire N__50251;
    wire N__50250;
    wire N__50249;
    wire N__50248;
    wire N__50247;
    wire N__50246;
    wire N__50245;
    wire N__50244;
    wire N__50243;
    wire N__50242;
    wire N__50241;
    wire N__50240;
    wire N__50239;
    wire N__50238;
    wire N__50237;
    wire N__50236;
    wire N__50235;
    wire N__50234;
    wire N__50233;
    wire N__50232;
    wire N__50231;
    wire N__50230;
    wire N__50229;
    wire N__50228;
    wire N__50227;
    wire N__50226;
    wire N__50225;
    wire N__50224;
    wire N__50223;
    wire N__50222;
    wire N__50221;
    wire N__50220;
    wire N__50219;
    wire N__50218;
    wire N__50217;
    wire N__50216;
    wire N__50215;
    wire N__50214;
    wire N__50213;
    wire N__50212;
    wire N__50211;
    wire N__50210;
    wire N__50209;
    wire N__50208;
    wire N__50207;
    wire N__50206;
    wire N__50205;
    wire N__50204;
    wire N__50203;
    wire N__50202;
    wire N__50201;
    wire N__50200;
    wire N__50199;
    wire N__50198;
    wire N__50197;
    wire N__50196;
    wire N__50195;
    wire N__50194;
    wire N__50193;
    wire N__50192;
    wire N__50191;
    wire N__50190;
    wire N__50189;
    wire N__50188;
    wire N__50187;
    wire N__50186;
    wire N__50185;
    wire N__50184;
    wire N__50183;
    wire N__50182;
    wire N__50181;
    wire N__50180;
    wire N__50179;
    wire N__50178;
    wire N__50177;
    wire N__50176;
    wire N__50175;
    wire N__50174;
    wire N__50173;
    wire N__50172;
    wire N__50171;
    wire N__50170;
    wire N__50169;
    wire N__50166;
    wire N__50165;
    wire N__49856;
    wire N__49853;
    wire N__49852;
    wire N__49851;
    wire N__49850;
    wire N__49849;
    wire N__49848;
    wire N__49847;
    wire N__49840;
    wire N__49839;
    wire N__49838;
    wire N__49837;
    wire N__49836;
    wire N__49835;
    wire N__49834;
    wire N__49833;
    wire N__49832;
    wire N__49823;
    wire N__49820;
    wire N__49811;
    wire N__49808;
    wire N__49807;
    wire N__49806;
    wire N__49805;
    wire N__49804;
    wire N__49803;
    wire N__49800;
    wire N__49799;
    wire N__49796;
    wire N__49793;
    wire N__49792;
    wire N__49791;
    wire N__49790;
    wire N__49789;
    wire N__49788;
    wire N__49781;
    wire N__49778;
    wire N__49777;
    wire N__49776;
    wire N__49775;
    wire N__49774;
    wire N__49773;
    wire N__49772;
    wire N__49771;
    wire N__49770;
    wire N__49769;
    wire N__49768;
    wire N__49767;
    wire N__49766;
    wire N__49763;
    wire N__49760;
    wire N__49757;
    wire N__49754;
    wire N__49751;
    wire N__49748;
    wire N__49747;
    wire N__49746;
    wire N__49745;
    wire N__49744;
    wire N__49741;
    wire N__49736;
    wire N__49735;
    wire N__49734;
    wire N__49733;
    wire N__49730;
    wire N__49727;
    wire N__49720;
    wire N__49715;
    wire N__49706;
    wire N__49697;
    wire N__49688;
    wire N__49685;
    wire N__49680;
    wire N__49677;
    wire N__49672;
    wire N__49663;
    wire N__49660;
    wire N__49657;
    wire N__49654;
    wire N__49651;
    wire N__49648;
    wire N__49645;
    wire N__49642;
    wire N__49631;
    wire N__49628;
    wire N__49625;
    wire N__49614;
    wire N__49611;
    wire N__49608;
    wire N__49603;
    wire N__49598;
    wire N__49595;
    wire N__49592;
    wire N__49589;
    wire N__49574;
    wire N__49573;
    wire N__49572;
    wire N__49571;
    wire N__49568;
    wire N__49565;
    wire N__49562;
    wire N__49559;
    wire N__49556;
    wire N__49553;
    wire N__49552;
    wire N__49551;
    wire N__49550;
    wire N__49549;
    wire N__49548;
    wire N__49545;
    wire N__49544;
    wire N__49541;
    wire N__49540;
    wire N__49539;
    wire N__49538;
    wire N__49537;
    wire N__49536;
    wire N__49535;
    wire N__49534;
    wire N__49533;
    wire N__49532;
    wire N__49531;
    wire N__49530;
    wire N__49529;
    wire N__49528;
    wire N__49527;
    wire N__49526;
    wire N__49525;
    wire N__49524;
    wire N__49523;
    wire N__49522;
    wire N__49521;
    wire N__49520;
    wire N__49519;
    wire N__49518;
    wire N__49517;
    wire N__49516;
    wire N__49515;
    wire N__49514;
    wire N__49513;
    wire N__49512;
    wire N__49511;
    wire N__49510;
    wire N__49509;
    wire N__49508;
    wire N__49507;
    wire N__49506;
    wire N__49505;
    wire N__49504;
    wire N__49503;
    wire N__49502;
    wire N__49501;
    wire N__49500;
    wire N__49499;
    wire N__49498;
    wire N__49497;
    wire N__49496;
    wire N__49495;
    wire N__49494;
    wire N__49493;
    wire N__49492;
    wire N__49491;
    wire N__49490;
    wire N__49489;
    wire N__49488;
    wire N__49487;
    wire N__49486;
    wire N__49485;
    wire N__49484;
    wire N__49483;
    wire N__49482;
    wire N__49481;
    wire N__49480;
    wire N__49479;
    wire N__49478;
    wire N__49477;
    wire N__49476;
    wire N__49475;
    wire N__49474;
    wire N__49473;
    wire N__49472;
    wire N__49471;
    wire N__49470;
    wire N__49469;
    wire N__49468;
    wire N__49467;
    wire N__49466;
    wire N__49465;
    wire N__49464;
    wire N__49463;
    wire N__49462;
    wire N__49461;
    wire N__49460;
    wire N__49459;
    wire N__49458;
    wire N__49457;
    wire N__49456;
    wire N__49455;
    wire N__49454;
    wire N__49453;
    wire N__49452;
    wire N__49451;
    wire N__49450;
    wire N__49449;
    wire N__49448;
    wire N__49447;
    wire N__49446;
    wire N__49445;
    wire N__49444;
    wire N__49443;
    wire N__49442;
    wire N__49441;
    wire N__49440;
    wire N__49439;
    wire N__49438;
    wire N__49437;
    wire N__49436;
    wire N__49435;
    wire N__49434;
    wire N__49433;
    wire N__49432;
    wire N__49431;
    wire N__49430;
    wire N__49429;
    wire N__49428;
    wire N__49427;
    wire N__49426;
    wire N__49425;
    wire N__49424;
    wire N__49423;
    wire N__49422;
    wire N__49421;
    wire N__49420;
    wire N__49419;
    wire N__49418;
    wire N__49417;
    wire N__49416;
    wire N__49415;
    wire N__49414;
    wire N__49413;
    wire N__49412;
    wire N__49411;
    wire N__49410;
    wire N__49409;
    wire N__49408;
    wire N__49407;
    wire N__49406;
    wire N__49405;
    wire N__49404;
    wire N__49403;
    wire N__49402;
    wire N__49401;
    wire N__49400;
    wire N__49399;
    wire N__49398;
    wire N__49397;
    wire N__49396;
    wire N__49395;
    wire N__49394;
    wire N__49393;
    wire N__49076;
    wire N__49073;
    wire N__49070;
    wire N__49067;
    wire N__49064;
    wire N__49061;
    wire N__49058;
    wire N__49055;
    wire N__49054;
    wire N__49049;
    wire N__49046;
    wire N__49045;
    wire N__49044;
    wire N__49039;
    wire N__49036;
    wire N__49033;
    wire N__49028;
    wire N__49027;
    wire N__49024;
    wire N__49021;
    wire N__49020;
    wire N__49015;
    wire N__49012;
    wire N__49009;
    wire N__49004;
    wire N__49003;
    wire N__48998;
    wire N__48995;
    wire N__48992;
    wire N__48989;
    wire N__48986;
    wire N__48983;
    wire N__48982;
    wire N__48979;
    wire N__48978;
    wire N__48975;
    wire N__48972;
    wire N__48969;
    wire N__48968;
    wire N__48965;
    wire N__48960;
    wire N__48957;
    wire N__48954;
    wire N__48949;
    wire N__48946;
    wire N__48943;
    wire N__48938;
    wire N__48937;
    wire N__48936;
    wire N__48935;
    wire N__48932;
    wire N__48931;
    wire N__48930;
    wire N__48927;
    wire N__48926;
    wire N__48925;
    wire N__48924;
    wire N__48923;
    wire N__48922;
    wire N__48921;
    wire N__48920;
    wire N__48911;
    wire N__48910;
    wire N__48909;
    wire N__48908;
    wire N__48907;
    wire N__48906;
    wire N__48905;
    wire N__48904;
    wire N__48903;
    wire N__48902;
    wire N__48901;
    wire N__48894;
    wire N__48893;
    wire N__48892;
    wire N__48891;
    wire N__48890;
    wire N__48889;
    wire N__48888;
    wire N__48887;
    wire N__48886;
    wire N__48885;
    wire N__48884;
    wire N__48881;
    wire N__48880;
    wire N__48879;
    wire N__48878;
    wire N__48877;
    wire N__48876;
    wire N__48875;
    wire N__48874;
    wire N__48873;
    wire N__48872;
    wire N__48871;
    wire N__48870;
    wire N__48869;
    wire N__48864;
    wire N__48863;
    wire N__48862;
    wire N__48861;
    wire N__48860;
    wire N__48859;
    wire N__48858;
    wire N__48857;
    wire N__48856;
    wire N__48855;
    wire N__48854;
    wire N__48851;
    wire N__48846;
    wire N__48843;
    wire N__48840;
    wire N__48839;
    wire N__48836;
    wire N__48835;
    wire N__48834;
    wire N__48833;
    wire N__48832;
    wire N__48831;
    wire N__48830;
    wire N__48829;
    wire N__48828;
    wire N__48827;
    wire N__48826;
    wire N__48823;
    wire N__48820;
    wire N__48817;
    wire N__48814;
    wire N__48805;
    wire N__48802;
    wire N__48795;
    wire N__48788;
    wire N__48779;
    wire N__48778;
    wire N__48777;
    wire N__48776;
    wire N__48773;
    wire N__48770;
    wire N__48765;
    wire N__48760;
    wire N__48759;
    wire N__48758;
    wire N__48757;
    wire N__48752;
    wire N__48749;
    wire N__48744;
    wire N__48739;
    wire N__48736;
    wire N__48727;
    wire N__48724;
    wire N__48719;
    wire N__48716;
    wire N__48711;
    wire N__48702;
    wire N__48699;
    wire N__48696;
    wire N__48693;
    wire N__48692;
    wire N__48691;
    wire N__48690;
    wire N__48689;
    wire N__48678;
    wire N__48677;
    wire N__48676;
    wire N__48675;
    wire N__48674;
    wire N__48673;
    wire N__48672;
    wire N__48671;
    wire N__48670;
    wire N__48669;
    wire N__48668;
    wire N__48667;
    wire N__48666;
    wire N__48665;
    wire N__48662;
    wire N__48657;
    wire N__48654;
    wire N__48653;
    wire N__48652;
    wire N__48651;
    wire N__48644;
    wire N__48631;
    wire N__48624;
    wire N__48619;
    wire N__48614;
    wire N__48607;
    wire N__48590;
    wire N__48583;
    wire N__48580;
    wire N__48575;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48549;
    wire N__48540;
    wire N__48533;
    wire N__48526;
    wire N__48519;
    wire N__48512;
    wire N__48507;
    wire N__48500;
    wire N__48495;
    wire N__48488;
    wire N__48467;
    wire N__48464;
    wire N__48463;
    wire N__48462;
    wire N__48459;
    wire N__48456;
    wire N__48453;
    wire N__48450;
    wire N__48447;
    wire N__48440;
    wire N__48439;
    wire N__48438;
    wire N__48437;
    wire N__48436;
    wire N__48435;
    wire N__48432;
    wire N__48431;
    wire N__48428;
    wire N__48425;
    wire N__48422;
    wire N__48419;
    wire N__48418;
    wire N__48417;
    wire N__48416;
    wire N__48415;
    wire N__48414;
    wire N__48413;
    wire N__48412;
    wire N__48411;
    wire N__48410;
    wire N__48409;
    wire N__48408;
    wire N__48407;
    wire N__48406;
    wire N__48405;
    wire N__48404;
    wire N__48397;
    wire N__48388;
    wire N__48381;
    wire N__48372;
    wire N__48371;
    wire N__48368;
    wire N__48363;
    wire N__48360;
    wire N__48355;
    wire N__48352;
    wire N__48349;
    wire N__48348;
    wire N__48345;
    wire N__48344;
    wire N__48343;
    wire N__48342;
    wire N__48341;
    wire N__48340;
    wire N__48339;
    wire N__48338;
    wire N__48337;
    wire N__48336;
    wire N__48335;
    wire N__48334;
    wire N__48333;
    wire N__48326;
    wire N__48323;
    wire N__48312;
    wire N__48309;
    wire N__48306;
    wire N__48305;
    wire N__48304;
    wire N__48303;
    wire N__48302;
    wire N__48301;
    wire N__48300;
    wire N__48299;
    wire N__48296;
    wire N__48295;
    wire N__48292;
    wire N__48291;
    wire N__48288;
    wire N__48287;
    wire N__48284;
    wire N__48283;
    wire N__48280;
    wire N__48279;
    wire N__48276;
    wire N__48275;
    wire N__48272;
    wire N__48271;
    wire N__48268;
    wire N__48267;
    wire N__48264;
    wire N__48263;
    wire N__48260;
    wire N__48259;
    wire N__48256;
    wire N__48255;
    wire N__48252;
    wire N__48251;
    wire N__48250;
    wire N__48249;
    wire N__48248;
    wire N__48245;
    wire N__48238;
    wire N__48235;
    wire N__48232;
    wire N__48225;
    wire N__48216;
    wire N__48213;
    wire N__48198;
    wire N__48181;
    wire N__48164;
    wire N__48163;
    wire N__48160;
    wire N__48159;
    wire N__48156;
    wire N__48155;
    wire N__48152;
    wire N__48151;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48139;
    wire N__48134;
    wire N__48129;
    wire N__48126;
    wire N__48123;
    wire N__48108;
    wire N__48105;
    wire N__48102;
    wire N__48095;
    wire N__48084;
    wire N__48081;
    wire N__48078;
    wire N__48075;
    wire N__48072;
    wire N__48065;
    wire N__48064;
    wire N__48063;
    wire N__48060;
    wire N__48057;
    wire N__48054;
    wire N__48051;
    wire N__48048;
    wire N__48047;
    wire N__48044;
    wire N__48041;
    wire N__48038;
    wire N__48035;
    wire N__48032;
    wire N__48027;
    wire N__48020;
    wire N__48017;
    wire N__48014;
    wire N__48013;
    wire N__48010;
    wire N__48007;
    wire N__48004;
    wire N__48001;
    wire N__48000;
    wire N__47997;
    wire N__47996;
    wire N__47993;
    wire N__47990;
    wire N__47987;
    wire N__47984;
    wire N__47981;
    wire N__47978;
    wire N__47969;
    wire N__47966;
    wire N__47963;
    wire N__47962;
    wire N__47959;
    wire N__47956;
    wire N__47953;
    wire N__47950;
    wire N__47945;
    wire N__47944;
    wire N__47943;
    wire N__47940;
    wire N__47937;
    wire N__47934;
    wire N__47931;
    wire N__47924;
    wire N__47923;
    wire N__47922;
    wire N__47919;
    wire N__47916;
    wire N__47913;
    wire N__47908;
    wire N__47907;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47891;
    wire N__47890;
    wire N__47885;
    wire N__47882;
    wire N__47879;
    wire N__47876;
    wire N__47873;
    wire N__47872;
    wire N__47871;
    wire N__47870;
    wire N__47869;
    wire N__47868;
    wire N__47867;
    wire N__47866;
    wire N__47865;
    wire N__47864;
    wire N__47863;
    wire N__47862;
    wire N__47861;
    wire N__47860;
    wire N__47831;
    wire N__47828;
    wire N__47825;
    wire N__47824;
    wire N__47823;
    wire N__47820;
    wire N__47817;
    wire N__47814;
    wire N__47807;
    wire N__47804;
    wire N__47803;
    wire N__47802;
    wire N__47799;
    wire N__47796;
    wire N__47793;
    wire N__47792;
    wire N__47789;
    wire N__47784;
    wire N__47781;
    wire N__47778;
    wire N__47775;
    wire N__47772;
    wire N__47765;
    wire N__47764;
    wire N__47759;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47749;
    wire N__47748;
    wire N__47745;
    wire N__47742;
    wire N__47739;
    wire N__47734;
    wire N__47729;
    wire N__47728;
    wire N__47727;
    wire N__47724;
    wire N__47721;
    wire N__47720;
    wire N__47717;
    wire N__47714;
    wire N__47711;
    wire N__47708;
    wire N__47705;
    wire N__47700;
    wire N__47697;
    wire N__47690;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47675;
    wire N__47672;
    wire N__47669;
    wire N__47668;
    wire N__47665;
    wire N__47662;
    wire N__47657;
    wire N__47656;
    wire N__47655;
    wire N__47650;
    wire N__47647;
    wire N__47644;
    wire N__47643;
    wire N__47640;
    wire N__47637;
    wire N__47634;
    wire N__47629;
    wire N__47626;
    wire N__47621;
    wire N__47618;
    wire N__47617;
    wire N__47612;
    wire N__47609;
    wire N__47608;
    wire N__47603;
    wire N__47602;
    wire N__47599;
    wire N__47596;
    wire N__47593;
    wire N__47588;
    wire N__47587;
    wire N__47584;
    wire N__47581;
    wire N__47576;
    wire N__47575;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47561;
    wire N__47560;
    wire N__47555;
    wire N__47552;
    wire N__47549;
    wire N__47546;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47533;
    wire N__47530;
    wire N__47527;
    wire N__47522;
    wire N__47521;
    wire N__47520;
    wire N__47515;
    wire N__47512;
    wire N__47509;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47492;
    wire N__47489;
    wire N__47486;
    wire N__47483;
    wire N__47480;
    wire N__47477;
    wire N__47476;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47466;
    wire N__47461;
    wire N__47456;
    wire N__47455;
    wire N__47452;
    wire N__47449;
    wire N__47448;
    wire N__47447;
    wire N__47444;
    wire N__47441;
    wire N__47438;
    wire N__47435;
    wire N__47430;
    wire N__47427;
    wire N__47424;
    wire N__47419;
    wire N__47416;
    wire N__47413;
    wire N__47408;
    wire N__47405;
    wire N__47402;
    wire N__47399;
    wire N__47396;
    wire N__47395;
    wire N__47394;
    wire N__47389;
    wire N__47386;
    wire N__47383;
    wire N__47378;
    wire N__47375;
    wire N__47374;
    wire N__47373;
    wire N__47368;
    wire N__47365;
    wire N__47362;
    wire N__47357;
    wire N__47354;
    wire N__47353;
    wire N__47348;
    wire N__47345;
    wire N__47342;
    wire N__47339;
    wire N__47336;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47324;
    wire N__47323;
    wire N__47320;
    wire N__47317;
    wire N__47312;
    wire N__47311;
    wire N__47306;
    wire N__47305;
    wire N__47302;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47284;
    wire N__47281;
    wire N__47278;
    wire N__47273;
    wire N__47270;
    wire N__47269;
    wire N__47264;
    wire N__47261;
    wire N__47260;
    wire N__47255;
    wire N__47252;
    wire N__47249;
    wire N__47248;
    wire N__47245;
    wire N__47242;
    wire N__47237;
    wire N__47234;
    wire N__47231;
    wire N__47228;
    wire N__47227;
    wire N__47224;
    wire N__47221;
    wire N__47216;
    wire N__47215;
    wire N__47210;
    wire N__47209;
    wire N__47206;
    wire N__47203;
    wire N__47200;
    wire N__47199;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47183;
    wire N__47180;
    wire N__47179;
    wire N__47178;
    wire N__47175;
    wire N__47170;
    wire N__47165;
    wire N__47162;
    wire N__47161;
    wire N__47158;
    wire N__47155;
    wire N__47150;
    wire N__47149;
    wire N__47146;
    wire N__47143;
    wire N__47140;
    wire N__47135;
    wire N__47132;
    wire N__47131;
    wire N__47126;
    wire N__47123;
    wire N__47120;
    wire N__47117;
    wire N__47114;
    wire N__47111;
    wire N__47108;
    wire N__47107;
    wire N__47104;
    wire N__47101;
    wire N__47098;
    wire N__47093;
    wire N__47092;
    wire N__47091;
    wire N__47086;
    wire N__47083;
    wire N__47080;
    wire N__47079;
    wire N__47076;
    wire N__47073;
    wire N__47070;
    wire N__47063;
    wire N__47060;
    wire N__47057;
    wire N__47054;
    wire N__47051;
    wire N__47048;
    wire N__47047;
    wire N__47042;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47032;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47018;
    wire N__47015;
    wire N__47012;
    wire N__47009;
    wire N__47006;
    wire N__47003;
    wire N__47002;
    wire N__46999;
    wire N__46996;
    wire N__46993;
    wire N__46988;
    wire N__46987;
    wire N__46986;
    wire N__46985;
    wire N__46982;
    wire N__46981;
    wire N__46974;
    wire N__46971;
    wire N__46968;
    wire N__46965;
    wire N__46958;
    wire N__46957;
    wire N__46954;
    wire N__46951;
    wire N__46950;
    wire N__46947;
    wire N__46942;
    wire N__46939;
    wire N__46936;
    wire N__46931;
    wire N__46930;
    wire N__46927;
    wire N__46926;
    wire N__46923;
    wire N__46920;
    wire N__46917;
    wire N__46916;
    wire N__46913;
    wire N__46910;
    wire N__46907;
    wire N__46904;
    wire N__46901;
    wire N__46896;
    wire N__46895;
    wire N__46894;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46880;
    wire N__46871;
    wire N__46868;
    wire N__46865;
    wire N__46862;
    wire N__46859;
    wire N__46856;
    wire N__46853;
    wire N__46852;
    wire N__46851;
    wire N__46850;
    wire N__46845;
    wire N__46840;
    wire N__46835;
    wire N__46834;
    wire N__46833;
    wire N__46828;
    wire N__46825;
    wire N__46822;
    wire N__46821;
    wire N__46820;
    wire N__46817;
    wire N__46814;
    wire N__46809;
    wire N__46802;
    wire N__46799;
    wire N__46796;
    wire N__46793;
    wire N__46790;
    wire N__46787;
    wire N__46784;
    wire N__46781;
    wire N__46778;
    wire N__46777;
    wire N__46776;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46762;
    wire N__46757;
    wire N__46754;
    wire N__46751;
    wire N__46748;
    wire N__46747;
    wire N__46744;
    wire N__46741;
    wire N__46740;
    wire N__46735;
    wire N__46732;
    wire N__46729;
    wire N__46724;
    wire N__46721;
    wire N__46718;
    wire N__46717;
    wire N__46714;
    wire N__46711;
    wire N__46708;
    wire N__46703;
    wire N__46700;
    wire N__46699;
    wire N__46698;
    wire N__46697;
    wire N__46696;
    wire N__46695;
    wire N__46694;
    wire N__46693;
    wire N__46684;
    wire N__46675;
    wire N__46674;
    wire N__46673;
    wire N__46672;
    wire N__46671;
    wire N__46670;
    wire N__46669;
    wire N__46668;
    wire N__46667;
    wire N__46666;
    wire N__46665;
    wire N__46664;
    wire N__46663;
    wire N__46662;
    wire N__46661;
    wire N__46660;
    wire N__46659;
    wire N__46658;
    wire N__46657;
    wire N__46656;
    wire N__46655;
    wire N__46654;
    wire N__46653;
    wire N__46648;
    wire N__46639;
    wire N__46634;
    wire N__46625;
    wire N__46616;
    wire N__46607;
    wire N__46598;
    wire N__46591;
    wire N__46582;
    wire N__46577;
    wire N__46574;
    wire N__46571;
    wire N__46568;
    wire N__46567;
    wire N__46564;
    wire N__46561;
    wire N__46558;
    wire N__46553;
    wire N__46552;
    wire N__46551;
    wire N__46548;
    wire N__46545;
    wire N__46544;
    wire N__46541;
    wire N__46538;
    wire N__46535;
    wire N__46532;
    wire N__46529;
    wire N__46526;
    wire N__46523;
    wire N__46520;
    wire N__46517;
    wire N__46514;
    wire N__46509;
    wire N__46502;
    wire N__46499;
    wire N__46498;
    wire N__46495;
    wire N__46492;
    wire N__46487;
    wire N__46484;
    wire N__46483;
    wire N__46480;
    wire N__46477;
    wire N__46476;
    wire N__46471;
    wire N__46468;
    wire N__46465;
    wire N__46460;
    wire N__46459;
    wire N__46458;
    wire N__46455;
    wire N__46452;
    wire N__46449;
    wire N__46448;
    wire N__46445;
    wire N__46442;
    wire N__46439;
    wire N__46436;
    wire N__46431;
    wire N__46428;
    wire N__46421;
    wire N__46418;
    wire N__46415;
    wire N__46414;
    wire N__46413;
    wire N__46410;
    wire N__46409;
    wire N__46406;
    wire N__46403;
    wire N__46400;
    wire N__46397;
    wire N__46394;
    wire N__46385;
    wire N__46384;
    wire N__46383;
    wire N__46380;
    wire N__46379;
    wire N__46376;
    wire N__46373;
    wire N__46370;
    wire N__46367;
    wire N__46364;
    wire N__46361;
    wire N__46358;
    wire N__46355;
    wire N__46350;
    wire N__46347;
    wire N__46340;
    wire N__46339;
    wire N__46336;
    wire N__46335;
    wire N__46332;
    wire N__46331;
    wire N__46328;
    wire N__46325;
    wire N__46322;
    wire N__46319;
    wire N__46316;
    wire N__46309;
    wire N__46304;
    wire N__46301;
    wire N__46298;
    wire N__46297;
    wire N__46296;
    wire N__46293;
    wire N__46290;
    wire N__46287;
    wire N__46282;
    wire N__46277;
    wire N__46274;
    wire N__46271;
    wire N__46270;
    wire N__46265;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46250;
    wire N__46247;
    wire N__46244;
    wire N__46243;
    wire N__46240;
    wire N__46237;
    wire N__46236;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46220;
    wire N__46217;
    wire N__46216;
    wire N__46213;
    wire N__46210;
    wire N__46205;
    wire N__46204;
    wire N__46201;
    wire N__46198;
    wire N__46195;
    wire N__46190;
    wire N__46187;
    wire N__46186;
    wire N__46181;
    wire N__46180;
    wire N__46177;
    wire N__46174;
    wire N__46171;
    wire N__46166;
    wire N__46163;
    wire N__46162;
    wire N__46157;
    wire N__46156;
    wire N__46153;
    wire N__46150;
    wire N__46147;
    wire N__46142;
    wire N__46139;
    wire N__46138;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46126;
    wire N__46125;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46103;
    wire N__46100;
    wire N__46099;
    wire N__46096;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46064;
    wire N__46061;
    wire N__46058;
    wire N__46057;
    wire N__46054;
    wire N__46051;
    wire N__46050;
    wire N__46047;
    wire N__46044;
    wire N__46041;
    wire N__46038;
    wire N__46035;
    wire N__46028;
    wire N__46025;
    wire N__46024;
    wire N__46023;
    wire N__46018;
    wire N__46015;
    wire N__46012;
    wire N__46007;
    wire N__46004;
    wire N__46001;
    wire N__46000;
    wire N__45995;
    wire N__45994;
    wire N__45991;
    wire N__45988;
    wire N__45985;
    wire N__45980;
    wire N__45977;
    wire N__45976;
    wire N__45973;
    wire N__45970;
    wire N__45965;
    wire N__45964;
    wire N__45961;
    wire N__45958;
    wire N__45955;
    wire N__45950;
    wire N__45947;
    wire N__45946;
    wire N__45943;
    wire N__45940;
    wire N__45935;
    wire N__45934;
    wire N__45931;
    wire N__45928;
    wire N__45925;
    wire N__45920;
    wire N__45917;
    wire N__45916;
    wire N__45911;
    wire N__45910;
    wire N__45907;
    wire N__45904;
    wire N__45901;
    wire N__45896;
    wire N__45893;
    wire N__45890;
    wire N__45889;
    wire N__45886;
    wire N__45883;
    wire N__45882;
    wire N__45877;
    wire N__45874;
    wire N__45871;
    wire N__45866;
    wire N__45863;
    wire N__45862;
    wire N__45859;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45849;
    wire N__45846;
    wire N__45843;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45820;
    wire N__45817;
    wire N__45814;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45798;
    wire N__45791;
    wire N__45790;
    wire N__45787;
    wire N__45784;
    wire N__45783;
    wire N__45780;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45764;
    wire N__45761;
    wire N__45760;
    wire N__45757;
    wire N__45754;
    wire N__45753;
    wire N__45748;
    wire N__45745;
    wire N__45742;
    wire N__45737;
    wire N__45734;
    wire N__45731;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45719;
    wire N__45718;
    wire N__45715;
    wire N__45712;
    wire N__45709;
    wire N__45704;
    wire N__45701;
    wire N__45698;
    wire N__45697;
    wire N__45694;
    wire N__45691;
    wire N__45690;
    wire N__45685;
    wire N__45682;
    wire N__45679;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45667;
    wire N__45664;
    wire N__45661;
    wire N__45660;
    wire N__45655;
    wire N__45652;
    wire N__45649;
    wire N__45644;
    wire N__45641;
    wire N__45638;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45630;
    wire N__45625;
    wire N__45622;
    wire N__45619;
    wire N__45614;
    wire N__45611;
    wire N__45608;
    wire N__45607;
    wire N__45604;
    wire N__45601;
    wire N__45600;
    wire N__45595;
    wire N__45592;
    wire N__45589;
    wire N__45584;
    wire N__45581;
    wire N__45578;
    wire N__45577;
    wire N__45574;
    wire N__45571;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45555;
    wire N__45548;
    wire N__45545;
    wire N__45544;
    wire N__45539;
    wire N__45536;
    wire N__45533;
    wire N__45532;
    wire N__45527;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45512;
    wire N__45511;
    wire N__45506;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45496;
    wire N__45491;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45481;
    wire N__45480;
    wire N__45477;
    wire N__45474;
    wire N__45471;
    wire N__45468;
    wire N__45461;
    wire N__45458;
    wire N__45455;
    wire N__45454;
    wire N__45453;
    wire N__45452;
    wire N__45451;
    wire N__45450;
    wire N__45449;
    wire N__45448;
    wire N__45447;
    wire N__45446;
    wire N__45445;
    wire N__45444;
    wire N__45443;
    wire N__45442;
    wire N__45441;
    wire N__45440;
    wire N__45439;
    wire N__45438;
    wire N__45437;
    wire N__45436;
    wire N__45435;
    wire N__45434;
    wire N__45433;
    wire N__45432;
    wire N__45431;
    wire N__45426;
    wire N__45425;
    wire N__45424;
    wire N__45419;
    wire N__45418;
    wire N__45417;
    wire N__45416;
    wire N__45415;
    wire N__45414;
    wire N__45411;
    wire N__45410;
    wire N__45409;
    wire N__45408;
    wire N__45407;
    wire N__45406;
    wire N__45405;
    wire N__45404;
    wire N__45401;
    wire N__45400;
    wire N__45399;
    wire N__45398;
    wire N__45397;
    wire N__45396;
    wire N__45393;
    wire N__45392;
    wire N__45391;
    wire N__45390;
    wire N__45387;
    wire N__45386;
    wire N__45385;
    wire N__45384;
    wire N__45383;
    wire N__45382;
    wire N__45379;
    wire N__45378;
    wire N__45377;
    wire N__45376;
    wire N__45369;
    wire N__45362;
    wire N__45359;
    wire N__45352;
    wire N__45339;
    wire N__45336;
    wire N__45335;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45319;
    wire N__45304;
    wire N__45297;
    wire N__45294;
    wire N__45285;
    wire N__45284;
    wire N__45283;
    wire N__45282;
    wire N__45281;
    wire N__45280;
    wire N__45279;
    wire N__45278;
    wire N__45277;
    wire N__45262;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45236;
    wire N__45233;
    wire N__45228;
    wire N__45225;
    wire N__45224;
    wire N__45223;
    wire N__45222;
    wire N__45221;
    wire N__45220;
    wire N__45219;
    wire N__45218;
    wire N__45209;
    wire N__45206;
    wire N__45203;
    wire N__45198;
    wire N__45195;
    wire N__45190;
    wire N__45185;
    wire N__45178;
    wire N__45173;
    wire N__45170;
    wire N__45165;
    wire N__45158;
    wire N__45151;
    wire N__45142;
    wire N__45139;
    wire N__45132;
    wire N__45107;
    wire N__45104;
    wire N__45103;
    wire N__45102;
    wire N__45101;
    wire N__45098;
    wire N__45095;
    wire N__45090;
    wire N__45083;
    wire N__45080;
    wire N__45077;
    wire N__45076;
    wire N__45073;
    wire N__45070;
    wire N__45067;
    wire N__45062;
    wire N__45059;
    wire N__45058;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45044;
    wire N__45043;
    wire N__45042;
    wire N__45041;
    wire N__45038;
    wire N__45035;
    wire N__45034;
    wire N__45033;
    wire N__45028;
    wire N__45023;
    wire N__45020;
    wire N__45017;
    wire N__45014;
    wire N__45011;
    wire N__45002;
    wire N__45001;
    wire N__44998;
    wire N__44997;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44982;
    wire N__44979;
    wire N__44976;
    wire N__44971;
    wire N__44966;
    wire N__44963;
    wire N__44960;
    wire N__44959;
    wire N__44958;
    wire N__44957;
    wire N__44956;
    wire N__44955;
    wire N__44954;
    wire N__44953;
    wire N__44936;
    wire N__44933;
    wire N__44930;
    wire N__44929;
    wire N__44928;
    wire N__44923;
    wire N__44920;
    wire N__44917;
    wire N__44916;
    wire N__44915;
    wire N__44914;
    wire N__44913;
    wire N__44912;
    wire N__44911;
    wire N__44910;
    wire N__44909;
    wire N__44908;
    wire N__44907;
    wire N__44906;
    wire N__44905;
    wire N__44904;
    wire N__44903;
    wire N__44902;
    wire N__44901;
    wire N__44900;
    wire N__44899;
    wire N__44898;
    wire N__44893;
    wire N__44884;
    wire N__44873;
    wire N__44866;
    wire N__44865;
    wire N__44864;
    wire N__44863;
    wire N__44860;
    wire N__44849;
    wire N__44846;
    wire N__44837;
    wire N__44834;
    wire N__44829;
    wire N__44816;
    wire N__44813;
    wire N__44812;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44802;
    wire N__44799;
    wire N__44794;
    wire N__44789;
    wire N__44786;
    wire N__44783;
    wire N__44780;
    wire N__44777;
    wire N__44776;
    wire N__44775;
    wire N__44774;
    wire N__44771;
    wire N__44768;
    wire N__44763;
    wire N__44760;
    wire N__44757;
    wire N__44754;
    wire N__44751;
    wire N__44746;
    wire N__44741;
    wire N__44738;
    wire N__44735;
    wire N__44732;
    wire N__44731;
    wire N__44728;
    wire N__44725;
    wire N__44724;
    wire N__44721;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44705;
    wire N__44702;
    wire N__44699;
    wire N__44696;
    wire N__44693;
    wire N__44692;
    wire N__44689;
    wire N__44686;
    wire N__44681;
    wire N__44680;
    wire N__44677;
    wire N__44674;
    wire N__44671;
    wire N__44666;
    wire N__44663;
    wire N__44660;
    wire N__44659;
    wire N__44654;
    wire N__44653;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44639;
    wire N__44636;
    wire N__44633;
    wire N__44630;
    wire N__44627;
    wire N__44624;
    wire N__44623;
    wire N__44620;
    wire N__44615;
    wire N__44614;
    wire N__44611;
    wire N__44608;
    wire N__44605;
    wire N__44600;
    wire N__44597;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44589;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44561;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44549;
    wire N__44548;
    wire N__44547;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44531;
    wire N__44528;
    wire N__44527;
    wire N__44526;
    wire N__44521;
    wire N__44518;
    wire N__44515;
    wire N__44510;
    wire N__44507;
    wire N__44506;
    wire N__44503;
    wire N__44502;
    wire N__44497;
    wire N__44494;
    wire N__44491;
    wire N__44486;
    wire N__44483;
    wire N__44480;
    wire N__44479;
    wire N__44478;
    wire N__44475;
    wire N__44472;
    wire N__44469;
    wire N__44464;
    wire N__44459;
    wire N__44456;
    wire N__44453;
    wire N__44450;
    wire N__44449;
    wire N__44448;
    wire N__44445;
    wire N__44440;
    wire N__44435;
    wire N__44432;
    wire N__44431;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44419;
    wire N__44414;
    wire N__44411;
    wire N__44408;
    wire N__44407;
    wire N__44404;
    wire N__44401;
    wire N__44396;
    wire N__44393;
    wire N__44392;
    wire N__44389;
    wire N__44386;
    wire N__44381;
    wire N__44378;
    wire N__44375;
    wire N__44374;
    wire N__44371;
    wire N__44368;
    wire N__44365;
    wire N__44360;
    wire N__44357;
    wire N__44356;
    wire N__44353;
    wire N__44350;
    wire N__44345;
    wire N__44342;
    wire N__44341;
    wire N__44338;
    wire N__44335;
    wire N__44330;
    wire N__44327;
    wire N__44326;
    wire N__44323;
    wire N__44320;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44306;
    wire N__44303;
    wire N__44300;
    wire N__44297;
    wire N__44296;
    wire N__44293;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44267;
    wire N__44266;
    wire N__44263;
    wire N__44260;
    wire N__44255;
    wire N__44252;
    wire N__44249;
    wire N__44246;
    wire N__44243;
    wire N__44242;
    wire N__44239;
    wire N__44236;
    wire N__44231;
    wire N__44228;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44216;
    wire N__44213;
    wire N__44212;
    wire N__44209;
    wire N__44206;
    wire N__44201;
    wire N__44198;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44186;
    wire N__44183;
    wire N__44182;
    wire N__44179;
    wire N__44176;
    wire N__44171;
    wire N__44168;
    wire N__44167;
    wire N__44164;
    wire N__44161;
    wire N__44156;
    wire N__44153;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44141;
    wire N__44138;
    wire N__44135;
    wire N__44132;
    wire N__44129;
    wire N__44126;
    wire N__44123;
    wire N__44120;
    wire N__44119;
    wire N__44116;
    wire N__44113;
    wire N__44108;
    wire N__44105;
    wire N__44104;
    wire N__44103;
    wire N__44100;
    wire N__44095;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44085;
    wire N__44080;
    wire N__44077;
    wire N__44072;
    wire N__44071;
    wire N__44068;
    wire N__44063;
    wire N__44060;
    wire N__44059;
    wire N__44056;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44039;
    wire N__44036;
    wire N__44035;
    wire N__44032;
    wire N__44029;
    wire N__44028;
    wire N__44027;
    wire N__44022;
    wire N__44017;
    wire N__44012;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__44002;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43985;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43973;
    wire N__43972;
    wire N__43967;
    wire N__43964;
    wire N__43963;
    wire N__43960;
    wire N__43957;
    wire N__43952;
    wire N__43949;
    wire N__43946;
    wire N__43943;
    wire N__43940;
    wire N__43939;
    wire N__43938;
    wire N__43935;
    wire N__43932;
    wire N__43929;
    wire N__43926;
    wire N__43923;
    wire N__43920;
    wire N__43919;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43907;
    wire N__43904;
    wire N__43901;
    wire N__43898;
    wire N__43889;
    wire N__43886;
    wire N__43885;
    wire N__43882;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43865;
    wire N__43862;
    wire N__43861;
    wire N__43858;
    wire N__43855;
    wire N__43854;
    wire N__43851;
    wire N__43848;
    wire N__43845;
    wire N__43838;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43828;
    wire N__43825;
    wire N__43824;
    wire N__43821;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43805;
    wire N__43802;
    wire N__43801;
    wire N__43800;
    wire N__43797;
    wire N__43794;
    wire N__43793;
    wire N__43792;
    wire N__43789;
    wire N__43784;
    wire N__43781;
    wire N__43778;
    wire N__43775;
    wire N__43772;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43758;
    wire N__43755;
    wire N__43748;
    wire N__43745;
    wire N__43744;
    wire N__43741;
    wire N__43740;
    wire N__43737;
    wire N__43734;
    wire N__43731;
    wire N__43724;
    wire N__43721;
    wire N__43720;
    wire N__43717;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43700;
    wire N__43697;
    wire N__43696;
    wire N__43693;
    wire N__43692;
    wire N__43689;
    wire N__43686;
    wire N__43683;
    wire N__43676;
    wire N__43673;
    wire N__43670;
    wire N__43667;
    wire N__43664;
    wire N__43661;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43649;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43637;
    wire N__43634;
    wire N__43631;
    wire N__43628;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43610;
    wire N__43607;
    wire N__43604;
    wire N__43601;
    wire N__43598;
    wire N__43595;
    wire N__43592;
    wire N__43591;
    wire N__43590;
    wire N__43589;
    wire N__43586;
    wire N__43583;
    wire N__43582;
    wire N__43581;
    wire N__43580;
    wire N__43579;
    wire N__43578;
    wire N__43577;
    wire N__43576;
    wire N__43575;
    wire N__43574;
    wire N__43573;
    wire N__43572;
    wire N__43571;
    wire N__43568;
    wire N__43567;
    wire N__43566;
    wire N__43563;
    wire N__43562;
    wire N__43561;
    wire N__43560;
    wire N__43559;
    wire N__43558;
    wire N__43557;
    wire N__43556;
    wire N__43555;
    wire N__43554;
    wire N__43553;
    wire N__43552;
    wire N__43551;
    wire N__43546;
    wire N__43543;
    wire N__43532;
    wire N__43529;
    wire N__43520;
    wire N__43517;
    wire N__43516;
    wire N__43515;
    wire N__43512;
    wire N__43501;
    wire N__43496;
    wire N__43491;
    wire N__43488;
    wire N__43477;
    wire N__43466;
    wire N__43463;
    wire N__43458;
    wire N__43451;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43433;
    wire N__43430;
    wire N__43427;
    wire N__43424;
    wire N__43419;
    wire N__43412;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43394;
    wire N__43391;
    wire N__43388;
    wire N__43385;
    wire N__43382;
    wire N__43379;
    wire N__43376;
    wire N__43373;
    wire N__43370;
    wire N__43367;
    wire N__43364;
    wire N__43361;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43349;
    wire N__43346;
    wire N__43343;
    wire N__43340;
    wire N__43337;
    wire N__43334;
    wire N__43331;
    wire N__43328;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43310;
    wire N__43307;
    wire N__43304;
    wire N__43301;
    wire N__43298;
    wire N__43295;
    wire N__43292;
    wire N__43289;
    wire N__43286;
    wire N__43283;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43259;
    wire N__43256;
    wire N__43253;
    wire N__43250;
    wire N__43247;
    wire N__43244;
    wire N__43241;
    wire N__43238;
    wire N__43235;
    wire N__43232;
    wire N__43229;
    wire N__43226;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43214;
    wire N__43211;
    wire N__43208;
    wire N__43205;
    wire N__43202;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43187;
    wire N__43184;
    wire N__43181;
    wire N__43178;
    wire N__43175;
    wire N__43172;
    wire N__43169;
    wire N__43166;
    wire N__43163;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43148;
    wire N__43145;
    wire N__43142;
    wire N__43139;
    wire N__43138;
    wire N__43137;
    wire N__43136;
    wire N__43133;
    wire N__43130;
    wire N__43125;
    wire N__43122;
    wire N__43119;
    wire N__43116;
    wire N__43113;
    wire N__43108;
    wire N__43105;
    wire N__43102;
    wire N__43097;
    wire N__43094;
    wire N__43091;
    wire N__43090;
    wire N__43089;
    wire N__43086;
    wire N__43083;
    wire N__43080;
    wire N__43073;
    wire N__43070;
    wire N__43069;
    wire N__43068;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43055;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43041;
    wire N__43034;
    wire N__43033;
    wire N__43030;
    wire N__43029;
    wire N__43026;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43008;
    wire N__43001;
    wire N__43000;
    wire N__42997;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42975;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42952;
    wire N__42949;
    wire N__42948;
    wire N__42945;
    wire N__42940;
    wire N__42935;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42911;
    wire N__42910;
    wire N__42909;
    wire N__42908;
    wire N__42907;
    wire N__42906;
    wire N__42903;
    wire N__42902;
    wire N__42899;
    wire N__42898;
    wire N__42897;
    wire N__42896;
    wire N__42895;
    wire N__42894;
    wire N__42893;
    wire N__42892;
    wire N__42891;
    wire N__42890;
    wire N__42889;
    wire N__42888;
    wire N__42887;
    wire N__42884;
    wire N__42883;
    wire N__42882;
    wire N__42881;
    wire N__42880;
    wire N__42879;
    wire N__42878;
    wire N__42877;
    wire N__42876;
    wire N__42871;
    wire N__42866;
    wire N__42865;
    wire N__42864;
    wire N__42863;
    wire N__42862;
    wire N__42861;
    wire N__42860;
    wire N__42859;
    wire N__42858;
    wire N__42857;
    wire N__42856;
    wire N__42855;
    wire N__42854;
    wire N__42851;
    wire N__42848;
    wire N__42847;
    wire N__42846;
    wire N__42843;
    wire N__42842;
    wire N__42841;
    wire N__42840;
    wire N__42839;
    wire N__42838;
    wire N__42837;
    wire N__42834;
    wire N__42833;
    wire N__42832;
    wire N__42831;
    wire N__42828;
    wire N__42827;
    wire N__42826;
    wire N__42825;
    wire N__42824;
    wire N__42823;
    wire N__42820;
    wire N__42819;
    wire N__42816;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42808;
    wire N__42805;
    wire N__42804;
    wire N__42801;
    wire N__42800;
    wire N__42797;
    wire N__42796;
    wire N__42795;
    wire N__42794;
    wire N__42793;
    wire N__42792;
    wire N__42789;
    wire N__42788;
    wire N__42787;
    wire N__42786;
    wire N__42785;
    wire N__42784;
    wire N__42783;
    wire N__42782;
    wire N__42781;
    wire N__42780;
    wire N__42779;
    wire N__42778;
    wire N__42773;
    wire N__42772;
    wire N__42771;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42757;
    wire N__42754;
    wire N__42753;
    wire N__42750;
    wire N__42749;
    wire N__42746;
    wire N__42745;
    wire N__42740;
    wire N__42737;
    wire N__42734;
    wire N__42731;
    wire N__42730;
    wire N__42727;
    wire N__42724;
    wire N__42723;
    wire N__42722;
    wire N__42721;
    wire N__42720;
    wire N__42719;
    wire N__42718;
    wire N__42717;
    wire N__42716;
    wire N__42713;
    wire N__42710;
    wire N__42697;
    wire N__42694;
    wire N__42689;
    wire N__42674;
    wire N__42659;
    wire N__42656;
    wire N__42641;
    wire N__42624;
    wire N__42621;
    wire N__42620;
    wire N__42617;
    wire N__42616;
    wire N__42613;
    wire N__42612;
    wire N__42609;
    wire N__42608;
    wire N__42607;
    wire N__42606;
    wire N__42605;
    wire N__42602;
    wire N__42595;
    wire N__42592;
    wire N__42591;
    wire N__42588;
    wire N__42587;
    wire N__42584;
    wire N__42583;
    wire N__42580;
    wire N__42579;
    wire N__42576;
    wire N__42575;
    wire N__42572;
    wire N__42571;
    wire N__42568;
    wire N__42567;
    wire N__42564;
    wire N__42563;
    wire N__42560;
    wire N__42553;
    wire N__42550;
    wire N__42545;
    wire N__42532;
    wire N__42529;
    wire N__42524;
    wire N__42513;
    wire N__42512;
    wire N__42511;
    wire N__42508;
    wire N__42505;
    wire N__42504;
    wire N__42503;
    wire N__42502;
    wire N__42499;
    wire N__42498;
    wire N__42495;
    wire N__42494;
    wire N__42491;
    wire N__42490;
    wire N__42487;
    wire N__42486;
    wire N__42483;
    wire N__42482;
    wire N__42475;
    wire N__42460;
    wire N__42443;
    wire N__42440;
    wire N__42439;
    wire N__42436;
    wire N__42435;
    wire N__42432;
    wire N__42431;
    wire N__42426;
    wire N__42423;
    wire N__42408;
    wire N__42391;
    wire N__42380;
    wire N__42377;
    wire N__42372;
    wire N__42359;
    wire N__42352;
    wire N__42335;
    wire N__42328;
    wire N__42315;
    wire N__42304;
    wire N__42287;
    wire N__42286;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42276;
    wire N__42273;
    wire N__42270;
    wire N__42263;
    wire N__42260;
    wire N__42257;
    wire N__42256;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42245;
    wire N__42242;
    wire N__42239;
    wire N__42236;
    wire N__42233;
    wire N__42224;
    wire N__42221;
    wire N__42218;
    wire N__42215;
    wire N__42212;
    wire N__42209;
    wire N__42208;
    wire N__42205;
    wire N__42202;
    wire N__42199;
    wire N__42198;
    wire N__42195;
    wire N__42192;
    wire N__42189;
    wire N__42188;
    wire N__42185;
    wire N__42180;
    wire N__42177;
    wire N__42170;
    wire N__42169;
    wire N__42166;
    wire N__42163;
    wire N__42162;
    wire N__42159;
    wire N__42156;
    wire N__42153;
    wire N__42146;
    wire N__42145;
    wire N__42142;
    wire N__42139;
    wire N__42136;
    wire N__42133;
    wire N__42132;
    wire N__42131;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42113;
    wire N__42110;
    wire N__42109;
    wire N__42108;
    wire N__42105;
    wire N__42102;
    wire N__42099;
    wire N__42094;
    wire N__42091;
    wire N__42086;
    wire N__42083;
    wire N__42080;
    wire N__42077;
    wire N__42076;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42066;
    wire N__42065;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42047;
    wire N__42044;
    wire N__42041;
    wire N__42038;
    wire N__42035;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42023;
    wire N__42022;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42007;
    wire N__42004;
    wire N__41999;
    wire N__41998;
    wire N__41993;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41981;
    wire N__41978;
    wire N__41975;
    wire N__41974;
    wire N__41971;
    wire N__41968;
    wire N__41965;
    wire N__41962;
    wire N__41959;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41948;
    wire N__41945;
    wire N__41942;
    wire N__41939;
    wire N__41936;
    wire N__41927;
    wire N__41926;
    wire N__41923;
    wire N__41920;
    wire N__41917;
    wire N__41916;
    wire N__41911;
    wire N__41908;
    wire N__41903;
    wire N__41900;
    wire N__41897;
    wire N__41896;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41885;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41867;
    wire N__41864;
    wire N__41861;
    wire N__41858;
    wire N__41857;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41843;
    wire N__41840;
    wire N__41837;
    wire N__41834;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41820;
    wire N__41813;
    wire N__41810;
    wire N__41809;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41799;
    wire N__41792;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41782;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41772;
    wire N__41771;
    wire N__41766;
    wire N__41763;
    wire N__41760;
    wire N__41753;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41742;
    wire N__41739;
    wire N__41736;
    wire N__41733;
    wire N__41726;
    wire N__41725;
    wire N__41722;
    wire N__41721;
    wire N__41716;
    wire N__41713;
    wire N__41708;
    wire N__41707;
    wire N__41706;
    wire N__41705;
    wire N__41700;
    wire N__41695;
    wire N__41692;
    wire N__41689;
    wire N__41684;
    wire N__41681;
    wire N__41678;
    wire N__41675;
    wire N__41672;
    wire N__41671;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41660;
    wire N__41657;
    wire N__41654;
    wire N__41651;
    wire N__41648;
    wire N__41639;
    wire N__41638;
    wire N__41635;
    wire N__41632;
    wire N__41631;
    wire N__41628;
    wire N__41625;
    wire N__41622;
    wire N__41615;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41607;
    wire N__41604;
    wire N__41599;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41589;
    wire N__41586;
    wire N__41583;
    wire N__41580;
    wire N__41573;
    wire N__41570;
    wire N__41567;
    wire N__41566;
    wire N__41565;
    wire N__41562;
    wire N__41557;
    wire N__41552;
    wire N__41549;
    wire N__41546;
    wire N__41543;
    wire N__41540;
    wire N__41537;
    wire N__41536;
    wire N__41535;
    wire N__41532;
    wire N__41529;
    wire N__41526;
    wire N__41519;
    wire N__41518;
    wire N__41517;
    wire N__41514;
    wire N__41513;
    wire N__41508;
    wire N__41505;
    wire N__41502;
    wire N__41499;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41483;
    wire N__41480;
    wire N__41479;
    wire N__41476;
    wire N__41473;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41463;
    wire N__41456;
    wire N__41453;
    wire N__41450;
    wire N__41447;
    wire N__41444;
    wire N__41441;
    wire N__41440;
    wire N__41437;
    wire N__41434;
    wire N__41431;
    wire N__41428;
    wire N__41427;
    wire N__41422;
    wire N__41419;
    wire N__41418;
    wire N__41413;
    wire N__41410;
    wire N__41405;
    wire N__41402;
    wire N__41401;
    wire N__41398;
    wire N__41397;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41381;
    wire N__41378;
    wire N__41377;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41369;
    wire N__41366;
    wire N__41361;
    wire N__41358;
    wire N__41355;
    wire N__41350;
    wire N__41345;
    wire N__41344;
    wire N__41341;
    wire N__41338;
    wire N__41337;
    wire N__41334;
    wire N__41331;
    wire N__41328;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41303;
    wire N__41302;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41283;
    wire N__41280;
    wire N__41275;
    wire N__41274;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41251;
    wire N__41250;
    wire N__41247;
    wire N__41244;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41231;
    wire N__41228;
    wire N__41225;
    wire N__41222;
    wire N__41219;
    wire N__41210;
    wire N__41209;
    wire N__41206;
    wire N__41203;
    wire N__41200;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41183;
    wire N__41180;
    wire N__41179;
    wire N__41176;
    wire N__41173;
    wire N__41170;
    wire N__41167;
    wire N__41164;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41147;
    wire N__41144;
    wire N__41141;
    wire N__41138;
    wire N__41135;
    wire N__41134;
    wire N__41133;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41121;
    wire N__41116;
    wire N__41113;
    wire N__41108;
    wire N__41105;
    wire N__41104;
    wire N__41103;
    wire N__41100;
    wire N__41097;
    wire N__41094;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41080;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41065;
    wire N__41060;
    wire N__41059;
    wire N__41056;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41048;
    wire N__41045;
    wire N__41042;
    wire N__41039;
    wire N__41036;
    wire N__41033;
    wire N__41030;
    wire N__41025;
    wire N__41018;
    wire N__41017;
    wire N__41014;
    wire N__41011;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__40999;
    wire N__40998;
    wire N__40993;
    wire N__40990;
    wire N__40985;
    wire N__40984;
    wire N__40983;
    wire N__40980;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40964;
    wire N__40957;
    wire N__40954;
    wire N__40949;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40933;
    wire N__40932;
    wire N__40929;
    wire N__40926;
    wire N__40923;
    wire N__40916;
    wire N__40913;
    wire N__40910;
    wire N__40909;
    wire N__40906;
    wire N__40903;
    wire N__40900;
    wire N__40899;
    wire N__40896;
    wire N__40893;
    wire N__40890;
    wire N__40887;
    wire N__40886;
    wire N__40883;
    wire N__40880;
    wire N__40877;
    wire N__40874;
    wire N__40869;
    wire N__40862;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40847;
    wire N__40844;
    wire N__40841;
    wire N__40838;
    wire N__40837;
    wire N__40836;
    wire N__40835;
    wire N__40832;
    wire N__40829;
    wire N__40824;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40810;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40793;
    wire N__40790;
    wire N__40787;
    wire N__40784;
    wire N__40781;
    wire N__40778;
    wire N__40775;
    wire N__40772;
    wire N__40769;
    wire N__40766;
    wire N__40763;
    wire N__40760;
    wire N__40757;
    wire N__40754;
    wire N__40751;
    wire N__40750;
    wire N__40747;
    wire N__40746;
    wire N__40739;
    wire N__40736;
    wire N__40733;
    wire N__40730;
    wire N__40727;
    wire N__40724;
    wire N__40721;
    wire N__40718;
    wire N__40715;
    wire N__40712;
    wire N__40709;
    wire N__40706;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40691;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40679;
    wire N__40678;
    wire N__40675;
    wire N__40672;
    wire N__40671;
    wire N__40670;
    wire N__40667;
    wire N__40664;
    wire N__40659;
    wire N__40656;
    wire N__40651;
    wire N__40648;
    wire N__40643;
    wire N__40640;
    wire N__40639;
    wire N__40636;
    wire N__40631;
    wire N__40628;
    wire N__40627;
    wire N__40626;
    wire N__40623;
    wire N__40622;
    wire N__40619;
    wire N__40616;
    wire N__40613;
    wire N__40610;
    wire N__40607;
    wire N__40604;
    wire N__40601;
    wire N__40598;
    wire N__40595;
    wire N__40586;
    wire N__40583;
    wire N__40582;
    wire N__40579;
    wire N__40578;
    wire N__40575;
    wire N__40572;
    wire N__40569;
    wire N__40566;
    wire N__40563;
    wire N__40556;
    wire N__40555;
    wire N__40550;
    wire N__40547;
    wire N__40544;
    wire N__40541;
    wire N__40538;
    wire N__40535;
    wire N__40532;
    wire N__40529;
    wire N__40526;
    wire N__40523;
    wire N__40520;
    wire N__40517;
    wire N__40514;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40502;
    wire N__40499;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40478;
    wire N__40475;
    wire N__40472;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40454;
    wire N__40451;
    wire N__40448;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40436;
    wire N__40433;
    wire N__40430;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40418;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40388;
    wire N__40385;
    wire N__40382;
    wire N__40379;
    wire N__40376;
    wire N__40373;
    wire N__40370;
    wire N__40367;
    wire N__40364;
    wire N__40361;
    wire N__40358;
    wire N__40357;
    wire N__40352;
    wire N__40349;
    wire N__40346;
    wire N__40343;
    wire N__40342;
    wire N__40337;
    wire N__40334;
    wire N__40331;
    wire N__40328;
    wire N__40325;
    wire N__40324;
    wire N__40323;
    wire N__40322;
    wire N__40319;
    wire N__40316;
    wire N__40313;
    wire N__40310;
    wire N__40301;
    wire N__40298;
    wire N__40297;
    wire N__40294;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40277;
    wire N__40276;
    wire N__40275;
    wire N__40272;
    wire N__40269;
    wire N__40266;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40247;
    wire N__40244;
    wire N__40241;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40220;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40196;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40169;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40154;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40142;
    wire N__40139;
    wire N__40136;
    wire N__40133;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40120;
    wire N__40119;
    wire N__40118;
    wire N__40115;
    wire N__40112;
    wire N__40109;
    wire N__40106;
    wire N__40097;
    wire N__40094;
    wire N__40093;
    wire N__40090;
    wire N__40089;
    wire N__40086;
    wire N__40083;
    wire N__40080;
    wire N__40073;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40065;
    wire N__40064;
    wire N__40061;
    wire N__40058;
    wire N__40055;
    wire N__40052;
    wire N__40043;
    wire N__40040;
    wire N__40039;
    wire N__40036;
    wire N__40035;
    wire N__40032;
    wire N__40029;
    wire N__40026;
    wire N__40019;
    wire N__40016;
    wire N__40013;
    wire N__40010;
    wire N__40009;
    wire N__40008;
    wire N__40003;
    wire N__40002;
    wire N__39999;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39985;
    wire N__39980;
    wire N__39979;
    wire N__39978;
    wire N__39975;
    wire N__39972;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39953;
    wire N__39950;
    wire N__39949;
    wire N__39946;
    wire N__39943;
    wire N__39940;
    wire N__39939;
    wire N__39938;
    wire N__39935;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39923;
    wire N__39920;
    wire N__39915;
    wire N__39908;
    wire N__39905;
    wire N__39904;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39886;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39863;
    wire N__39860;
    wire N__39857;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39847;
    wire N__39846;
    wire N__39845;
    wire N__39840;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39818;
    wire N__39815;
    wire N__39812;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39800;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39792;
    wire N__39789;
    wire N__39786;
    wire N__39783;
    wire N__39780;
    wire N__39777;
    wire N__39770;
    wire N__39769;
    wire N__39768;
    wire N__39767;
    wire N__39764;
    wire N__39761;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39747;
    wire N__39744;
    wire N__39739;
    wire N__39736;
    wire N__39731;
    wire N__39728;
    wire N__39725;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39713;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39700;
    wire N__39699;
    wire N__39696;
    wire N__39691;
    wire N__39690;
    wire N__39687;
    wire N__39684;
    wire N__39681;
    wire N__39674;
    wire N__39671;
    wire N__39668;
    wire N__39665;
    wire N__39662;
    wire N__39659;
    wire N__39656;
    wire N__39655;
    wire N__39652;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39642;
    wire N__39641;
    wire N__39636;
    wire N__39633;
    wire N__39630;
    wire N__39623;
    wire N__39620;
    wire N__39619;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39606;
    wire N__39599;
    wire N__39598;
    wire N__39597;
    wire N__39594;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39545;
    wire N__39542;
    wire N__39539;
    wire N__39536;
    wire N__39533;
    wire N__39530;
    wire N__39527;
    wire N__39524;
    wire N__39521;
    wire N__39518;
    wire N__39515;
    wire N__39512;
    wire N__39509;
    wire N__39506;
    wire N__39503;
    wire N__39500;
    wire N__39497;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39467;
    wire N__39464;
    wire N__39461;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39442;
    wire N__39439;
    wire N__39436;
    wire N__39435;
    wire N__39432;
    wire N__39427;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39359;
    wire N__39356;
    wire N__39353;
    wire N__39350;
    wire N__39347;
    wire N__39344;
    wire N__39341;
    wire N__39338;
    wire N__39335;
    wire N__39332;
    wire N__39329;
    wire N__39326;
    wire N__39323;
    wire N__39320;
    wire N__39317;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39305;
    wire N__39302;
    wire N__39299;
    wire N__39296;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39284;
    wire N__39281;
    wire N__39278;
    wire N__39275;
    wire N__39272;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39260;
    wire N__39257;
    wire N__39254;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39239;
    wire N__39236;
    wire N__39233;
    wire N__39230;
    wire N__39227;
    wire N__39224;
    wire N__39221;
    wire N__39218;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39203;
    wire N__39200;
    wire N__39199;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39184;
    wire N__39179;
    wire N__39176;
    wire N__39175;
    wire N__39174;
    wire N__39173;
    wire N__39170;
    wire N__39167;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39128;
    wire N__39125;
    wire N__39124;
    wire N__39121;
    wire N__39116;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39101;
    wire N__39100;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39088;
    wire N__39083;
    wire N__39080;
    wire N__39077;
    wire N__39074;
    wire N__39071;
    wire N__39070;
    wire N__39065;
    wire N__39062;
    wire N__39059;
    wire N__39056;
    wire N__39053;
    wire N__39050;
    wire N__39049;
    wire N__39048;
    wire N__39043;
    wire N__39040;
    wire N__39037;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39025;
    wire N__39024;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39010;
    wire N__39005;
    wire N__39002;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38977;
    wire N__38972;
    wire N__38969;
    wire N__38968;
    wire N__38963;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38948;
    wire N__38945;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38933;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38918;
    wire N__38915;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38901;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38885;
    wire N__38882;
    wire N__38879;
    wire N__38878;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38863;
    wire N__38858;
    wire N__38855;
    wire N__38854;
    wire N__38853;
    wire N__38848;
    wire N__38845;
    wire N__38842;
    wire N__38837;
    wire N__38834;
    wire N__38833;
    wire N__38830;
    wire N__38827;
    wire N__38824;
    wire N__38819;
    wire N__38816;
    wire N__38815;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38797;
    wire N__38796;
    wire N__38791;
    wire N__38788;
    wire N__38783;
    wire N__38780;
    wire N__38779;
    wire N__38774;
    wire N__38773;
    wire N__38770;
    wire N__38767;
    wire N__38764;
    wire N__38759;
    wire N__38756;
    wire N__38755;
    wire N__38752;
    wire N__38749;
    wire N__38748;
    wire N__38743;
    wire N__38740;
    wire N__38737;
    wire N__38732;
    wire N__38729;
    wire N__38728;
    wire N__38725;
    wire N__38722;
    wire N__38721;
    wire N__38716;
    wire N__38713;
    wire N__38710;
    wire N__38705;
    wire N__38702;
    wire N__38701;
    wire N__38696;
    wire N__38695;
    wire N__38692;
    wire N__38689;
    wire N__38686;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38674;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38659;
    wire N__38654;
    wire N__38651;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38640;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38624;
    wire N__38621;
    wire N__38618;
    wire N__38617;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38602;
    wire N__38597;
    wire N__38594;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38586;
    wire N__38581;
    wire N__38578;
    wire N__38575;
    wire N__38570;
    wire N__38567;
    wire N__38566;
    wire N__38563;
    wire N__38560;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38545;
    wire N__38540;
    wire N__38537;
    wire N__38536;
    wire N__38531;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38516;
    wire N__38513;
    wire N__38512;
    wire N__38509;
    wire N__38506;
    wire N__38505;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38483;
    wire N__38480;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38472;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38456;
    wire N__38453;
    wire N__38452;
    wire N__38449;
    wire N__38446;
    wire N__38445;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38429;
    wire N__38426;
    wire N__38425;
    wire N__38420;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38405;
    wire N__38404;
    wire N__38401;
    wire N__38400;
    wire N__38399;
    wire N__38396;
    wire N__38393;
    wire N__38390;
    wire N__38387;
    wire N__38384;
    wire N__38381;
    wire N__38378;
    wire N__38369;
    wire N__38366;
    wire N__38365;
    wire N__38360;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38345;
    wire N__38342;
    wire N__38339;
    wire N__38338;
    wire N__38337;
    wire N__38336;
    wire N__38333;
    wire N__38328;
    wire N__38325;
    wire N__38318;
    wire N__38315;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38301;
    wire N__38296;
    wire N__38293;
    wire N__38290;
    wire N__38285;
    wire N__38284;
    wire N__38281;
    wire N__38278;
    wire N__38275;
    wire N__38274;
    wire N__38273;
    wire N__38270;
    wire N__38267;
    wire N__38262;
    wire N__38255;
    wire N__38252;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38238;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38222;
    wire N__38219;
    wire N__38218;
    wire N__38213;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38189;
    wire N__38186;
    wire N__38183;
    wire N__38182;
    wire N__38181;
    wire N__38180;
    wire N__38179;
    wire N__38178;
    wire N__38177;
    wire N__38176;
    wire N__38175;
    wire N__38174;
    wire N__38173;
    wire N__38172;
    wire N__38171;
    wire N__38170;
    wire N__38169;
    wire N__38168;
    wire N__38167;
    wire N__38166;
    wire N__38165;
    wire N__38164;
    wire N__38163;
    wire N__38162;
    wire N__38161;
    wire N__38160;
    wire N__38159;
    wire N__38158;
    wire N__38157;
    wire N__38156;
    wire N__38155;
    wire N__38154;
    wire N__38149;
    wire N__38140;
    wire N__38131;
    wire N__38122;
    wire N__38113;
    wire N__38104;
    wire N__38095;
    wire N__38086;
    wire N__38081;
    wire N__38068;
    wire N__38063;
    wire N__38060;
    wire N__38057;
    wire N__38056;
    wire N__38055;
    wire N__38054;
    wire N__38051;
    wire N__38048;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38036;
    wire N__38033;
    wire N__38030;
    wire N__38027;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38009;
    wire N__38006;
    wire N__38003;
    wire N__38000;
    wire N__37997;
    wire N__37994;
    wire N__37991;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37979;
    wire N__37976;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37964;
    wire N__37961;
    wire N__37958;
    wire N__37955;
    wire N__37952;
    wire N__37949;
    wire N__37948;
    wire N__37947;
    wire N__37944;
    wire N__37943;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37931;
    wire N__37922;
    wire N__37919;
    wire N__37916;
    wire N__37913;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37880;
    wire N__37877;
    wire N__37874;
    wire N__37871;
    wire N__37868;
    wire N__37865;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37838;
    wire N__37835;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37808;
    wire N__37805;
    wire N__37802;
    wire N__37799;
    wire N__37796;
    wire N__37793;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37778;
    wire N__37775;
    wire N__37772;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37754;
    wire N__37751;
    wire N__37748;
    wire N__37745;
    wire N__37742;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37706;
    wire N__37703;
    wire N__37700;
    wire N__37697;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37657;
    wire N__37656;
    wire N__37653;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37628;
    wire N__37625;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37594;
    wire N__37591;
    wire N__37588;
    wire N__37585;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37571;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37561;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37505;
    wire N__37502;
    wire N__37499;
    wire N__37496;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37481;
    wire N__37478;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37436;
    wire N__37433;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37399;
    wire N__37396;
    wire N__37393;
    wire N__37390;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37327;
    wire N__37324;
    wire N__37321;
    wire N__37318;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37297;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37258;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37232;
    wire N__37229;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37210;
    wire N__37205;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37171;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37156;
    wire N__37153;
    wire N__37152;
    wire N__37149;
    wire N__37146;
    wire N__37143;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37117;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37087;
    wire N__37084;
    wire N__37081;
    wire N__37078;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36991;
    wire N__36988;
    wire N__36987;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36965;
    wire N__36964;
    wire N__36961;
    wire N__36960;
    wire N__36955;
    wire N__36952;
    wire N__36949;
    wire N__36944;
    wire N__36941;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36933;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36917;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36905;
    wire N__36902;
    wire N__36901;
    wire N__36896;
    wire N__36893;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36885;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36869;
    wire N__36868;
    wire N__36865;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36851;
    wire N__36850;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36838;
    wire N__36833;
    wire N__36832;
    wire N__36831;
    wire N__36828;
    wire N__36823;
    wire N__36818;
    wire N__36815;
    wire N__36812;
    wire N__36809;
    wire N__36806;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36781;
    wire N__36778;
    wire N__36775;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36751;
    wire N__36750;
    wire N__36749;
    wire N__36744;
    wire N__36741;
    wire N__36738;
    wire N__36733;
    wire N__36728;
    wire N__36727;
    wire N__36726;
    wire N__36725;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36685;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36675;
    wire N__36670;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36614;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36587;
    wire N__36584;
    wire N__36581;
    wire N__36578;
    wire N__36575;
    wire N__36572;
    wire N__36569;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36533;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36449;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36425;
    wire N__36422;
    wire N__36419;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36395;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36320;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36287;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36277;
    wire N__36276;
    wire N__36273;
    wire N__36268;
    wire N__36263;
    wire N__36260;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36247;
    wire N__36246;
    wire N__36243;
    wire N__36238;
    wire N__36233;
    wire N__36230;
    wire N__36229;
    wire N__36228;
    wire N__36227;
    wire N__36226;
    wire N__36225;
    wire N__36224;
    wire N__36223;
    wire N__36222;
    wire N__36221;
    wire N__36220;
    wire N__36219;
    wire N__36218;
    wire N__36217;
    wire N__36216;
    wire N__36213;
    wire N__36206;
    wire N__36197;
    wire N__36196;
    wire N__36195;
    wire N__36194;
    wire N__36193;
    wire N__36186;
    wire N__36177;
    wire N__36176;
    wire N__36175;
    wire N__36174;
    wire N__36173;
    wire N__36170;
    wire N__36169;
    wire N__36168;
    wire N__36167;
    wire N__36166;
    wire N__36165;
    wire N__36164;
    wire N__36163;
    wire N__36162;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36146;
    wire N__36141;
    wire N__36132;
    wire N__36129;
    wire N__36126;
    wire N__36117;
    wire N__36108;
    wire N__36097;
    wire N__36094;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36065;
    wire N__36062;
    wire N__36061;
    wire N__36058;
    wire N__36057;
    wire N__36054;
    wire N__36049;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36022;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36010;
    wire N__36005;
    wire N__36002;
    wire N__36001;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35989;
    wire N__35984;
    wire N__35981;
    wire N__35980;
    wire N__35977;
    wire N__35976;
    wire N__35973;
    wire N__35968;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35932;
    wire N__35929;
    wire N__35928;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35876;
    wire N__35873;
    wire N__35870;
    wire N__35867;
    wire N__35864;
    wire N__35861;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35853;
    wire N__35852;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35838;
    wire N__35831;
    wire N__35828;
    wire N__35827;
    wire N__35826;
    wire N__35823;
    wire N__35818;
    wire N__35817;
    wire N__35812;
    wire N__35809;
    wire N__35806;
    wire N__35801;
    wire N__35798;
    wire N__35797;
    wire N__35796;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35782;
    wire N__35777;
    wire N__35774;
    wire N__35773;
    wire N__35770;
    wire N__35769;
    wire N__35766;
    wire N__35763;
    wire N__35760;
    wire N__35753;
    wire N__35750;
    wire N__35747;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35693;
    wire N__35690;
    wire N__35687;
    wire N__35684;
    wire N__35681;
    wire N__35680;
    wire N__35677;
    wire N__35676;
    wire N__35673;
    wire N__35670;
    wire N__35667;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35642;
    wire N__35641;
    wire N__35638;
    wire N__35635;
    wire N__35630;
    wire N__35629;
    wire N__35628;
    wire N__35625;
    wire N__35624;
    wire N__35623;
    wire N__35618;
    wire N__35615;
    wire N__35610;
    wire N__35603;
    wire N__35602;
    wire N__35601;
    wire N__35598;
    wire N__35593;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35575;
    wire N__35574;
    wire N__35571;
    wire N__35568;
    wire N__35565;
    wire N__35558;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35546;
    wire N__35543;
    wire N__35540;
    wire N__35537;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35525;
    wire N__35522;
    wire N__35519;
    wire N__35516;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35498;
    wire N__35495;
    wire N__35492;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35444;
    wire N__35441;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35282;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35251;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35239;
    wire N__35234;
    wire N__35231;
    wire N__35228;
    wire N__35227;
    wire N__35222;
    wire N__35219;
    wire N__35218;
    wire N__35213;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35180;
    wire N__35179;
    wire N__35174;
    wire N__35171;
    wire N__35170;
    wire N__35169;
    wire N__35168;
    wire N__35165;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35135;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35111;
    wire N__35108;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35096;
    wire N__35093;
    wire N__35092;
    wire N__35091;
    wire N__35088;
    wire N__35083;
    wire N__35078;
    wire N__35075;
    wire N__35074;
    wire N__35071;
    wire N__35068;
    wire N__35067;
    wire N__35066;
    wire N__35061;
    wire N__35056;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35039;
    wire N__35038;
    wire N__35037;
    wire N__35036;
    wire N__35031;
    wire N__35026;
    wire N__35021;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35013;
    wire N__35012;
    wire N__35011;
    wire N__35008;
    wire N__35005;
    wire N__35000;
    wire N__34997;
    wire N__34988;
    wire N__34987;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34969;
    wire N__34964;
    wire N__34961;
    wire N__34958;
    wire N__34955;
    wire N__34954;
    wire N__34949;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34922;
    wire N__34921;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34909;
    wire N__34906;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34889;
    wire N__34886;
    wire N__34885;
    wire N__34882;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34871;
    wire N__34868;
    wire N__34863;
    wire N__34860;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34843;
    wire N__34842;
    wire N__34841;
    wire N__34840;
    wire N__34839;
    wire N__34838;
    wire N__34837;
    wire N__34836;
    wire N__34835;
    wire N__34834;
    wire N__34833;
    wire N__34832;
    wire N__34831;
    wire N__34830;
    wire N__34829;
    wire N__34828;
    wire N__34825;
    wire N__34818;
    wire N__34817;
    wire N__34816;
    wire N__34815;
    wire N__34810;
    wire N__34795;
    wire N__34786;
    wire N__34781;
    wire N__34780;
    wire N__34779;
    wire N__34778;
    wire N__34777;
    wire N__34776;
    wire N__34775;
    wire N__34774;
    wire N__34773;
    wire N__34772;
    wire N__34771;
    wire N__34770;
    wire N__34769;
    wire N__34768;
    wire N__34767;
    wire N__34766;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34758;
    wire N__34757;
    wire N__34756;
    wire N__34755;
    wire N__34754;
    wire N__34753;
    wire N__34752;
    wire N__34751;
    wire N__34750;
    wire N__34749;
    wire N__34748;
    wire N__34747;
    wire N__34746;
    wire N__34743;
    wire N__34742;
    wire N__34741;
    wire N__34740;
    wire N__34739;
    wire N__34738;
    wire N__34737;
    wire N__34736;
    wire N__34735;
    wire N__34734;
    wire N__34733;
    wire N__34732;
    wire N__34723;
    wire N__34712;
    wire N__34711;
    wire N__34710;
    wire N__34709;
    wire N__34704;
    wire N__34691;
    wire N__34686;
    wire N__34685;
    wire N__34684;
    wire N__34683;
    wire N__34680;
    wire N__34679;
    wire N__34674;
    wire N__34673;
    wire N__34672;
    wire N__34671;
    wire N__34670;
    wire N__34669;
    wire N__34668;
    wire N__34667;
    wire N__34666;
    wire N__34663;
    wire N__34660;
    wire N__34647;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34623;
    wire N__34620;
    wire N__34615;
    wire N__34614;
    wire N__34613;
    wire N__34612;
    wire N__34611;
    wire N__34610;
    wire N__34609;
    wire N__34608;
    wire N__34607;
    wire N__34606;
    wire N__34605;
    wire N__34604;
    wire N__34603;
    wire N__34602;
    wire N__34601;
    wire N__34600;
    wire N__34599;
    wire N__34590;
    wire N__34585;
    wire N__34582;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34568;
    wire N__34557;
    wire N__34554;
    wire N__34551;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34525;
    wire N__34520;
    wire N__34517;
    wire N__34512;
    wire N__34507;
    wire N__34504;
    wire N__34491;
    wire N__34486;
    wire N__34475;
    wire N__34472;
    wire N__34469;
    wire N__34464;
    wire N__34459;
    wire N__34452;
    wire N__34435;
    wire N__34412;
    wire N__34409;
    wire N__34408;
    wire N__34405;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34390;
    wire N__34385;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34365;
    wire N__34364;
    wire N__34361;
    wire N__34356;
    wire N__34353;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34333;
    wire N__34332;
    wire N__34331;
    wire N__34330;
    wire N__34329;
    wire N__34328;
    wire N__34327;
    wire N__34326;
    wire N__34325;
    wire N__34324;
    wire N__34323;
    wire N__34322;
    wire N__34321;
    wire N__34320;
    wire N__34319;
    wire N__34318;
    wire N__34317;
    wire N__34316;
    wire N__34313;
    wire N__34312;
    wire N__34311;
    wire N__34310;
    wire N__34309;
    wire N__34302;
    wire N__34293;
    wire N__34284;
    wire N__34281;
    wire N__34280;
    wire N__34277;
    wire N__34276;
    wire N__34267;
    wire N__34264;
    wire N__34263;
    wire N__34262;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34254;
    wire N__34247;
    wire N__34238;
    wire N__34237;
    wire N__34236;
    wire N__34235;
    wire N__34234;
    wire N__34233;
    wire N__34232;
    wire N__34231;
    wire N__34230;
    wire N__34229;
    wire N__34228;
    wire N__34227;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34217;
    wire N__34212;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34202;
    wire N__34197;
    wire N__34194;
    wire N__34189;
    wire N__34180;
    wire N__34171;
    wire N__34162;
    wire N__34159;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34145;
    wire N__34142;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34121;
    wire N__34118;
    wire N__34115;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34099;
    wire N__34094;
    wire N__34089;
    wire N__34076;
    wire N__34075;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34054;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34039;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34019;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34001;
    wire N__33998;
    wire N__33997;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33955;
    wire N__33954;
    wire N__33951;
    wire N__33946;
    wire N__33941;
    wire N__33938;
    wire N__33937;
    wire N__33936;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33901;
    wire N__33900;
    wire N__33897;
    wire N__33894;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33878;
    wire N__33875;
    wire N__33874;
    wire N__33871;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33860;
    wire N__33857;
    wire N__33852;
    wire N__33849;
    wire N__33842;
    wire N__33839;
    wire N__33838;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33761;
    wire N__33758;
    wire N__33755;
    wire N__33752;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33740;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33546;
    wire N__33545;
    wire N__33540;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33506;
    wire N__33503;
    wire N__33500;
    wire N__33497;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33469;
    wire N__33468;
    wire N__33461;
    wire N__33458;
    wire N__33457;
    wire N__33454;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33437;
    wire N__33434;
    wire N__33431;
    wire N__33428;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33416;
    wire N__33413;
    wire N__33412;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33400;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33355;
    wire N__33354;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33338;
    wire N__33335;
    wire N__33334;
    wire N__33329;
    wire N__33326;
    wire N__33325;
    wire N__33324;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33308;
    wire N__33305;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33293;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33281;
    wire N__33278;
    wire N__33277;
    wire N__33276;
    wire N__33273;
    wire N__33268;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33242;
    wire N__33239;
    wire N__33238;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33217;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33200;
    wire N__33197;
    wire N__33196;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33184;
    wire N__33179;
    wire N__33176;
    wire N__33175;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33163;
    wire N__33158;
    wire N__33155;
    wire N__33154;
    wire N__33153;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33137;
    wire N__33134;
    wire N__33133;
    wire N__33132;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33116;
    wire N__33113;
    wire N__33112;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33079;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33066;
    wire N__33059;
    wire N__33056;
    wire N__33055;
    wire N__33052;
    wire N__33049;
    wire N__33046;
    wire N__33041;
    wire N__33038;
    wire N__33037;
    wire N__33036;
    wire N__33033;
    wire N__33028;
    wire N__33023;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32985;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32969;
    wire N__32966;
    wire N__32965;
    wire N__32964;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32948;
    wire N__32945;
    wire N__32944;
    wire N__32941;
    wire N__32940;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32924;
    wire N__32921;
    wire N__32920;
    wire N__32919;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32903;
    wire N__32900;
    wire N__32899;
    wire N__32898;
    wire N__32893;
    wire N__32890;
    wire N__32887;
    wire N__32882;
    wire N__32879;
    wire N__32878;
    wire N__32877;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32851;
    wire N__32848;
    wire N__32845;
    wire N__32840;
    wire N__32837;
    wire N__32836;
    wire N__32833;
    wire N__32830;
    wire N__32825;
    wire N__32822;
    wire N__32821;
    wire N__32818;
    wire N__32815;
    wire N__32810;
    wire N__32807;
    wire N__32806;
    wire N__32803;
    wire N__32800;
    wire N__32795;
    wire N__32792;
    wire N__32791;
    wire N__32788;
    wire N__32785;
    wire N__32780;
    wire N__32777;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32765;
    wire N__32762;
    wire N__32761;
    wire N__32758;
    wire N__32755;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32737;
    wire N__32734;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32717;
    wire N__32714;
    wire N__32713;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32700;
    wire N__32697;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32680;
    wire N__32677;
    wire N__32674;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32651;
    wire N__32648;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32636;
    wire N__32633;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32621;
    wire N__32618;
    wire N__32617;
    wire N__32614;
    wire N__32611;
    wire N__32606;
    wire N__32603;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32591;
    wire N__32588;
    wire N__32587;
    wire N__32584;
    wire N__32581;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32536;
    wire N__32533;
    wire N__32530;
    wire N__32527;
    wire N__32522;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32510;
    wire N__32507;
    wire N__32506;
    wire N__32505;
    wire N__32504;
    wire N__32503;
    wire N__32502;
    wire N__32501;
    wire N__32498;
    wire N__32491;
    wire N__32484;
    wire N__32477;
    wire N__32474;
    wire N__32471;
    wire N__32470;
    wire N__32469;
    wire N__32468;
    wire N__32467;
    wire N__32466;
    wire N__32465;
    wire N__32464;
    wire N__32463;
    wire N__32462;
    wire N__32461;
    wire N__32460;
    wire N__32459;
    wire N__32458;
    wire N__32457;
    wire N__32440;
    wire N__32425;
    wire N__32424;
    wire N__32423;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32411;
    wire N__32410;
    wire N__32409;
    wire N__32408;
    wire N__32407;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32396;
    wire N__32395;
    wire N__32394;
    wire N__32393;
    wire N__32392;
    wire N__32391;
    wire N__32390;
    wire N__32389;
    wire N__32386;
    wire N__32381;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32367;
    wire N__32364;
    wire N__32347;
    wire N__32344;
    wire N__32339;
    wire N__32336;
    wire N__32333;
    wire N__32330;
    wire N__32321;
    wire N__32318;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32288;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32257;
    wire N__32254;
    wire N__32253;
    wire N__32250;
    wire N__32247;
    wire N__32244;
    wire N__32243;
    wire N__32240;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32219;
    wire N__32216;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32186;
    wire N__32183;
    wire N__32180;
    wire N__32179;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32168;
    wire N__32165;
    wire N__32160;
    wire N__32157;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32065;
    wire N__32062;
    wire N__32059;
    wire N__32054;
    wire N__32051;
    wire N__32048;
    wire N__32045;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32012;
    wire N__32009;
    wire N__32006;
    wire N__32003;
    wire N__32000;
    wire N__31997;
    wire N__31994;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31925;
    wire N__31922;
    wire N__31919;
    wire N__31916;
    wire N__31913;
    wire N__31910;
    wire N__31907;
    wire N__31904;
    wire N__31901;
    wire N__31898;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31883;
    wire N__31880;
    wire N__31877;
    wire N__31874;
    wire N__31871;
    wire N__31868;
    wire N__31865;
    wire N__31862;
    wire N__31859;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31847;
    wire N__31844;
    wire N__31841;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31768;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31748;
    wire N__31745;
    wire N__31742;
    wire N__31739;
    wire N__31736;
    wire N__31733;
    wire N__31730;
    wire N__31727;
    wire N__31724;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31691;
    wire N__31688;
    wire N__31685;
    wire N__31682;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31634;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31615;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31604;
    wire N__31599;
    wire N__31596;
    wire N__31595;
    wire N__31592;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31574;
    wire N__31573;
    wire N__31570;
    wire N__31569;
    wire N__31566;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31541;
    wire N__31540;
    wire N__31539;
    wire N__31538;
    wire N__31537;
    wire N__31536;
    wire N__31535;
    wire N__31534;
    wire N__31533;
    wire N__31532;
    wire N__31531;
    wire N__31530;
    wire N__31529;
    wire N__31528;
    wire N__31527;
    wire N__31526;
    wire N__31525;
    wire N__31524;
    wire N__31523;
    wire N__31522;
    wire N__31521;
    wire N__31520;
    wire N__31519;
    wire N__31516;
    wire N__31515;
    wire N__31514;
    wire N__31513;
    wire N__31512;
    wire N__31511;
    wire N__31510;
    wire N__31509;
    wire N__31508;
    wire N__31499;
    wire N__31492;
    wire N__31483;
    wire N__31476;
    wire N__31467;
    wire N__31458;
    wire N__31455;
    wire N__31446;
    wire N__31437;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31418;
    wire N__31411;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31391;
    wire N__31390;
    wire N__31389;
    wire N__31386;
    wire N__31381;
    wire N__31380;
    wire N__31379;
    wire N__31376;
    wire N__31373;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31355;
    wire N__31352;
    wire N__31351;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31327;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31312;
    wire N__31307;
    wire N__31304;
    wire N__31303;
    wire N__31298;
    wire N__31295;
    wire N__31294;
    wire N__31291;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31280;
    wire N__31277;
    wire N__31272;
    wire N__31269;
    wire N__31264;
    wire N__31259;
    wire N__31256;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31244;
    wire N__31243;
    wire N__31242;
    wire N__31241;
    wire N__31238;
    wire N__31231;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31205;
    wire N__31202;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31174;
    wire N__31173;
    wire N__31170;
    wire N__31165;
    wire N__31164;
    wire N__31159;
    wire N__31156;
    wire N__31153;
    wire N__31150;
    wire N__31145;
    wire N__31144;
    wire N__31139;
    wire N__31136;
    wire N__31135;
    wire N__31132;
    wire N__31129;
    wire N__31124;
    wire N__31121;
    wire N__31120;
    wire N__31119;
    wire N__31116;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31088;
    wire N__31087;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31058;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31037;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30977;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30944;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30917;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30857;
    wire N__30854;
    wire N__30853;
    wire N__30848;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30831;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30815;
    wire N__30814;
    wire N__30811;
    wire N__30808;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30800;
    wire N__30797;
    wire N__30792;
    wire N__30787;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30725;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30641;
    wire N__30638;
    wire N__30635;
    wire N__30632;
    wire N__30629;
    wire N__30626;
    wire N__30623;
    wire N__30620;
    wire N__30617;
    wire N__30614;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30569;
    wire N__30566;
    wire N__30563;
    wire N__30560;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30545;
    wire N__30542;
    wire N__30539;
    wire N__30536;
    wire N__30533;
    wire N__30530;
    wire N__30529;
    wire N__30526;
    wire N__30525;
    wire N__30522;
    wire N__30521;
    wire N__30520;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30507;
    wire N__30504;
    wire N__30503;
    wire N__30502;
    wire N__30501;
    wire N__30500;
    wire N__30499;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30487;
    wire N__30482;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30465;
    wire N__30462;
    wire N__30457;
    wire N__30454;
    wire N__30449;
    wire N__30440;
    wire N__30437;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30395;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30236;
    wire N__30233;
    wire N__30230;
    wire N__30227;
    wire N__30224;
    wire N__30221;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30200;
    wire N__30197;
    wire N__30194;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30005;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29909;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29893;
    wire N__29888;
    wire N__29887;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29873;
    wire N__29870;
    wire N__29869;
    wire N__29864;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29842;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29830;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29818;
    wire N__29817;
    wire N__29814;
    wire N__29809;
    wire N__29804;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29792;
    wire N__29789;
    wire N__29788;
    wire N__29785;
    wire N__29782;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29767;
    wire N__29766;
    wire N__29765;
    wire N__29764;
    wire N__29763;
    wire N__29762;
    wire N__29761;
    wire N__29760;
    wire N__29759;
    wire N__29758;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29716;
    wire N__29713;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29693;
    wire N__29690;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29680;
    wire N__29679;
    wire N__29678;
    wire N__29675;
    wire N__29668;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29645;
    wire N__29642;
    wire N__29641;
    wire N__29640;
    wire N__29637;
    wire N__29632;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29615;
    wire N__29612;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29593;
    wire N__29592;
    wire N__29589;
    wire N__29584;
    wire N__29579;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29567;
    wire N__29564;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29531;
    wire N__29528;
    wire N__29527;
    wire N__29522;
    wire N__29519;
    wire N__29518;
    wire N__29517;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29501;
    wire N__29500;
    wire N__29497;
    wire N__29496;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29480;
    wire N__29479;
    wire N__29476;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29458;
    wire N__29455;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29441;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29423;
    wire N__29420;
    wire N__29419;
    wire N__29416;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29377;
    wire N__29372;
    wire N__29369;
    wire N__29368;
    wire N__29363;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29348;
    wire N__29347;
    wire N__29344;
    wire N__29339;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29308;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29293;
    wire N__29288;
    wire N__29287;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29261;
    wire N__29258;
    wire N__29249;
    wire N__29246;
    wire N__29245;
    wire N__29240;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29217;
    wire N__29212;
    wire N__29209;
    wire N__29206;
    wire N__29201;
    wire N__29198;
    wire N__29197;
    wire N__29194;
    wire N__29191;
    wire N__29190;
    wire N__29189;
    wire N__29184;
    wire N__29179;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29162;
    wire N__29161;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29132;
    wire N__29131;
    wire N__29126;
    wire N__29123;
    wire N__29122;
    wire N__29119;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29107;
    wire N__29106;
    wire N__29105;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29085;
    wire N__29082;
    wire N__29075;
    wire N__29074;
    wire N__29071;
    wire N__29070;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29054;
    wire N__29053;
    wire N__29048;
    wire N__29045;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29026;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29011;
    wire N__29006;
    wire N__29005;
    wire N__29002;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28994;
    wire N__28991;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28977;
    wire N__28970;
    wire N__28967;
    wire N__28966;
    wire N__28963;
    wire N__28962;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28946;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28928;
    wire N__28925;
    wire N__28922;
    wire N__28919;
    wire N__28916;
    wire N__28907;
    wire N__28906;
    wire N__28903;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28886;
    wire N__28885;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28844;
    wire N__28841;
    wire N__28840;
    wire N__28837;
    wire N__28834;
    wire N__28829;
    wire N__28828;
    wire N__28827;
    wire N__28824;
    wire N__28819;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28784;
    wire N__28783;
    wire N__28782;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28770;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28740;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28728;
    wire N__28721;
    wire N__28720;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28705;
    wire N__28700;
    wire N__28699;
    wire N__28698;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28682;
    wire N__28681;
    wire N__28680;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28647;
    wire N__28640;
    wire N__28639;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28622;
    wire N__28619;
    wire N__28618;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28607;
    wire N__28604;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28541;
    wire N__28538;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28493;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28468;
    wire N__28467;
    wire N__28466;
    wire N__28465;
    wire N__28464;
    wire N__28457;
    wire N__28454;
    wire N__28453;
    wire N__28452;
    wire N__28451;
    wire N__28450;
    wire N__28445;
    wire N__28442;
    wire N__28439;
    wire N__28430;
    wire N__28427;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28244;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28172;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28145;
    wire N__28142;
    wire N__28141;
    wire N__28138;
    wire N__28135;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28061;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28049;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28028;
    wire N__28025;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27992;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27913;
    wire N__27910;
    wire N__27907;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27893;
    wire N__27892;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27866;
    wire N__27863;
    wire N__27860;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27836;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27826;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27767;
    wire N__27764;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27686;
    wire N__27683;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27673;
    wire N__27670;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27653;
    wire N__27650;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27596;
    wire N__27593;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27550;
    wire N__27547;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27530;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27505;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27446;
    wire N__27443;
    wire N__27440;
    wire N__27437;
    wire N__27434;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27409;
    wire N__27408;
    wire N__27405;
    wire N__27400;
    wire N__27397;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27332;
    wire N__27329;
    wire N__27328;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27295;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27271;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27247;
    wire N__27244;
    wire N__27241;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27161;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27025;
    wire N__27022;
    wire N__27019;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26992;
    wire N__26989;
    wire N__26986;
    wire N__26981;
    wire N__26978;
    wire N__26975;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26945;
    wire N__26942;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26923;
    wire N__26922;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26906;
    wire N__26905;
    wire N__26902;
    wire N__26897;
    wire N__26894;
    wire N__26893;
    wire N__26890;
    wire N__26885;
    wire N__26884;
    wire N__26881;
    wire N__26878;
    wire N__26875;
    wire N__26870;
    wire N__26869;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26831;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26810;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26789;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26735;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26723;
    wire N__26722;
    wire N__26719;
    wire N__26718;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26706;
    wire N__26703;
    wire N__26696;
    wire N__26693;
    wire N__26692;
    wire N__26691;
    wire N__26690;
    wire N__26687;
    wire N__26682;
    wire N__26679;
    wire N__26672;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26660;
    wire N__26659;
    wire N__26654;
    wire N__26651;
    wire N__26650;
    wire N__26649;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26633;
    wire N__26630;
    wire N__26629;
    wire N__26628;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26612;
    wire N__26609;
    wire N__26608;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26596;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26584;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26527;
    wire N__26522;
    wire N__26519;
    wire N__26518;
    wire N__26515;
    wire N__26510;
    wire N__26507;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26492;
    wire N__26491;
    wire N__26486;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26471;
    wire N__26470;
    wire N__26467;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26446;
    wire N__26443;
    wire N__26440;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26425;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26413;
    wire N__26408;
    wire N__26407;
    wire N__26406;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26381;
    wire N__26380;
    wire N__26379;
    wire N__26376;
    wire N__26373;
    wire N__26372;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26353;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26337;
    wire N__26330;
    wire N__26329;
    wire N__26328;
    wire N__26327;
    wire N__26324;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26306;
    wire N__26303;
    wire N__26302;
    wire N__26299;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26289;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26269;
    wire N__26268;
    wire N__26265;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26218;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26189;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26158;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26146;
    wire N__26141;
    wire N__26138;
    wire N__26137;
    wire N__26136;
    wire N__26133;
    wire N__26128;
    wire N__26123;
    wire N__26120;
    wire N__26119;
    wire N__26118;
    wire N__26115;
    wire N__26110;
    wire N__26105;
    wire N__26102;
    wire N__26101;
    wire N__26100;
    wire N__26097;
    wire N__26094;
    wire N__26089;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26074;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25988;
    wire N__25985;
    wire N__25984;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25967;
    wire N__25964;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25952;
    wire N__25949;
    wire N__25948;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25891;
    wire N__25890;
    wire N__25887;
    wire N__25884;
    wire N__25881;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25867;
    wire N__25866;
    wire N__25863;
    wire N__25860;
    wire N__25857;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25843;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25819;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25795;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25771;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25747;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25723;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25699;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25682;
    wire N__25679;
    wire N__25678;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25654;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25630;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25606;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25582;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25558;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25534;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25510;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25493;
    wire N__25490;
    wire N__25489;
    wire N__25486;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25469;
    wire N__25468;
    wire N__25465;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25441;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25417;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25393;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25369;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25345;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25321;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25297;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25280;
    wire N__25277;
    wire N__25276;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25241;
    wire N__25238;
    wire N__25237;
    wire N__25232;
    wire N__25229;
    wire N__25228;
    wire N__25225;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25207;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25186;
    wire N__25185;
    wire N__25182;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25149;
    wire N__25148;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25129;
    wire N__25124;
    wire N__25121;
    wire N__25120;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25108;
    wire N__25103;
    wire N__25102;
    wire N__25101;
    wire N__25100;
    wire N__25099;
    wire N__25098;
    wire N__25097;
    wire N__25096;
    wire N__25095;
    wire N__25092;
    wire N__25083;
    wire N__25082;
    wire N__25081;
    wire N__25080;
    wire N__25079;
    wire N__25078;
    wire N__25077;
    wire N__25076;
    wire N__25075;
    wire N__25074;
    wire N__25073;
    wire N__25072;
    wire N__25071;
    wire N__25070;
    wire N__25069;
    wire N__25068;
    wire N__25067;
    wire N__25066;
    wire N__25065;
    wire N__25064;
    wire N__25063;
    wire N__25054;
    wire N__25049;
    wire N__25040;
    wire N__25031;
    wire N__25022;
    wire N__25013;
    wire N__25004;
    wire N__24997;
    wire N__24988;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24976;
    wire N__24975;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24950;
    wire N__24949;
    wire N__24946;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24853;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24833;
    wire N__24830;
    wire N__24829;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24806;
    wire N__24803;
    wire N__24802;
    wire N__24801;
    wire N__24800;
    wire N__24799;
    wire N__24798;
    wire N__24797;
    wire N__24796;
    wire N__24795;
    wire N__24794;
    wire N__24785;
    wire N__24780;
    wire N__24771;
    wire N__24766;
    wire N__24761;
    wire N__24758;
    wire N__24757;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24709;
    wire N__24706;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24696;
    wire N__24689;
    wire N__24686;
    wire N__24685;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24665;
    wire N__24662;
    wire N__24661;
    wire N__24658;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24641;
    wire N__24638;
    wire N__24637;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24617;
    wire N__24614;
    wire N__24613;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24593;
    wire N__24590;
    wire N__24589;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24569;
    wire N__24566;
    wire N__24565;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24238;
    wire N__24235;
    wire N__24232;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24165;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24146;
    wire N__24143;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24135;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24109;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24083;
    wire N__24080;
    wire N__24077;
    wire N__24076;
    wire N__24075;
    wire N__24074;
    wire N__24073;
    wire N__24072;
    wire N__24071;
    wire N__24070;
    wire N__24069;
    wire N__24066;
    wire N__24049;
    wire N__24044;
    wire N__24043;
    wire N__24042;
    wire N__24041;
    wire N__24040;
    wire N__24039;
    wire N__24038;
    wire N__24035;
    wire N__24034;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24000;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23983;
    wire N__23980;
    wire N__23977;
    wire N__23976;
    wire N__23973;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23878;
    wire N__23877;
    wire N__23874;
    wire N__23873;
    wire N__23872;
    wire N__23871;
    wire N__23870;
    wire N__23869;
    wire N__23868;
    wire N__23867;
    wire N__23866;
    wire N__23865;
    wire N__23860;
    wire N__23857;
    wire N__23852;
    wire N__23851;
    wire N__23850;
    wire N__23849;
    wire N__23848;
    wire N__23847;
    wire N__23846;
    wire N__23845;
    wire N__23844;
    wire N__23843;
    wire N__23842;
    wire N__23839;
    wire N__23838;
    wire N__23837;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23820;
    wire N__23813;
    wire N__23810;
    wire N__23805;
    wire N__23804;
    wire N__23803;
    wire N__23802;
    wire N__23801;
    wire N__23800;
    wire N__23785;
    wire N__23782;
    wire N__23775;
    wire N__23766;
    wire N__23763;
    wire N__23762;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23743;
    wire N__23738;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23718;
    wire N__23705;
    wire N__23704;
    wire N__23703;
    wire N__23702;
    wire N__23701;
    wire N__23700;
    wire N__23699;
    wire N__23698;
    wire N__23691;
    wire N__23690;
    wire N__23689;
    wire N__23688;
    wire N__23687;
    wire N__23686;
    wire N__23685;
    wire N__23684;
    wire N__23683;
    wire N__23682;
    wire N__23679;
    wire N__23678;
    wire N__23675;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23661;
    wire N__23660;
    wire N__23659;
    wire N__23658;
    wire N__23657;
    wire N__23656;
    wire N__23655;
    wire N__23654;
    wire N__23653;
    wire N__23652;
    wire N__23651;
    wire N__23648;
    wire N__23647;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23630;
    wire N__23625;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23593;
    wire N__23584;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23563;
    wire N__23556;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23521;
    wire N__23520;
    wire N__23519;
    wire N__23518;
    wire N__23517;
    wire N__23516;
    wire N__23515;
    wire N__23514;
    wire N__23513;
    wire N__23512;
    wire N__23511;
    wire N__23510;
    wire N__23509;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23505;
    wire N__23504;
    wire N__23503;
    wire N__23502;
    wire N__23501;
    wire N__23500;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23484;
    wire N__23477;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23461;
    wire N__23460;
    wire N__23459;
    wire N__23456;
    wire N__23455;
    wire N__23454;
    wire N__23453;
    wire N__23452;
    wire N__23447;
    wire N__23440;
    wire N__23435;
    wire N__23420;
    wire N__23415;
    wire N__23408;
    wire N__23401;
    wire N__23394;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23372;
    wire N__23367;
    wire N__23364;
    wire N__23351;
    wire N__23350;
    wire N__23349;
    wire N__23346;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23293;
    wire N__23290;
    wire N__23289;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23264;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23179;
    wire N__23176;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23141;
    wire N__23138;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23116;
    wire N__23113;
    wire N__23112;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23087;
    wire N__23086;
    wire N__23083;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23065;
    wire N__23064;
    wire N__23061;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23043;
    wire N__23036;
    wire N__23035;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23010;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22985;
    wire N__22984;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22955;
    wire N__22952;
    wire N__22947;
    wire N__22944;
    wire N__22937;
    wire N__22936;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22911;
    wire N__22908;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22886;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22867;
    wire N__22864;
    wire N__22863;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22838;
    wire N__22837;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22819;
    wire N__22818;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22796;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22765;
    wire N__22764;
    wire N__22761;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22743;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22705;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22694;
    wire N__22691;
    wire N__22686;
    wire N__22683;
    wire N__22676;
    wire N__22675;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22660;
    wire N__22657;
    wire N__22656;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22631;
    wire N__22628;
    wire N__22627;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22612;
    wire N__22609;
    wire N__22608;
    wire N__22605;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22587;
    wire N__22584;
    wire N__22577;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22546;
    wire N__22543;
    wire N__22542;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22517;
    wire N__22514;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22495;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22463;
    wire N__22462;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22435;
    wire N__22432;
    wire N__22431;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22408;
    wire N__22403;
    wire N__22402;
    wire N__22399;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22371;
    wire N__22368;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22350;
    wire N__22343;
    wire N__22340;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22309;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22280;
    wire N__22277;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22256;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22238;
    wire N__22235;
    wire N__22234;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22199;
    wire N__22196;
    wire N__22195;
    wire N__22194;
    wire N__22191;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22161;
    wire N__22154;
    wire N__22153;
    wire N__22150;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22105;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22081;
    wire N__22078;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22061;
    wire N__22060;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22002;
    wire N__21999;
    wire N__21992;
    wire N__21991;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21979;
    wire N__21978;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21952;
    wire N__21947;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21919;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21888;
    wire N__21885;
    wire N__21878;
    wire N__21875;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21856;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21848;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21835;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21811;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21793;
    wire N__21790;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21739;
    wire N__21736;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21721;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21695;
    wire N__21692;
    wire N__21691;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21655;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21638;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21611;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21594;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21577;
    wire N__21576;
    wire N__21573;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21544;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21487;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21454;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21442;
    wire N__21441;
    wire N__21438;
    wire N__21435;
    wire N__21432;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21397;
    wire N__21394;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21334;
    wire N__21329;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21311;
    wire N__21310;
    wire N__21307;
    wire N__21306;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21281;
    wire N__21278;
    wire N__21277;
    wire N__21276;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21251;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21211;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21064;
    wire N__21063;
    wire N__21062;
    wire N__21061;
    wire N__21060;
    wire N__21059;
    wire N__21056;
    wire N__21051;
    wire N__21044;
    wire N__21041;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20884;
    wire N__20881;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20785;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20722;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20705;
    wire N__20702;
    wire N__20701;
    wire N__20698;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20681;
    wire N__20680;
    wire N__20677;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20653;
    wire N__20652;
    wire N__20651;
    wire N__20650;
    wire N__20647;
    wire N__20640;
    wire N__20639;
    wire N__20638;
    wire N__20637;
    wire N__20632;
    wire N__20629;
    wire N__20622;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20601;
    wire N__20598;
    wire N__20593;
    wire N__20588;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20573;
    wire N__20570;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20555;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20540;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20530;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20167;
    wire N__20166;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19492;
    wire N__19491;
    wire N__19490;
    wire N__19489;
    wire N__19488;
    wire N__19487;
    wire N__19486;
    wire N__19485;
    wire N__19484;
    wire N__19483;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19443;
    wire N__19436;
    wire N__19427;
    wire N__19422;
    wire N__19417;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire bfn_1_11_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire bfn_1_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire bfn_1_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire bfn_1_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire bfn_1_15_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire bfn_1_16_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_98_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_96_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.N_94 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.N_161 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_1_24_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_1_25_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire bfn_1_26_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_43_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire rgb_drv_RNOZ0;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_44_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.N_77 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.N_159 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire bfn_3_23_0_;
    wire \pwm_generator_inst.un19_threshold_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_7 ;
    wire \pwm_generator_inst.un19_threshold_axb_8 ;
    wire bfn_3_24_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_axb_3 ;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire pwm_duty_input_9;
    wire pwm_duty_input_8;
    wire pwm_duty_input_6;
    wire pwm_duty_input_7;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un19_threshold_axb_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire bfn_4_17_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire bfn_4_18_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire bfn_4_19_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire bfn_4_20_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ;
    wire \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ;
    wire pwm_duty_input_3;
    wire pwm_duty_input_4;
    wire pwm_duty_input_5;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.N_16 ;
    wire \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ;
    wire \pwm_generator_inst.N_17_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un19_threshold_axb_0 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_46 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.N_47 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire \pwm_generator_inst.threshold_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_5_23_0_;
    wire \pwm_generator_inst.un14_counter_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.threshold_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.threshold_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.threshold_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.threshold_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.un14_counter_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.un14_counter_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.un14_counter_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_5_24_0_;
    wire \pwm_generator_inst.threshold_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire N_38_i_i;
    wire \pwm_generator_inst.un1_counterlto9_2_cascade_ ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire bfn_5_26_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire bfn_5_27_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire bfn_7_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_7_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_7_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_7_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \phase_controller_inst2.start_timer_tr_RNO_0_0 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ;
    wire il_max_comp2_c;
    wire \delay_measurement_inst.delay_tr_timer.N_201_i ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_8_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_8_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_8_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_8_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire bfn_8_11_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire bfn_8_12_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_8_13_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_8_14_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst2.state_RNIG7JFZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_200_i ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire s3_phy_c;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire s4_phy_c;
    wire GB_BUFFER_clock_output_0_THRU_CO;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21_cascade_;
    wire elapsed_time_ns_1_RNI5FOBB_0_18_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14_cascade_;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_9_12_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_9_13_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire bfn_9_14_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_9_15_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire bfn_9_16_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_16 ;
    wire bfn_9_17_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_16 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_17 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_18 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_19 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_20 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_23 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_24 ;
    wire bfn_9_18_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_24 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_25 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_26 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_27 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_28 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_30 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire bfn_9_26_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ;
    wire bfn_9_27_0_;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire bfn_9_28_0_;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire il_min_comp1_c;
    wire il_min_comp1_D1;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire elapsed_time_ns_1_RNIU7OBB_0_11_cascade_;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10_cascade_;
    wire elapsed_time_ns_1_RNILK91B_0_9_cascade_;
    wire elapsed_time_ns_1_RNIU8PBB_0_20_cascade_;
    wire elapsed_time_ns_1_RNI2COBB_0_15_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_start_g ;
    wire \current_shift_inst.control_input_axb_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire bfn_10_26_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ;
    wire bfn_10_27_0_;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire bfn_10_28_0_;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_11_8_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_11_9_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire bfn_11_10_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire elapsed_time_ns_1_RNI5GPBB_0_27_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire elapsed_time_ns_1_RNI4FPBB_0_26_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire T45_c;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.N_1269_i ;
    wire \current_shift_inst.control_input_1 ;
    wire bfn_11_15_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_11_16_0_;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ;
    wire \current_shift_inst.control_input_cry_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ;
    wire \current_shift_inst.control_input_cry_14 ;
    wire \current_shift_inst.control_input_cry_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ;
    wire bfn_11_17_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ;
    wire \current_shift_inst.control_input_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ;
    wire \current_shift_inst.control_input_cry_17 ;
    wire \current_shift_inst.control_input_axb_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ;
    wire \current_shift_inst.control_input_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ;
    wire \current_shift_inst.control_input_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ;
    wire \current_shift_inst.control_input_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ;
    wire \current_shift_inst.control_input_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ;
    wire \current_shift_inst.control_input_cry_22 ;
    wire \current_shift_inst.control_input_cry_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ;
    wire bfn_11_18_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ;
    wire \current_shift_inst.control_input_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ;
    wire \current_shift_inst.control_input_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ;
    wire \current_shift_inst.control_input_cry_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ;
    wire \current_shift_inst.control_input_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ;
    wire \current_shift_inst.control_input_cry_28 ;
    wire \current_shift_inst.control_input_cry_29 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.control_input_axb_27 ;
    wire \current_shift_inst.control_input_axb_18 ;
    wire \current_shift_inst.control_input_axb_17 ;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire N_19_1;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire il_max_comp1_c;
    wire il_max_comp1_D1;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire bfn_12_7_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_12_8_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_12_9_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_12_10_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire elapsed_time_ns_1_RNI4EOBB_0_17_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_ ;
    wire state_ns_i_a3_1;
    wire start_stop_c;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire bfn_12_16_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ;
    wire \current_shift_inst.un38_control_input_0_s0_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_8 ;
    wire bfn_12_17_0_;
    wire \current_shift_inst.un38_control_input_0_s0_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire bfn_12_18_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire bfn_12_19_0_;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_28 ;
    wire \current_shift_inst.control_input_axb_29 ;
    wire \pll_inst.red_c_i ;
    wire delay_hc_input_c_g;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire elapsed_time_ns_1_RNI2DPBB_0_24_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.state_RNI7NN7Z0Z_0 ;
    wire \phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ;
    wire \current_shift_inst.un38_control_input_0_s0_10 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ;
    wire \current_shift_inst.un38_control_input_0_s0_14 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.un38_control_input_0_s0_15 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.un38_control_input_0_s0_16 ;
    wire \current_shift_inst.control_input_axb_13 ;
    wire \current_shift_inst.un38_control_input_0_s0_17 ;
    wire \current_shift_inst.control_input_axb_14 ;
    wire \current_shift_inst.un38_control_input_0_s0_18 ;
    wire \current_shift_inst.control_input_axb_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ;
    wire \current_shift_inst.un38_control_input_0_s0_19 ;
    wire \current_shift_inst.control_input_axb_16 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.control_input_axb_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.control_input_axb_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.control_input_axb_26 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.control_input_axb_20 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire \current_shift_inst.control_input_axb_21 ;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.control_input_axb_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.control_input_axb_23 ;
    wire il_max_comp1_D2;
    wire T01_c;
    wire state_3;
    wire s1_phy_c;
    wire \current_shift_inst.timer_s1.N_162_i ;
    wire s2_phy_c;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire bfn_14_11_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_14_12_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_14_13_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_14_14_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ;
    wire \current_shift_inst.un38_control_input_0_s1_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_8 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.un38_control_input_0_s1_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_16 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.un38_control_input_0_s1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_14_18_0_;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire elapsed_time_ns_1_RNITUBN9_0_10_cascade_;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_15_13_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_15_14_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire bfn_15_15_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire bfn_16_5_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_16_6_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_16_7_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_16_8_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.N_199_i ;
    wire bfn_16_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire bfn_16_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_16_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_16_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ;
    wire bfn_16_15_0_;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire bfn_16_16_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire bfn_16_17_0_;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire bfn_16_18_0_;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire bfn_16_19_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire bfn_16_20_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire bfn_16_21_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire bfn_16_22_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_17 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire T23_c;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_17_10_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_17_11_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire bfn_17_12_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire elapsed_time_ns_1_RNI36DN9_0_25_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire bfn_17_20_0_;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_17_21_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire bfn_17_22_0_;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire bfn_17_23_0_;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.N_198_i ;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire elapsed_time_ns_1_RNI68CN9_0_19_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_18_11_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_18_12_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_18_13_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_18_14_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.timer_s1.N_162_i_g ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_18_17_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_18_18_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_18_19_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_18_20_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_163_i ;
    wire T12_c;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire phase_controller_inst1_state_4;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17_cascade_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire elapsed_time_ns_1_RNI13CN9_0_14_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt28 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.state_RNIE87FZ0Z_2 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_start_g ;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt22 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire clock_output_0;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire red_c_g;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__23894),
            .RESETB(N__34067),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clock_output_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__48411),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__48408),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__27998,N__28024,N__28055,N__28082,N__28115,N__28141,N__28175,N__28208,N__27737,N__27763,N__27800,N__27833,N__27859,N__27899,N__27929,N__27962}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__48410,dangling_wire_45,N__48409}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__48348),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__48299),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__32470,N__32463,N__32468,N__32462,N__32469,N__32461,N__32471,N__32458,N__32464,N__32457,N__32465,N__32459,N__32466,N__32460,N__32467}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,N__48305,N__48302,dangling_wire_102,dangling_wire_103,dangling_wire_104,N__48300,N__48304,N__48301,N__48303}),
            .OHOLDTOP(),
            .O({dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__48436),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__48412),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .ADDSUBBOT(),
            .A({dangling_wire_136,N__32406,N__32409,N__32407,N__32410,N__32408,N__21328,N__21306,N__21250,N__21276,N__24108,N__24135,N__24165,N__20555,N__20573,N__20588}),
            .C({dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}),
            .B({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,N__48418,N__48415,dangling_wire_160,dangling_wire_161,dangling_wire_162,N__48413,N__48417,N__48414,N__48416}),
            .OHOLDTOP(),
            .O({dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__48371),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__48405),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .ADDSUBBOT(),
            .A({dangling_wire_185,N__27470,N__27493,N__27527,N__27557,N__27593,N__27626,N__27650,N__27680,N__27704,N__27271,N__27299,N__27329,N__27359,N__27385,N__29726}),
            .C({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201}),
            .B({dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,N__48407,dangling_wire_215,N__48406}),
            .OHOLDTOP(),
            .O({dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__50562),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__50564),
            .DIN(N__50563),
            .DOUT(N__50562),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__50564),
            .PADOUT(N__50563),
            .PADIN(N__50562),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clock_output_obuf_iopad (
            .OE(N__50553),
            .DIN(N__50552),
            .DOUT(N__50551),
            .PACKAGEPIN(clock_output));
    defparam clock_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam clock_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO clock_output_obuf_preio (
            .PADOEN(N__50553),
            .PADOUT(N__50552),
            .PADIN(N__50551),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26171),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T01_obuf_iopad (
            .OE(N__50544),
            .DIN(N__50543),
            .DOUT(N__50542),
            .PACKAGEPIN(T01));
    defparam T01_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T01_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T01_obuf_preio (
            .PADOEN(N__50544),
            .PADOUT(N__50543),
            .PADIN(N__50542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35654),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__50535),
            .DIN(N__50534),
            .DOUT(N__50533),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__50535),
            .PADOUT(N__50534),
            .PADIN(N__50533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__50526),
            .DIN(N__50525),
            .DOUT(N__50524),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__50526),
            .PADOUT(N__50525),
            .PADIN(N__50524),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__50517),
            .DIN(N__50516),
            .DOUT(N__50515),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__50517),
            .PADOUT(N__50516),
            .PADIN(N__50515),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__39818),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__50508),
            .DIN(N__50507),
            .DOUT(N__50506),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__50508),
            .PADOUT(N__50507),
            .PADIN(N__50506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24476),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__50499),
            .DIN(N__50498),
            .DOUT(N__50497),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__50499),
            .PADOUT(N__50498),
            .PADIN(N__50497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__50490),
            .DIN(N__50489),
            .DOUT(N__50488),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__50490),
            .PADOUT(N__50489),
            .PADIN(N__50488),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35870),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__50481),
            .DIN(N__50480),
            .DOUT(N__50479),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__50481),
            .PADOUT(N__50480),
            .PADIN(N__50479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__46502),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__50472),
            .DIN(N__50471),
            .DOUT(N__50470),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__50472),
            .PADOUT(N__50471),
            .PADIN(N__50470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__50463),
            .DIN(N__50462),
            .DOUT(N__50461),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__50463),
            .PADOUT(N__50462),
            .PADIN(N__50461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35588),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__50454),
            .DIN(N__50453),
            .DOUT(N__50452),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__50454),
            .PADOUT(N__50453),
            .PADIN(N__50452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26180),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__50445),
            .DIN(N__50444),
            .DOUT(N__50443),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__50445),
            .PADOUT(N__50444),
            .PADIN(N__50443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__50436),
            .DIN(N__50435),
            .DOUT(N__50434),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__50436),
            .PADOUT(N__50435),
            .PADIN(N__50434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26234),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T45_obuf_iopad (
            .OE(N__50427),
            .DIN(N__50426),
            .DOUT(N__50425),
            .PACKAGEPIN(T45));
    defparam T45_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T45_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T45_obuf_preio (
            .PADOEN(N__50427),
            .PADOUT(N__50426),
            .PADIN(N__50425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31802),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__50418),
            .DIN(N__50417),
            .DOUT(N__50416),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__50418),
            .PADOUT(N__50417),
            .PADIN(N__50416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__50409),
            .DIN(N__50408),
            .DOUT(N__50407),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__50409),
            .PADOUT(N__50408),
            .PADIN(N__50407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11986 (
            .O(N__50390),
            .I(N__50387));
    LocalMux I__11985 (
            .O(N__50387),
            .I(N__50382));
    InMux I__11984 (
            .O(N__50386),
            .I(N__50379));
    InMux I__11983 (
            .O(N__50385),
            .I(N__50376));
    Span4Mux_v I__11982 (
            .O(N__50382),
            .I(N__50371));
    LocalMux I__11981 (
            .O(N__50379),
            .I(N__50371));
    LocalMux I__11980 (
            .O(N__50376),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    Odrv4 I__11979 (
            .O(N__50371),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    InMux I__11978 (
            .O(N__50366),
            .I(N__50363));
    LocalMux I__11977 (
            .O(N__50363),
            .I(N__50359));
    InMux I__11976 (
            .O(N__50362),
            .I(N__50356));
    Span4Mux_v I__11975 (
            .O(N__50359),
            .I(N__50349));
    LocalMux I__11974 (
            .O(N__50356),
            .I(N__50349));
    InMux I__11973 (
            .O(N__50355),
            .I(N__50346));
    InMux I__11972 (
            .O(N__50354),
            .I(N__50343));
    Span4Mux_v I__11971 (
            .O(N__50349),
            .I(N__50338));
    LocalMux I__11970 (
            .O(N__50346),
            .I(N__50338));
    LocalMux I__11969 (
            .O(N__50343),
            .I(N__50335));
    Span4Mux_h I__11968 (
            .O(N__50338),
            .I(N__50332));
    Span4Mux_h I__11967 (
            .O(N__50335),
            .I(N__50329));
    Odrv4 I__11966 (
            .O(N__50332),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__11965 (
            .O(N__50329),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__11964 (
            .O(N__50324),
            .I(N__50321));
    LocalMux I__11963 (
            .O(N__50321),
            .I(N__50166));
    ClkMux I__11962 (
            .O(N__50320),
            .I(N__49856));
    ClkMux I__11961 (
            .O(N__50319),
            .I(N__49856));
    ClkMux I__11960 (
            .O(N__50318),
            .I(N__49856));
    ClkMux I__11959 (
            .O(N__50317),
            .I(N__49856));
    ClkMux I__11958 (
            .O(N__50316),
            .I(N__49856));
    ClkMux I__11957 (
            .O(N__50315),
            .I(N__49856));
    ClkMux I__11956 (
            .O(N__50314),
            .I(N__49856));
    ClkMux I__11955 (
            .O(N__50313),
            .I(N__49856));
    ClkMux I__11954 (
            .O(N__50312),
            .I(N__49856));
    ClkMux I__11953 (
            .O(N__50311),
            .I(N__49856));
    ClkMux I__11952 (
            .O(N__50310),
            .I(N__49856));
    ClkMux I__11951 (
            .O(N__50309),
            .I(N__49856));
    ClkMux I__11950 (
            .O(N__50308),
            .I(N__49856));
    ClkMux I__11949 (
            .O(N__50307),
            .I(N__49856));
    ClkMux I__11948 (
            .O(N__50306),
            .I(N__49856));
    ClkMux I__11947 (
            .O(N__50305),
            .I(N__49856));
    ClkMux I__11946 (
            .O(N__50304),
            .I(N__49856));
    ClkMux I__11945 (
            .O(N__50303),
            .I(N__49856));
    ClkMux I__11944 (
            .O(N__50302),
            .I(N__49856));
    ClkMux I__11943 (
            .O(N__50301),
            .I(N__49856));
    ClkMux I__11942 (
            .O(N__50300),
            .I(N__49856));
    ClkMux I__11941 (
            .O(N__50299),
            .I(N__49856));
    ClkMux I__11940 (
            .O(N__50298),
            .I(N__49856));
    ClkMux I__11939 (
            .O(N__50297),
            .I(N__49856));
    ClkMux I__11938 (
            .O(N__50296),
            .I(N__49856));
    ClkMux I__11937 (
            .O(N__50295),
            .I(N__49856));
    ClkMux I__11936 (
            .O(N__50294),
            .I(N__49856));
    ClkMux I__11935 (
            .O(N__50293),
            .I(N__49856));
    ClkMux I__11934 (
            .O(N__50292),
            .I(N__49856));
    ClkMux I__11933 (
            .O(N__50291),
            .I(N__49856));
    ClkMux I__11932 (
            .O(N__50290),
            .I(N__49856));
    ClkMux I__11931 (
            .O(N__50289),
            .I(N__49856));
    ClkMux I__11930 (
            .O(N__50288),
            .I(N__49856));
    ClkMux I__11929 (
            .O(N__50287),
            .I(N__49856));
    ClkMux I__11928 (
            .O(N__50286),
            .I(N__49856));
    ClkMux I__11927 (
            .O(N__50285),
            .I(N__49856));
    ClkMux I__11926 (
            .O(N__50284),
            .I(N__49856));
    ClkMux I__11925 (
            .O(N__50283),
            .I(N__49856));
    ClkMux I__11924 (
            .O(N__50282),
            .I(N__49856));
    ClkMux I__11923 (
            .O(N__50281),
            .I(N__49856));
    ClkMux I__11922 (
            .O(N__50280),
            .I(N__49856));
    ClkMux I__11921 (
            .O(N__50279),
            .I(N__49856));
    ClkMux I__11920 (
            .O(N__50278),
            .I(N__49856));
    ClkMux I__11919 (
            .O(N__50277),
            .I(N__49856));
    ClkMux I__11918 (
            .O(N__50276),
            .I(N__49856));
    ClkMux I__11917 (
            .O(N__50275),
            .I(N__49856));
    ClkMux I__11916 (
            .O(N__50274),
            .I(N__49856));
    ClkMux I__11915 (
            .O(N__50273),
            .I(N__49856));
    ClkMux I__11914 (
            .O(N__50272),
            .I(N__49856));
    ClkMux I__11913 (
            .O(N__50271),
            .I(N__49856));
    ClkMux I__11912 (
            .O(N__50270),
            .I(N__49856));
    ClkMux I__11911 (
            .O(N__50269),
            .I(N__49856));
    ClkMux I__11910 (
            .O(N__50268),
            .I(N__49856));
    ClkMux I__11909 (
            .O(N__50267),
            .I(N__49856));
    ClkMux I__11908 (
            .O(N__50266),
            .I(N__49856));
    ClkMux I__11907 (
            .O(N__50265),
            .I(N__49856));
    ClkMux I__11906 (
            .O(N__50264),
            .I(N__49856));
    ClkMux I__11905 (
            .O(N__50263),
            .I(N__49856));
    ClkMux I__11904 (
            .O(N__50262),
            .I(N__49856));
    ClkMux I__11903 (
            .O(N__50261),
            .I(N__49856));
    ClkMux I__11902 (
            .O(N__50260),
            .I(N__49856));
    ClkMux I__11901 (
            .O(N__50259),
            .I(N__49856));
    ClkMux I__11900 (
            .O(N__50258),
            .I(N__49856));
    ClkMux I__11899 (
            .O(N__50257),
            .I(N__49856));
    ClkMux I__11898 (
            .O(N__50256),
            .I(N__49856));
    ClkMux I__11897 (
            .O(N__50255),
            .I(N__49856));
    ClkMux I__11896 (
            .O(N__50254),
            .I(N__49856));
    ClkMux I__11895 (
            .O(N__50253),
            .I(N__49856));
    ClkMux I__11894 (
            .O(N__50252),
            .I(N__49856));
    ClkMux I__11893 (
            .O(N__50251),
            .I(N__49856));
    ClkMux I__11892 (
            .O(N__50250),
            .I(N__49856));
    ClkMux I__11891 (
            .O(N__50249),
            .I(N__49856));
    ClkMux I__11890 (
            .O(N__50248),
            .I(N__49856));
    ClkMux I__11889 (
            .O(N__50247),
            .I(N__49856));
    ClkMux I__11888 (
            .O(N__50246),
            .I(N__49856));
    ClkMux I__11887 (
            .O(N__50245),
            .I(N__49856));
    ClkMux I__11886 (
            .O(N__50244),
            .I(N__49856));
    ClkMux I__11885 (
            .O(N__50243),
            .I(N__49856));
    ClkMux I__11884 (
            .O(N__50242),
            .I(N__49856));
    ClkMux I__11883 (
            .O(N__50241),
            .I(N__49856));
    ClkMux I__11882 (
            .O(N__50240),
            .I(N__49856));
    ClkMux I__11881 (
            .O(N__50239),
            .I(N__49856));
    ClkMux I__11880 (
            .O(N__50238),
            .I(N__49856));
    ClkMux I__11879 (
            .O(N__50237),
            .I(N__49856));
    ClkMux I__11878 (
            .O(N__50236),
            .I(N__49856));
    ClkMux I__11877 (
            .O(N__50235),
            .I(N__49856));
    ClkMux I__11876 (
            .O(N__50234),
            .I(N__49856));
    ClkMux I__11875 (
            .O(N__50233),
            .I(N__49856));
    ClkMux I__11874 (
            .O(N__50232),
            .I(N__49856));
    ClkMux I__11873 (
            .O(N__50231),
            .I(N__49856));
    ClkMux I__11872 (
            .O(N__50230),
            .I(N__49856));
    ClkMux I__11871 (
            .O(N__50229),
            .I(N__49856));
    ClkMux I__11870 (
            .O(N__50228),
            .I(N__49856));
    ClkMux I__11869 (
            .O(N__50227),
            .I(N__49856));
    ClkMux I__11868 (
            .O(N__50226),
            .I(N__49856));
    ClkMux I__11867 (
            .O(N__50225),
            .I(N__49856));
    ClkMux I__11866 (
            .O(N__50224),
            .I(N__49856));
    ClkMux I__11865 (
            .O(N__50223),
            .I(N__49856));
    ClkMux I__11864 (
            .O(N__50222),
            .I(N__49856));
    ClkMux I__11863 (
            .O(N__50221),
            .I(N__49856));
    ClkMux I__11862 (
            .O(N__50220),
            .I(N__49856));
    ClkMux I__11861 (
            .O(N__50219),
            .I(N__49856));
    ClkMux I__11860 (
            .O(N__50218),
            .I(N__49856));
    ClkMux I__11859 (
            .O(N__50217),
            .I(N__49856));
    ClkMux I__11858 (
            .O(N__50216),
            .I(N__49856));
    ClkMux I__11857 (
            .O(N__50215),
            .I(N__49856));
    ClkMux I__11856 (
            .O(N__50214),
            .I(N__49856));
    ClkMux I__11855 (
            .O(N__50213),
            .I(N__49856));
    ClkMux I__11854 (
            .O(N__50212),
            .I(N__49856));
    ClkMux I__11853 (
            .O(N__50211),
            .I(N__49856));
    ClkMux I__11852 (
            .O(N__50210),
            .I(N__49856));
    ClkMux I__11851 (
            .O(N__50209),
            .I(N__49856));
    ClkMux I__11850 (
            .O(N__50208),
            .I(N__49856));
    ClkMux I__11849 (
            .O(N__50207),
            .I(N__49856));
    ClkMux I__11848 (
            .O(N__50206),
            .I(N__49856));
    ClkMux I__11847 (
            .O(N__50205),
            .I(N__49856));
    ClkMux I__11846 (
            .O(N__50204),
            .I(N__49856));
    ClkMux I__11845 (
            .O(N__50203),
            .I(N__49856));
    ClkMux I__11844 (
            .O(N__50202),
            .I(N__49856));
    ClkMux I__11843 (
            .O(N__50201),
            .I(N__49856));
    ClkMux I__11842 (
            .O(N__50200),
            .I(N__49856));
    ClkMux I__11841 (
            .O(N__50199),
            .I(N__49856));
    ClkMux I__11840 (
            .O(N__50198),
            .I(N__49856));
    ClkMux I__11839 (
            .O(N__50197),
            .I(N__49856));
    ClkMux I__11838 (
            .O(N__50196),
            .I(N__49856));
    ClkMux I__11837 (
            .O(N__50195),
            .I(N__49856));
    ClkMux I__11836 (
            .O(N__50194),
            .I(N__49856));
    ClkMux I__11835 (
            .O(N__50193),
            .I(N__49856));
    ClkMux I__11834 (
            .O(N__50192),
            .I(N__49856));
    ClkMux I__11833 (
            .O(N__50191),
            .I(N__49856));
    ClkMux I__11832 (
            .O(N__50190),
            .I(N__49856));
    ClkMux I__11831 (
            .O(N__50189),
            .I(N__49856));
    ClkMux I__11830 (
            .O(N__50188),
            .I(N__49856));
    ClkMux I__11829 (
            .O(N__50187),
            .I(N__49856));
    ClkMux I__11828 (
            .O(N__50186),
            .I(N__49856));
    ClkMux I__11827 (
            .O(N__50185),
            .I(N__49856));
    ClkMux I__11826 (
            .O(N__50184),
            .I(N__49856));
    ClkMux I__11825 (
            .O(N__50183),
            .I(N__49856));
    ClkMux I__11824 (
            .O(N__50182),
            .I(N__49856));
    ClkMux I__11823 (
            .O(N__50181),
            .I(N__49856));
    ClkMux I__11822 (
            .O(N__50180),
            .I(N__49856));
    ClkMux I__11821 (
            .O(N__50179),
            .I(N__49856));
    ClkMux I__11820 (
            .O(N__50178),
            .I(N__49856));
    ClkMux I__11819 (
            .O(N__50177),
            .I(N__49856));
    ClkMux I__11818 (
            .O(N__50176),
            .I(N__49856));
    ClkMux I__11817 (
            .O(N__50175),
            .I(N__49856));
    ClkMux I__11816 (
            .O(N__50174),
            .I(N__49856));
    ClkMux I__11815 (
            .O(N__50173),
            .I(N__49856));
    ClkMux I__11814 (
            .O(N__50172),
            .I(N__49856));
    ClkMux I__11813 (
            .O(N__50171),
            .I(N__49856));
    ClkMux I__11812 (
            .O(N__50170),
            .I(N__49856));
    ClkMux I__11811 (
            .O(N__50169),
            .I(N__49856));
    Glb2LocalMux I__11810 (
            .O(N__50166),
            .I(N__49856));
    ClkMux I__11809 (
            .O(N__50165),
            .I(N__49856));
    GlobalMux I__11808 (
            .O(N__49856),
            .I(clock_output_0));
    InMux I__11807 (
            .O(N__49853),
            .I(N__49840));
    InMux I__11806 (
            .O(N__49852),
            .I(N__49840));
    InMux I__11805 (
            .O(N__49851),
            .I(N__49840));
    InMux I__11804 (
            .O(N__49850),
            .I(N__49823));
    InMux I__11803 (
            .O(N__49849),
            .I(N__49823));
    InMux I__11802 (
            .O(N__49848),
            .I(N__49823));
    InMux I__11801 (
            .O(N__49847),
            .I(N__49823));
    LocalMux I__11800 (
            .O(N__49840),
            .I(N__49820));
    InMux I__11799 (
            .O(N__49839),
            .I(N__49811));
    InMux I__11798 (
            .O(N__49838),
            .I(N__49811));
    InMux I__11797 (
            .O(N__49837),
            .I(N__49811));
    InMux I__11796 (
            .O(N__49836),
            .I(N__49811));
    CEMux I__11795 (
            .O(N__49835),
            .I(N__49808));
    CEMux I__11794 (
            .O(N__49834),
            .I(N__49800));
    InMux I__11793 (
            .O(N__49833),
            .I(N__49796));
    CEMux I__11792 (
            .O(N__49832),
            .I(N__49793));
    LocalMux I__11791 (
            .O(N__49823),
            .I(N__49781));
    Span4Mux_h I__11790 (
            .O(N__49820),
            .I(N__49781));
    LocalMux I__11789 (
            .O(N__49811),
            .I(N__49781));
    LocalMux I__11788 (
            .O(N__49808),
            .I(N__49778));
    CEMux I__11787 (
            .O(N__49807),
            .I(N__49763));
    CEMux I__11786 (
            .O(N__49806),
            .I(N__49760));
    CEMux I__11785 (
            .O(N__49805),
            .I(N__49757));
    CEMux I__11784 (
            .O(N__49804),
            .I(N__49754));
    CEMux I__11783 (
            .O(N__49803),
            .I(N__49751));
    LocalMux I__11782 (
            .O(N__49800),
            .I(N__49748));
    CEMux I__11781 (
            .O(N__49799),
            .I(N__49741));
    LocalMux I__11780 (
            .O(N__49796),
            .I(N__49736));
    LocalMux I__11779 (
            .O(N__49793),
            .I(N__49736));
    CEMux I__11778 (
            .O(N__49792),
            .I(N__49730));
    CEMux I__11777 (
            .O(N__49791),
            .I(N__49727));
    InMux I__11776 (
            .O(N__49790),
            .I(N__49720));
    InMux I__11775 (
            .O(N__49789),
            .I(N__49720));
    InMux I__11774 (
            .O(N__49788),
            .I(N__49720));
    Span4Mux_v I__11773 (
            .O(N__49781),
            .I(N__49715));
    Span4Mux_v I__11772 (
            .O(N__49778),
            .I(N__49715));
    InMux I__11771 (
            .O(N__49777),
            .I(N__49706));
    InMux I__11770 (
            .O(N__49776),
            .I(N__49706));
    InMux I__11769 (
            .O(N__49775),
            .I(N__49706));
    InMux I__11768 (
            .O(N__49774),
            .I(N__49706));
    InMux I__11767 (
            .O(N__49773),
            .I(N__49697));
    InMux I__11766 (
            .O(N__49772),
            .I(N__49697));
    InMux I__11765 (
            .O(N__49771),
            .I(N__49697));
    InMux I__11764 (
            .O(N__49770),
            .I(N__49697));
    InMux I__11763 (
            .O(N__49769),
            .I(N__49688));
    InMux I__11762 (
            .O(N__49768),
            .I(N__49688));
    InMux I__11761 (
            .O(N__49767),
            .I(N__49688));
    InMux I__11760 (
            .O(N__49766),
            .I(N__49688));
    LocalMux I__11759 (
            .O(N__49763),
            .I(N__49685));
    LocalMux I__11758 (
            .O(N__49760),
            .I(N__49680));
    LocalMux I__11757 (
            .O(N__49757),
            .I(N__49680));
    LocalMux I__11756 (
            .O(N__49754),
            .I(N__49677));
    LocalMux I__11755 (
            .O(N__49751),
            .I(N__49672));
    Span4Mux_h I__11754 (
            .O(N__49748),
            .I(N__49672));
    InMux I__11753 (
            .O(N__49747),
            .I(N__49663));
    InMux I__11752 (
            .O(N__49746),
            .I(N__49663));
    InMux I__11751 (
            .O(N__49745),
            .I(N__49663));
    InMux I__11750 (
            .O(N__49744),
            .I(N__49663));
    LocalMux I__11749 (
            .O(N__49741),
            .I(N__49660));
    Span4Mux_v I__11748 (
            .O(N__49736),
            .I(N__49657));
    CEMux I__11747 (
            .O(N__49735),
            .I(N__49654));
    CEMux I__11746 (
            .O(N__49734),
            .I(N__49651));
    CEMux I__11745 (
            .O(N__49733),
            .I(N__49648));
    LocalMux I__11744 (
            .O(N__49730),
            .I(N__49645));
    LocalMux I__11743 (
            .O(N__49727),
            .I(N__49642));
    LocalMux I__11742 (
            .O(N__49720),
            .I(N__49631));
    Span4Mux_h I__11741 (
            .O(N__49715),
            .I(N__49631));
    LocalMux I__11740 (
            .O(N__49706),
            .I(N__49631));
    LocalMux I__11739 (
            .O(N__49697),
            .I(N__49631));
    LocalMux I__11738 (
            .O(N__49688),
            .I(N__49631));
    Span4Mux_h I__11737 (
            .O(N__49685),
            .I(N__49628));
    Sp12to4 I__11736 (
            .O(N__49680),
            .I(N__49625));
    Span4Mux_v I__11735 (
            .O(N__49677),
            .I(N__49614));
    Span4Mux_v I__11734 (
            .O(N__49672),
            .I(N__49614));
    LocalMux I__11733 (
            .O(N__49663),
            .I(N__49614));
    Span4Mux_v I__11732 (
            .O(N__49660),
            .I(N__49614));
    Span4Mux_h I__11731 (
            .O(N__49657),
            .I(N__49614));
    LocalMux I__11730 (
            .O(N__49654),
            .I(N__49611));
    LocalMux I__11729 (
            .O(N__49651),
            .I(N__49608));
    LocalMux I__11728 (
            .O(N__49648),
            .I(N__49603));
    Span4Mux_h I__11727 (
            .O(N__49645),
            .I(N__49603));
    Span4Mux_h I__11726 (
            .O(N__49642),
            .I(N__49598));
    Span4Mux_v I__11725 (
            .O(N__49631),
            .I(N__49598));
    Span4Mux_h I__11724 (
            .O(N__49628),
            .I(N__49595));
    Span12Mux_s9_v I__11723 (
            .O(N__49625),
            .I(N__49592));
    Span4Mux_h I__11722 (
            .O(N__49614),
            .I(N__49589));
    Odrv4 I__11721 (
            .O(N__49611),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv12 I__11720 (
            .O(N__49608),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11719 (
            .O(N__49603),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11718 (
            .O(N__49598),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11717 (
            .O(N__49595),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv12 I__11716 (
            .O(N__49592),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11715 (
            .O(N__49589),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__11714 (
            .O(N__49574),
            .I(N__49568));
    InMux I__11713 (
            .O(N__49573),
            .I(N__49565));
    InMux I__11712 (
            .O(N__49572),
            .I(N__49562));
    InMux I__11711 (
            .O(N__49571),
            .I(N__49559));
    LocalMux I__11710 (
            .O(N__49568),
            .I(N__49556));
    LocalMux I__11709 (
            .O(N__49565),
            .I(N__49553));
    LocalMux I__11708 (
            .O(N__49562),
            .I(N__49545));
    LocalMux I__11707 (
            .O(N__49559),
            .I(N__49541));
    Glb2LocalMux I__11706 (
            .O(N__49556),
            .I(N__49076));
    Glb2LocalMux I__11705 (
            .O(N__49553),
            .I(N__49076));
    SRMux I__11704 (
            .O(N__49552),
            .I(N__49076));
    SRMux I__11703 (
            .O(N__49551),
            .I(N__49076));
    SRMux I__11702 (
            .O(N__49550),
            .I(N__49076));
    SRMux I__11701 (
            .O(N__49549),
            .I(N__49076));
    SRMux I__11700 (
            .O(N__49548),
            .I(N__49076));
    Glb2LocalMux I__11699 (
            .O(N__49545),
            .I(N__49076));
    SRMux I__11698 (
            .O(N__49544),
            .I(N__49076));
    Glb2LocalMux I__11697 (
            .O(N__49541),
            .I(N__49076));
    SRMux I__11696 (
            .O(N__49540),
            .I(N__49076));
    SRMux I__11695 (
            .O(N__49539),
            .I(N__49076));
    SRMux I__11694 (
            .O(N__49538),
            .I(N__49076));
    SRMux I__11693 (
            .O(N__49537),
            .I(N__49076));
    SRMux I__11692 (
            .O(N__49536),
            .I(N__49076));
    SRMux I__11691 (
            .O(N__49535),
            .I(N__49076));
    SRMux I__11690 (
            .O(N__49534),
            .I(N__49076));
    SRMux I__11689 (
            .O(N__49533),
            .I(N__49076));
    SRMux I__11688 (
            .O(N__49532),
            .I(N__49076));
    SRMux I__11687 (
            .O(N__49531),
            .I(N__49076));
    SRMux I__11686 (
            .O(N__49530),
            .I(N__49076));
    SRMux I__11685 (
            .O(N__49529),
            .I(N__49076));
    SRMux I__11684 (
            .O(N__49528),
            .I(N__49076));
    SRMux I__11683 (
            .O(N__49527),
            .I(N__49076));
    SRMux I__11682 (
            .O(N__49526),
            .I(N__49076));
    SRMux I__11681 (
            .O(N__49525),
            .I(N__49076));
    SRMux I__11680 (
            .O(N__49524),
            .I(N__49076));
    SRMux I__11679 (
            .O(N__49523),
            .I(N__49076));
    SRMux I__11678 (
            .O(N__49522),
            .I(N__49076));
    SRMux I__11677 (
            .O(N__49521),
            .I(N__49076));
    SRMux I__11676 (
            .O(N__49520),
            .I(N__49076));
    SRMux I__11675 (
            .O(N__49519),
            .I(N__49076));
    SRMux I__11674 (
            .O(N__49518),
            .I(N__49076));
    SRMux I__11673 (
            .O(N__49517),
            .I(N__49076));
    SRMux I__11672 (
            .O(N__49516),
            .I(N__49076));
    SRMux I__11671 (
            .O(N__49515),
            .I(N__49076));
    SRMux I__11670 (
            .O(N__49514),
            .I(N__49076));
    SRMux I__11669 (
            .O(N__49513),
            .I(N__49076));
    SRMux I__11668 (
            .O(N__49512),
            .I(N__49076));
    SRMux I__11667 (
            .O(N__49511),
            .I(N__49076));
    SRMux I__11666 (
            .O(N__49510),
            .I(N__49076));
    SRMux I__11665 (
            .O(N__49509),
            .I(N__49076));
    SRMux I__11664 (
            .O(N__49508),
            .I(N__49076));
    SRMux I__11663 (
            .O(N__49507),
            .I(N__49076));
    SRMux I__11662 (
            .O(N__49506),
            .I(N__49076));
    SRMux I__11661 (
            .O(N__49505),
            .I(N__49076));
    SRMux I__11660 (
            .O(N__49504),
            .I(N__49076));
    SRMux I__11659 (
            .O(N__49503),
            .I(N__49076));
    SRMux I__11658 (
            .O(N__49502),
            .I(N__49076));
    SRMux I__11657 (
            .O(N__49501),
            .I(N__49076));
    SRMux I__11656 (
            .O(N__49500),
            .I(N__49076));
    SRMux I__11655 (
            .O(N__49499),
            .I(N__49076));
    SRMux I__11654 (
            .O(N__49498),
            .I(N__49076));
    SRMux I__11653 (
            .O(N__49497),
            .I(N__49076));
    SRMux I__11652 (
            .O(N__49496),
            .I(N__49076));
    SRMux I__11651 (
            .O(N__49495),
            .I(N__49076));
    SRMux I__11650 (
            .O(N__49494),
            .I(N__49076));
    SRMux I__11649 (
            .O(N__49493),
            .I(N__49076));
    SRMux I__11648 (
            .O(N__49492),
            .I(N__49076));
    SRMux I__11647 (
            .O(N__49491),
            .I(N__49076));
    SRMux I__11646 (
            .O(N__49490),
            .I(N__49076));
    SRMux I__11645 (
            .O(N__49489),
            .I(N__49076));
    SRMux I__11644 (
            .O(N__49488),
            .I(N__49076));
    SRMux I__11643 (
            .O(N__49487),
            .I(N__49076));
    SRMux I__11642 (
            .O(N__49486),
            .I(N__49076));
    SRMux I__11641 (
            .O(N__49485),
            .I(N__49076));
    SRMux I__11640 (
            .O(N__49484),
            .I(N__49076));
    SRMux I__11639 (
            .O(N__49483),
            .I(N__49076));
    SRMux I__11638 (
            .O(N__49482),
            .I(N__49076));
    SRMux I__11637 (
            .O(N__49481),
            .I(N__49076));
    SRMux I__11636 (
            .O(N__49480),
            .I(N__49076));
    SRMux I__11635 (
            .O(N__49479),
            .I(N__49076));
    SRMux I__11634 (
            .O(N__49478),
            .I(N__49076));
    SRMux I__11633 (
            .O(N__49477),
            .I(N__49076));
    SRMux I__11632 (
            .O(N__49476),
            .I(N__49076));
    SRMux I__11631 (
            .O(N__49475),
            .I(N__49076));
    SRMux I__11630 (
            .O(N__49474),
            .I(N__49076));
    SRMux I__11629 (
            .O(N__49473),
            .I(N__49076));
    SRMux I__11628 (
            .O(N__49472),
            .I(N__49076));
    SRMux I__11627 (
            .O(N__49471),
            .I(N__49076));
    SRMux I__11626 (
            .O(N__49470),
            .I(N__49076));
    SRMux I__11625 (
            .O(N__49469),
            .I(N__49076));
    SRMux I__11624 (
            .O(N__49468),
            .I(N__49076));
    SRMux I__11623 (
            .O(N__49467),
            .I(N__49076));
    SRMux I__11622 (
            .O(N__49466),
            .I(N__49076));
    SRMux I__11621 (
            .O(N__49465),
            .I(N__49076));
    SRMux I__11620 (
            .O(N__49464),
            .I(N__49076));
    SRMux I__11619 (
            .O(N__49463),
            .I(N__49076));
    SRMux I__11618 (
            .O(N__49462),
            .I(N__49076));
    SRMux I__11617 (
            .O(N__49461),
            .I(N__49076));
    SRMux I__11616 (
            .O(N__49460),
            .I(N__49076));
    SRMux I__11615 (
            .O(N__49459),
            .I(N__49076));
    SRMux I__11614 (
            .O(N__49458),
            .I(N__49076));
    SRMux I__11613 (
            .O(N__49457),
            .I(N__49076));
    SRMux I__11612 (
            .O(N__49456),
            .I(N__49076));
    SRMux I__11611 (
            .O(N__49455),
            .I(N__49076));
    SRMux I__11610 (
            .O(N__49454),
            .I(N__49076));
    SRMux I__11609 (
            .O(N__49453),
            .I(N__49076));
    SRMux I__11608 (
            .O(N__49452),
            .I(N__49076));
    SRMux I__11607 (
            .O(N__49451),
            .I(N__49076));
    SRMux I__11606 (
            .O(N__49450),
            .I(N__49076));
    SRMux I__11605 (
            .O(N__49449),
            .I(N__49076));
    SRMux I__11604 (
            .O(N__49448),
            .I(N__49076));
    SRMux I__11603 (
            .O(N__49447),
            .I(N__49076));
    SRMux I__11602 (
            .O(N__49446),
            .I(N__49076));
    SRMux I__11601 (
            .O(N__49445),
            .I(N__49076));
    SRMux I__11600 (
            .O(N__49444),
            .I(N__49076));
    SRMux I__11599 (
            .O(N__49443),
            .I(N__49076));
    SRMux I__11598 (
            .O(N__49442),
            .I(N__49076));
    SRMux I__11597 (
            .O(N__49441),
            .I(N__49076));
    SRMux I__11596 (
            .O(N__49440),
            .I(N__49076));
    SRMux I__11595 (
            .O(N__49439),
            .I(N__49076));
    SRMux I__11594 (
            .O(N__49438),
            .I(N__49076));
    SRMux I__11593 (
            .O(N__49437),
            .I(N__49076));
    SRMux I__11592 (
            .O(N__49436),
            .I(N__49076));
    SRMux I__11591 (
            .O(N__49435),
            .I(N__49076));
    SRMux I__11590 (
            .O(N__49434),
            .I(N__49076));
    SRMux I__11589 (
            .O(N__49433),
            .I(N__49076));
    SRMux I__11588 (
            .O(N__49432),
            .I(N__49076));
    SRMux I__11587 (
            .O(N__49431),
            .I(N__49076));
    SRMux I__11586 (
            .O(N__49430),
            .I(N__49076));
    SRMux I__11585 (
            .O(N__49429),
            .I(N__49076));
    SRMux I__11584 (
            .O(N__49428),
            .I(N__49076));
    SRMux I__11583 (
            .O(N__49427),
            .I(N__49076));
    SRMux I__11582 (
            .O(N__49426),
            .I(N__49076));
    SRMux I__11581 (
            .O(N__49425),
            .I(N__49076));
    SRMux I__11580 (
            .O(N__49424),
            .I(N__49076));
    SRMux I__11579 (
            .O(N__49423),
            .I(N__49076));
    SRMux I__11578 (
            .O(N__49422),
            .I(N__49076));
    SRMux I__11577 (
            .O(N__49421),
            .I(N__49076));
    SRMux I__11576 (
            .O(N__49420),
            .I(N__49076));
    SRMux I__11575 (
            .O(N__49419),
            .I(N__49076));
    SRMux I__11574 (
            .O(N__49418),
            .I(N__49076));
    SRMux I__11573 (
            .O(N__49417),
            .I(N__49076));
    SRMux I__11572 (
            .O(N__49416),
            .I(N__49076));
    SRMux I__11571 (
            .O(N__49415),
            .I(N__49076));
    SRMux I__11570 (
            .O(N__49414),
            .I(N__49076));
    SRMux I__11569 (
            .O(N__49413),
            .I(N__49076));
    SRMux I__11568 (
            .O(N__49412),
            .I(N__49076));
    SRMux I__11567 (
            .O(N__49411),
            .I(N__49076));
    SRMux I__11566 (
            .O(N__49410),
            .I(N__49076));
    SRMux I__11565 (
            .O(N__49409),
            .I(N__49076));
    SRMux I__11564 (
            .O(N__49408),
            .I(N__49076));
    SRMux I__11563 (
            .O(N__49407),
            .I(N__49076));
    SRMux I__11562 (
            .O(N__49406),
            .I(N__49076));
    SRMux I__11561 (
            .O(N__49405),
            .I(N__49076));
    SRMux I__11560 (
            .O(N__49404),
            .I(N__49076));
    SRMux I__11559 (
            .O(N__49403),
            .I(N__49076));
    SRMux I__11558 (
            .O(N__49402),
            .I(N__49076));
    SRMux I__11557 (
            .O(N__49401),
            .I(N__49076));
    SRMux I__11556 (
            .O(N__49400),
            .I(N__49076));
    SRMux I__11555 (
            .O(N__49399),
            .I(N__49076));
    SRMux I__11554 (
            .O(N__49398),
            .I(N__49076));
    SRMux I__11553 (
            .O(N__49397),
            .I(N__49076));
    SRMux I__11552 (
            .O(N__49396),
            .I(N__49076));
    SRMux I__11551 (
            .O(N__49395),
            .I(N__49076));
    SRMux I__11550 (
            .O(N__49394),
            .I(N__49076));
    SRMux I__11549 (
            .O(N__49393),
            .I(N__49076));
    GlobalMux I__11548 (
            .O(N__49076),
            .I(N__49073));
    gio2CtrlBuf I__11547 (
            .O(N__49073),
            .I(red_c_g));
    CascadeMux I__11546 (
            .O(N__49070),
            .I(N__49067));
    InMux I__11545 (
            .O(N__49067),
            .I(N__49064));
    LocalMux I__11544 (
            .O(N__49064),
            .I(N__49061));
    Span4Mux_h I__11543 (
            .O(N__49061),
            .I(N__49058));
    Odrv4 I__11542 (
            .O(N__49058),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt26 ));
    InMux I__11541 (
            .O(N__49055),
            .I(N__49049));
    InMux I__11540 (
            .O(N__49054),
            .I(N__49049));
    LocalMux I__11539 (
            .O(N__49049),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ));
    InMux I__11538 (
            .O(N__49046),
            .I(N__49039));
    InMux I__11537 (
            .O(N__49045),
            .I(N__49039));
    InMux I__11536 (
            .O(N__49044),
            .I(N__49036));
    LocalMux I__11535 (
            .O(N__49039),
            .I(N__49033));
    LocalMux I__11534 (
            .O(N__49036),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    Odrv4 I__11533 (
            .O(N__49033),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    CascadeMux I__11532 (
            .O(N__49028),
            .I(N__49024));
    CascadeMux I__11531 (
            .O(N__49027),
            .I(N__49021));
    InMux I__11530 (
            .O(N__49024),
            .I(N__49015));
    InMux I__11529 (
            .O(N__49021),
            .I(N__49015));
    InMux I__11528 (
            .O(N__49020),
            .I(N__49012));
    LocalMux I__11527 (
            .O(N__49015),
            .I(N__49009));
    LocalMux I__11526 (
            .O(N__49012),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    Odrv4 I__11525 (
            .O(N__49009),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__11524 (
            .O(N__49004),
            .I(N__48998));
    InMux I__11523 (
            .O(N__49003),
            .I(N__48998));
    LocalMux I__11522 (
            .O(N__48998),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ));
    InMux I__11521 (
            .O(N__48995),
            .I(N__48992));
    LocalMux I__11520 (
            .O(N__48992),
            .I(N__48989));
    Span4Mux_h I__11519 (
            .O(N__48989),
            .I(N__48986));
    Odrv4 I__11518 (
            .O(N__48986),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ));
    InMux I__11517 (
            .O(N__48983),
            .I(N__48979));
    InMux I__11516 (
            .O(N__48982),
            .I(N__48975));
    LocalMux I__11515 (
            .O(N__48979),
            .I(N__48972));
    InMux I__11514 (
            .O(N__48978),
            .I(N__48969));
    LocalMux I__11513 (
            .O(N__48975),
            .I(N__48965));
    Span4Mux_v I__11512 (
            .O(N__48972),
            .I(N__48960));
    LocalMux I__11511 (
            .O(N__48969),
            .I(N__48960));
    InMux I__11510 (
            .O(N__48968),
            .I(N__48957));
    Span4Mux_v I__11509 (
            .O(N__48965),
            .I(N__48954));
    Span4Mux_v I__11508 (
            .O(N__48960),
            .I(N__48949));
    LocalMux I__11507 (
            .O(N__48957),
            .I(N__48949));
    Span4Mux_h I__11506 (
            .O(N__48954),
            .I(N__48946));
    Span4Mux_h I__11505 (
            .O(N__48949),
            .I(N__48943));
    Odrv4 I__11504 (
            .O(N__48946),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__11503 (
            .O(N__48943),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    CascadeMux I__11502 (
            .O(N__48938),
            .I(N__48932));
    CascadeMux I__11501 (
            .O(N__48937),
            .I(N__48927));
    InMux I__11500 (
            .O(N__48936),
            .I(N__48911));
    InMux I__11499 (
            .O(N__48935),
            .I(N__48911));
    InMux I__11498 (
            .O(N__48932),
            .I(N__48911));
    InMux I__11497 (
            .O(N__48931),
            .I(N__48911));
    InMux I__11496 (
            .O(N__48930),
            .I(N__48894));
    InMux I__11495 (
            .O(N__48927),
            .I(N__48894));
    InMux I__11494 (
            .O(N__48926),
            .I(N__48894));
    InMux I__11493 (
            .O(N__48925),
            .I(N__48881));
    InMux I__11492 (
            .O(N__48924),
            .I(N__48864));
    InMux I__11491 (
            .O(N__48923),
            .I(N__48864));
    InMux I__11490 (
            .O(N__48922),
            .I(N__48851));
    InMux I__11489 (
            .O(N__48921),
            .I(N__48846));
    InMux I__11488 (
            .O(N__48920),
            .I(N__48846));
    LocalMux I__11487 (
            .O(N__48911),
            .I(N__48843));
    InMux I__11486 (
            .O(N__48910),
            .I(N__48840));
    InMux I__11485 (
            .O(N__48909),
            .I(N__48836));
    InMux I__11484 (
            .O(N__48908),
            .I(N__48823));
    InMux I__11483 (
            .O(N__48907),
            .I(N__48820));
    InMux I__11482 (
            .O(N__48906),
            .I(N__48817));
    InMux I__11481 (
            .O(N__48905),
            .I(N__48814));
    InMux I__11480 (
            .O(N__48904),
            .I(N__48805));
    InMux I__11479 (
            .O(N__48903),
            .I(N__48805));
    InMux I__11478 (
            .O(N__48902),
            .I(N__48805));
    InMux I__11477 (
            .O(N__48901),
            .I(N__48805));
    LocalMux I__11476 (
            .O(N__48894),
            .I(N__48802));
    InMux I__11475 (
            .O(N__48893),
            .I(N__48795));
    InMux I__11474 (
            .O(N__48892),
            .I(N__48795));
    InMux I__11473 (
            .O(N__48891),
            .I(N__48795));
    InMux I__11472 (
            .O(N__48890),
            .I(N__48788));
    InMux I__11471 (
            .O(N__48889),
            .I(N__48788));
    InMux I__11470 (
            .O(N__48888),
            .I(N__48788));
    InMux I__11469 (
            .O(N__48887),
            .I(N__48779));
    InMux I__11468 (
            .O(N__48886),
            .I(N__48779));
    InMux I__11467 (
            .O(N__48885),
            .I(N__48779));
    InMux I__11466 (
            .O(N__48884),
            .I(N__48779));
    LocalMux I__11465 (
            .O(N__48881),
            .I(N__48773));
    InMux I__11464 (
            .O(N__48880),
            .I(N__48770));
    InMux I__11463 (
            .O(N__48879),
            .I(N__48765));
    InMux I__11462 (
            .O(N__48878),
            .I(N__48765));
    InMux I__11461 (
            .O(N__48877),
            .I(N__48760));
    InMux I__11460 (
            .O(N__48876),
            .I(N__48760));
    InMux I__11459 (
            .O(N__48875),
            .I(N__48752));
    InMux I__11458 (
            .O(N__48874),
            .I(N__48752));
    InMux I__11457 (
            .O(N__48873),
            .I(N__48749));
    InMux I__11456 (
            .O(N__48872),
            .I(N__48744));
    InMux I__11455 (
            .O(N__48871),
            .I(N__48744));
    InMux I__11454 (
            .O(N__48870),
            .I(N__48739));
    InMux I__11453 (
            .O(N__48869),
            .I(N__48739));
    LocalMux I__11452 (
            .O(N__48864),
            .I(N__48736));
    InMux I__11451 (
            .O(N__48863),
            .I(N__48727));
    InMux I__11450 (
            .O(N__48862),
            .I(N__48727));
    InMux I__11449 (
            .O(N__48861),
            .I(N__48727));
    InMux I__11448 (
            .O(N__48860),
            .I(N__48727));
    InMux I__11447 (
            .O(N__48859),
            .I(N__48724));
    InMux I__11446 (
            .O(N__48858),
            .I(N__48719));
    InMux I__11445 (
            .O(N__48857),
            .I(N__48719));
    InMux I__11444 (
            .O(N__48856),
            .I(N__48716));
    InMux I__11443 (
            .O(N__48855),
            .I(N__48711));
    InMux I__11442 (
            .O(N__48854),
            .I(N__48711));
    LocalMux I__11441 (
            .O(N__48851),
            .I(N__48702));
    LocalMux I__11440 (
            .O(N__48846),
            .I(N__48702));
    Span4Mux_v I__11439 (
            .O(N__48843),
            .I(N__48702));
    LocalMux I__11438 (
            .O(N__48840),
            .I(N__48702));
    InMux I__11437 (
            .O(N__48839),
            .I(N__48699));
    LocalMux I__11436 (
            .O(N__48836),
            .I(N__48696));
    InMux I__11435 (
            .O(N__48835),
            .I(N__48693));
    InMux I__11434 (
            .O(N__48834),
            .I(N__48678));
    InMux I__11433 (
            .O(N__48833),
            .I(N__48678));
    InMux I__11432 (
            .O(N__48832),
            .I(N__48678));
    InMux I__11431 (
            .O(N__48831),
            .I(N__48678));
    InMux I__11430 (
            .O(N__48830),
            .I(N__48678));
    InMux I__11429 (
            .O(N__48829),
            .I(N__48662));
    InMux I__11428 (
            .O(N__48828),
            .I(N__48657));
    InMux I__11427 (
            .O(N__48827),
            .I(N__48657));
    InMux I__11426 (
            .O(N__48826),
            .I(N__48654));
    LocalMux I__11425 (
            .O(N__48823),
            .I(N__48644));
    LocalMux I__11424 (
            .O(N__48820),
            .I(N__48644));
    LocalMux I__11423 (
            .O(N__48817),
            .I(N__48644));
    LocalMux I__11422 (
            .O(N__48814),
            .I(N__48631));
    LocalMux I__11421 (
            .O(N__48805),
            .I(N__48631));
    Span4Mux_h I__11420 (
            .O(N__48802),
            .I(N__48631));
    LocalMux I__11419 (
            .O(N__48795),
            .I(N__48631));
    LocalMux I__11418 (
            .O(N__48788),
            .I(N__48631));
    LocalMux I__11417 (
            .O(N__48779),
            .I(N__48631));
    InMux I__11416 (
            .O(N__48778),
            .I(N__48624));
    InMux I__11415 (
            .O(N__48777),
            .I(N__48624));
    InMux I__11414 (
            .O(N__48776),
            .I(N__48624));
    Span4Mux_h I__11413 (
            .O(N__48773),
            .I(N__48619));
    LocalMux I__11412 (
            .O(N__48770),
            .I(N__48619));
    LocalMux I__11411 (
            .O(N__48765),
            .I(N__48614));
    LocalMux I__11410 (
            .O(N__48760),
            .I(N__48614));
    InMux I__11409 (
            .O(N__48759),
            .I(N__48607));
    InMux I__11408 (
            .O(N__48758),
            .I(N__48607));
    InMux I__11407 (
            .O(N__48757),
            .I(N__48607));
    LocalMux I__11406 (
            .O(N__48752),
            .I(N__48590));
    LocalMux I__11405 (
            .O(N__48749),
            .I(N__48590));
    LocalMux I__11404 (
            .O(N__48744),
            .I(N__48590));
    LocalMux I__11403 (
            .O(N__48739),
            .I(N__48590));
    Span4Mux_v I__11402 (
            .O(N__48736),
            .I(N__48590));
    LocalMux I__11401 (
            .O(N__48727),
            .I(N__48590));
    LocalMux I__11400 (
            .O(N__48724),
            .I(N__48590));
    LocalMux I__11399 (
            .O(N__48719),
            .I(N__48590));
    LocalMux I__11398 (
            .O(N__48716),
            .I(N__48583));
    LocalMux I__11397 (
            .O(N__48711),
            .I(N__48583));
    Span4Mux_v I__11396 (
            .O(N__48702),
            .I(N__48583));
    LocalMux I__11395 (
            .O(N__48699),
            .I(N__48580));
    Span4Mux_v I__11394 (
            .O(N__48696),
            .I(N__48575));
    LocalMux I__11393 (
            .O(N__48693),
            .I(N__48575));
    InMux I__11392 (
            .O(N__48692),
            .I(N__48568));
    InMux I__11391 (
            .O(N__48691),
            .I(N__48568));
    InMux I__11390 (
            .O(N__48690),
            .I(N__48568));
    InMux I__11389 (
            .O(N__48689),
            .I(N__48565));
    LocalMux I__11388 (
            .O(N__48678),
            .I(N__48562));
    InMux I__11387 (
            .O(N__48677),
            .I(N__48549));
    InMux I__11386 (
            .O(N__48676),
            .I(N__48549));
    InMux I__11385 (
            .O(N__48675),
            .I(N__48549));
    InMux I__11384 (
            .O(N__48674),
            .I(N__48549));
    InMux I__11383 (
            .O(N__48673),
            .I(N__48549));
    InMux I__11382 (
            .O(N__48672),
            .I(N__48549));
    InMux I__11381 (
            .O(N__48671),
            .I(N__48540));
    InMux I__11380 (
            .O(N__48670),
            .I(N__48540));
    InMux I__11379 (
            .O(N__48669),
            .I(N__48540));
    InMux I__11378 (
            .O(N__48668),
            .I(N__48540));
    InMux I__11377 (
            .O(N__48667),
            .I(N__48533));
    InMux I__11376 (
            .O(N__48666),
            .I(N__48533));
    InMux I__11375 (
            .O(N__48665),
            .I(N__48533));
    LocalMux I__11374 (
            .O(N__48662),
            .I(N__48526));
    LocalMux I__11373 (
            .O(N__48657),
            .I(N__48526));
    LocalMux I__11372 (
            .O(N__48654),
            .I(N__48526));
    InMux I__11371 (
            .O(N__48653),
            .I(N__48519));
    InMux I__11370 (
            .O(N__48652),
            .I(N__48519));
    InMux I__11369 (
            .O(N__48651),
            .I(N__48519));
    Span4Mux_v I__11368 (
            .O(N__48644),
            .I(N__48512));
    Span4Mux_v I__11367 (
            .O(N__48631),
            .I(N__48512));
    LocalMux I__11366 (
            .O(N__48624),
            .I(N__48512));
    Span4Mux_h I__11365 (
            .O(N__48619),
            .I(N__48507));
    Span4Mux_h I__11364 (
            .O(N__48614),
            .I(N__48507));
    LocalMux I__11363 (
            .O(N__48607),
            .I(N__48500));
    Span4Mux_v I__11362 (
            .O(N__48590),
            .I(N__48500));
    Span4Mux_h I__11361 (
            .O(N__48583),
            .I(N__48500));
    Span4Mux_v I__11360 (
            .O(N__48580),
            .I(N__48495));
    Span4Mux_h I__11359 (
            .O(N__48575),
            .I(N__48495));
    LocalMux I__11358 (
            .O(N__48568),
            .I(N__48488));
    LocalMux I__11357 (
            .O(N__48565),
            .I(N__48488));
    Span12Mux_s8_h I__11356 (
            .O(N__48562),
            .I(N__48488));
    LocalMux I__11355 (
            .O(N__48549),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11354 (
            .O(N__48540),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11353 (
            .O(N__48533),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11352 (
            .O(N__48526),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11351 (
            .O(N__48519),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11350 (
            .O(N__48512),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11349 (
            .O(N__48507),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11348 (
            .O(N__48500),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11347 (
            .O(N__48495),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__11346 (
            .O(N__48488),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    InMux I__11345 (
            .O(N__48467),
            .I(N__48464));
    LocalMux I__11344 (
            .O(N__48464),
            .I(N__48459));
    InMux I__11343 (
            .O(N__48463),
            .I(N__48456));
    InMux I__11342 (
            .O(N__48462),
            .I(N__48453));
    Span4Mux_v I__11341 (
            .O(N__48459),
            .I(N__48450));
    LocalMux I__11340 (
            .O(N__48456),
            .I(N__48447));
    LocalMux I__11339 (
            .O(N__48453),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__11338 (
            .O(N__48450),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__11337 (
            .O(N__48447),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    CascadeMux I__11336 (
            .O(N__48440),
            .I(N__48432));
    InMux I__11335 (
            .O(N__48439),
            .I(N__48428));
    InMux I__11334 (
            .O(N__48438),
            .I(N__48425));
    InMux I__11333 (
            .O(N__48437),
            .I(N__48422));
    InMux I__11332 (
            .O(N__48436),
            .I(N__48419));
    InMux I__11331 (
            .O(N__48435),
            .I(N__48397));
    InMux I__11330 (
            .O(N__48432),
            .I(N__48397));
    InMux I__11329 (
            .O(N__48431),
            .I(N__48397));
    LocalMux I__11328 (
            .O(N__48428),
            .I(N__48388));
    LocalMux I__11327 (
            .O(N__48425),
            .I(N__48388));
    LocalMux I__11326 (
            .O(N__48422),
            .I(N__48388));
    LocalMux I__11325 (
            .O(N__48419),
            .I(N__48388));
    InMux I__11324 (
            .O(N__48418),
            .I(N__48381));
    InMux I__11323 (
            .O(N__48417),
            .I(N__48381));
    InMux I__11322 (
            .O(N__48416),
            .I(N__48381));
    InMux I__11321 (
            .O(N__48415),
            .I(N__48372));
    InMux I__11320 (
            .O(N__48414),
            .I(N__48372));
    InMux I__11319 (
            .O(N__48413),
            .I(N__48372));
    InMux I__11318 (
            .O(N__48412),
            .I(N__48372));
    InMux I__11317 (
            .O(N__48411),
            .I(N__48368));
    InMux I__11316 (
            .O(N__48410),
            .I(N__48363));
    InMux I__11315 (
            .O(N__48409),
            .I(N__48363));
    InMux I__11314 (
            .O(N__48408),
            .I(N__48360));
    InMux I__11313 (
            .O(N__48407),
            .I(N__48355));
    InMux I__11312 (
            .O(N__48406),
            .I(N__48355));
    InMux I__11311 (
            .O(N__48405),
            .I(N__48352));
    InMux I__11310 (
            .O(N__48404),
            .I(N__48349));
    LocalMux I__11309 (
            .O(N__48397),
            .I(N__48345));
    Span12Mux_s6_v I__11308 (
            .O(N__48388),
            .I(N__48326));
    LocalMux I__11307 (
            .O(N__48381),
            .I(N__48326));
    LocalMux I__11306 (
            .O(N__48372),
            .I(N__48326));
    InMux I__11305 (
            .O(N__48371),
            .I(N__48323));
    LocalMux I__11304 (
            .O(N__48368),
            .I(N__48312));
    LocalMux I__11303 (
            .O(N__48363),
            .I(N__48312));
    LocalMux I__11302 (
            .O(N__48360),
            .I(N__48312));
    LocalMux I__11301 (
            .O(N__48355),
            .I(N__48312));
    LocalMux I__11300 (
            .O(N__48352),
            .I(N__48312));
    LocalMux I__11299 (
            .O(N__48349),
            .I(N__48309));
    InMux I__11298 (
            .O(N__48348),
            .I(N__48306));
    Span4Mux_h I__11297 (
            .O(N__48345),
            .I(N__48296));
    CascadeMux I__11296 (
            .O(N__48344),
            .I(N__48292));
    CascadeMux I__11295 (
            .O(N__48343),
            .I(N__48288));
    CascadeMux I__11294 (
            .O(N__48342),
            .I(N__48284));
    CascadeMux I__11293 (
            .O(N__48341),
            .I(N__48280));
    CascadeMux I__11292 (
            .O(N__48340),
            .I(N__48276));
    CascadeMux I__11291 (
            .O(N__48339),
            .I(N__48272));
    CascadeMux I__11290 (
            .O(N__48338),
            .I(N__48268));
    CascadeMux I__11289 (
            .O(N__48337),
            .I(N__48264));
    CascadeMux I__11288 (
            .O(N__48336),
            .I(N__48260));
    CascadeMux I__11287 (
            .O(N__48335),
            .I(N__48256));
    CascadeMux I__11286 (
            .O(N__48334),
            .I(N__48252));
    InMux I__11285 (
            .O(N__48333),
            .I(N__48245));
    Span12Mux_v I__11284 (
            .O(N__48326),
            .I(N__48238));
    LocalMux I__11283 (
            .O(N__48323),
            .I(N__48238));
    Span12Mux_s11_v I__11282 (
            .O(N__48312),
            .I(N__48238));
    Span4Mux_s1_h I__11281 (
            .O(N__48309),
            .I(N__48235));
    LocalMux I__11280 (
            .O(N__48306),
            .I(N__48232));
    InMux I__11279 (
            .O(N__48305),
            .I(N__48225));
    InMux I__11278 (
            .O(N__48304),
            .I(N__48225));
    InMux I__11277 (
            .O(N__48303),
            .I(N__48225));
    InMux I__11276 (
            .O(N__48302),
            .I(N__48216));
    InMux I__11275 (
            .O(N__48301),
            .I(N__48216));
    InMux I__11274 (
            .O(N__48300),
            .I(N__48216));
    InMux I__11273 (
            .O(N__48299),
            .I(N__48216));
    Span4Mux_h I__11272 (
            .O(N__48296),
            .I(N__48213));
    InMux I__11271 (
            .O(N__48295),
            .I(N__48198));
    InMux I__11270 (
            .O(N__48292),
            .I(N__48198));
    InMux I__11269 (
            .O(N__48291),
            .I(N__48198));
    InMux I__11268 (
            .O(N__48288),
            .I(N__48198));
    InMux I__11267 (
            .O(N__48287),
            .I(N__48198));
    InMux I__11266 (
            .O(N__48284),
            .I(N__48198));
    InMux I__11265 (
            .O(N__48283),
            .I(N__48198));
    InMux I__11264 (
            .O(N__48280),
            .I(N__48181));
    InMux I__11263 (
            .O(N__48279),
            .I(N__48181));
    InMux I__11262 (
            .O(N__48276),
            .I(N__48181));
    InMux I__11261 (
            .O(N__48275),
            .I(N__48181));
    InMux I__11260 (
            .O(N__48272),
            .I(N__48181));
    InMux I__11259 (
            .O(N__48271),
            .I(N__48181));
    InMux I__11258 (
            .O(N__48268),
            .I(N__48181));
    InMux I__11257 (
            .O(N__48267),
            .I(N__48181));
    InMux I__11256 (
            .O(N__48264),
            .I(N__48164));
    InMux I__11255 (
            .O(N__48263),
            .I(N__48164));
    InMux I__11254 (
            .O(N__48260),
            .I(N__48164));
    InMux I__11253 (
            .O(N__48259),
            .I(N__48164));
    InMux I__11252 (
            .O(N__48256),
            .I(N__48164));
    InMux I__11251 (
            .O(N__48255),
            .I(N__48164));
    InMux I__11250 (
            .O(N__48252),
            .I(N__48164));
    InMux I__11249 (
            .O(N__48251),
            .I(N__48164));
    CascadeMux I__11248 (
            .O(N__48250),
            .I(N__48160));
    CascadeMux I__11247 (
            .O(N__48249),
            .I(N__48156));
    CascadeMux I__11246 (
            .O(N__48248),
            .I(N__48152));
    LocalMux I__11245 (
            .O(N__48245),
            .I(N__48147));
    Span12Mux_h I__11244 (
            .O(N__48238),
            .I(N__48144));
    Span4Mux_v I__11243 (
            .O(N__48235),
            .I(N__48139));
    Span4Mux_s1_h I__11242 (
            .O(N__48232),
            .I(N__48139));
    LocalMux I__11241 (
            .O(N__48225),
            .I(N__48134));
    LocalMux I__11240 (
            .O(N__48216),
            .I(N__48134));
    Sp12to4 I__11239 (
            .O(N__48213),
            .I(N__48129));
    LocalMux I__11238 (
            .O(N__48198),
            .I(N__48129));
    LocalMux I__11237 (
            .O(N__48181),
            .I(N__48126));
    LocalMux I__11236 (
            .O(N__48164),
            .I(N__48123));
    InMux I__11235 (
            .O(N__48163),
            .I(N__48108));
    InMux I__11234 (
            .O(N__48160),
            .I(N__48108));
    InMux I__11233 (
            .O(N__48159),
            .I(N__48108));
    InMux I__11232 (
            .O(N__48156),
            .I(N__48108));
    InMux I__11231 (
            .O(N__48155),
            .I(N__48108));
    InMux I__11230 (
            .O(N__48152),
            .I(N__48108));
    InMux I__11229 (
            .O(N__48151),
            .I(N__48108));
    InMux I__11228 (
            .O(N__48150),
            .I(N__48105));
    Span4Mux_v I__11227 (
            .O(N__48147),
            .I(N__48102));
    Span12Mux_h I__11226 (
            .O(N__48144),
            .I(N__48095));
    Sp12to4 I__11225 (
            .O(N__48139),
            .I(N__48095));
    Span12Mux_s1_h I__11224 (
            .O(N__48134),
            .I(N__48095));
    Span12Mux_s9_v I__11223 (
            .O(N__48129),
            .I(N__48084));
    Sp12to4 I__11222 (
            .O(N__48126),
            .I(N__48084));
    Span12Mux_s8_h I__11221 (
            .O(N__48123),
            .I(N__48084));
    LocalMux I__11220 (
            .O(N__48108),
            .I(N__48084));
    LocalMux I__11219 (
            .O(N__48105),
            .I(N__48084));
    Span4Mux_v I__11218 (
            .O(N__48102),
            .I(N__48081));
    Span12Mux_v I__11217 (
            .O(N__48095),
            .I(N__48078));
    Span12Mux_v I__11216 (
            .O(N__48084),
            .I(N__48075));
    Span4Mux_h I__11215 (
            .O(N__48081),
            .I(N__48072));
    Odrv12 I__11214 (
            .O(N__48078),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__11213 (
            .O(N__48075),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__11212 (
            .O(N__48072),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__11211 (
            .O(N__48065),
            .I(N__48060));
    InMux I__11210 (
            .O(N__48064),
            .I(N__48057));
    InMux I__11209 (
            .O(N__48063),
            .I(N__48054));
    InMux I__11208 (
            .O(N__48060),
            .I(N__48051));
    LocalMux I__11207 (
            .O(N__48057),
            .I(N__48048));
    LocalMux I__11206 (
            .O(N__48054),
            .I(N__48044));
    LocalMux I__11205 (
            .O(N__48051),
            .I(N__48041));
    Span4Mux_h I__11204 (
            .O(N__48048),
            .I(N__48038));
    InMux I__11203 (
            .O(N__48047),
            .I(N__48035));
    Span12Mux_h I__11202 (
            .O(N__48044),
            .I(N__48032));
    Span4Mux_v I__11201 (
            .O(N__48041),
            .I(N__48027));
    Span4Mux_h I__11200 (
            .O(N__48038),
            .I(N__48027));
    LocalMux I__11199 (
            .O(N__48035),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv12 I__11198 (
            .O(N__48032),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__11197 (
            .O(N__48027),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__11196 (
            .O(N__48020),
            .I(N__48017));
    LocalMux I__11195 (
            .O(N__48017),
            .I(N__48014));
    Span4Mux_h I__11194 (
            .O(N__48014),
            .I(N__48010));
    InMux I__11193 (
            .O(N__48013),
            .I(N__48007));
    Span4Mux_h I__11192 (
            .O(N__48010),
            .I(N__48004));
    LocalMux I__11191 (
            .O(N__48007),
            .I(N__48001));
    Span4Mux_v I__11190 (
            .O(N__48004),
            .I(N__47997));
    Span4Mux_h I__11189 (
            .O(N__48001),
            .I(N__47993));
    InMux I__11188 (
            .O(N__48000),
            .I(N__47990));
    Span4Mux_v I__11187 (
            .O(N__47997),
            .I(N__47987));
    InMux I__11186 (
            .O(N__47996),
            .I(N__47984));
    Span4Mux_h I__11185 (
            .O(N__47993),
            .I(N__47981));
    LocalMux I__11184 (
            .O(N__47990),
            .I(N__47978));
    Odrv4 I__11183 (
            .O(N__47987),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__11182 (
            .O(N__47984),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__11181 (
            .O(N__47981),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv12 I__11180 (
            .O(N__47978),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__11179 (
            .O(N__47969),
            .I(N__47966));
    LocalMux I__11178 (
            .O(N__47966),
            .I(N__47963));
    Span4Mux_v I__11177 (
            .O(N__47963),
            .I(N__47959));
    InMux I__11176 (
            .O(N__47962),
            .I(N__47956));
    Span4Mux_h I__11175 (
            .O(N__47959),
            .I(N__47953));
    LocalMux I__11174 (
            .O(N__47956),
            .I(N__47950));
    Odrv4 I__11173 (
            .O(N__47953),
            .I(\phase_controller_inst1.state_RNIE87FZ0Z_2 ));
    Odrv12 I__11172 (
            .O(N__47950),
            .I(\phase_controller_inst1.state_RNIE87FZ0Z_2 ));
    InMux I__11171 (
            .O(N__47945),
            .I(N__47940));
    InMux I__11170 (
            .O(N__47944),
            .I(N__47937));
    InMux I__11169 (
            .O(N__47943),
            .I(N__47934));
    LocalMux I__11168 (
            .O(N__47940),
            .I(N__47931));
    LocalMux I__11167 (
            .O(N__47937),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    LocalMux I__11166 (
            .O(N__47934),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    Odrv4 I__11165 (
            .O(N__47931),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    InMux I__11164 (
            .O(N__47924),
            .I(N__47919));
    InMux I__11163 (
            .O(N__47923),
            .I(N__47916));
    InMux I__11162 (
            .O(N__47922),
            .I(N__47913));
    LocalMux I__11161 (
            .O(N__47919),
            .I(N__47908));
    LocalMux I__11160 (
            .O(N__47916),
            .I(N__47908));
    LocalMux I__11159 (
            .O(N__47913),
            .I(N__47904));
    Span4Mux_h I__11158 (
            .O(N__47908),
            .I(N__47901));
    InMux I__11157 (
            .O(N__47907),
            .I(N__47898));
    Odrv12 I__11156 (
            .O(N__47904),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    Odrv4 I__11155 (
            .O(N__47901),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    LocalMux I__11154 (
            .O(N__47898),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__11153 (
            .O(N__47891),
            .I(N__47885));
    InMux I__11152 (
            .O(N__47890),
            .I(N__47885));
    LocalMux I__11151 (
            .O(N__47885),
            .I(N__47882));
    Span4Mux_h I__11150 (
            .O(N__47882),
            .I(N__47879));
    Span4Mux_h I__11149 (
            .O(N__47879),
            .I(N__47876));
    Odrv4 I__11148 (
            .O(N__47876),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    CEMux I__11147 (
            .O(N__47873),
            .I(N__47831));
    CEMux I__11146 (
            .O(N__47872),
            .I(N__47831));
    CEMux I__11145 (
            .O(N__47871),
            .I(N__47831));
    CEMux I__11144 (
            .O(N__47870),
            .I(N__47831));
    CEMux I__11143 (
            .O(N__47869),
            .I(N__47831));
    CEMux I__11142 (
            .O(N__47868),
            .I(N__47831));
    CEMux I__11141 (
            .O(N__47867),
            .I(N__47831));
    CEMux I__11140 (
            .O(N__47866),
            .I(N__47831));
    CEMux I__11139 (
            .O(N__47865),
            .I(N__47831));
    CEMux I__11138 (
            .O(N__47864),
            .I(N__47831));
    CEMux I__11137 (
            .O(N__47863),
            .I(N__47831));
    CEMux I__11136 (
            .O(N__47862),
            .I(N__47831));
    CEMux I__11135 (
            .O(N__47861),
            .I(N__47831));
    CEMux I__11134 (
            .O(N__47860),
            .I(N__47831));
    GlobalMux I__11133 (
            .O(N__47831),
            .I(N__47828));
    gio2CtrlBuf I__11132 (
            .O(N__47828),
            .I(\phase_controller_inst2.stoper_hc.un1_start_g ));
    InMux I__11131 (
            .O(N__47825),
            .I(N__47820));
    InMux I__11130 (
            .O(N__47824),
            .I(N__47817));
    InMux I__11129 (
            .O(N__47823),
            .I(N__47814));
    LocalMux I__11128 (
            .O(N__47820),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    LocalMux I__11127 (
            .O(N__47817),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    LocalMux I__11126 (
            .O(N__47814),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    InMux I__11125 (
            .O(N__47807),
            .I(N__47804));
    LocalMux I__11124 (
            .O(N__47804),
            .I(N__47799));
    InMux I__11123 (
            .O(N__47803),
            .I(N__47796));
    InMux I__11122 (
            .O(N__47802),
            .I(N__47793));
    Span4Mux_v I__11121 (
            .O(N__47799),
            .I(N__47789));
    LocalMux I__11120 (
            .O(N__47796),
            .I(N__47784));
    LocalMux I__11119 (
            .O(N__47793),
            .I(N__47784));
    CascadeMux I__11118 (
            .O(N__47792),
            .I(N__47781));
    Span4Mux_h I__11117 (
            .O(N__47789),
            .I(N__47778));
    Span4Mux_v I__11116 (
            .O(N__47784),
            .I(N__47775));
    InMux I__11115 (
            .O(N__47781),
            .I(N__47772));
    Odrv4 I__11114 (
            .O(N__47778),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__11113 (
            .O(N__47775),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    LocalMux I__11112 (
            .O(N__47772),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__11111 (
            .O(N__47765),
            .I(N__47759));
    InMux I__11110 (
            .O(N__47764),
            .I(N__47759));
    LocalMux I__11109 (
            .O(N__47759),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__11108 (
            .O(N__47756),
            .I(N__47753));
    LocalMux I__11107 (
            .O(N__47753),
            .I(N__47750));
    Span4Mux_h I__11106 (
            .O(N__47750),
            .I(N__47745));
    InMux I__11105 (
            .O(N__47749),
            .I(N__47742));
    InMux I__11104 (
            .O(N__47748),
            .I(N__47739));
    Span4Mux_h I__11103 (
            .O(N__47745),
            .I(N__47734));
    LocalMux I__11102 (
            .O(N__47742),
            .I(N__47734));
    LocalMux I__11101 (
            .O(N__47739),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    Odrv4 I__11100 (
            .O(N__47734),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    InMux I__11099 (
            .O(N__47729),
            .I(N__47724));
    InMux I__11098 (
            .O(N__47728),
            .I(N__47721));
    InMux I__11097 (
            .O(N__47727),
            .I(N__47717));
    LocalMux I__11096 (
            .O(N__47724),
            .I(N__47714));
    LocalMux I__11095 (
            .O(N__47721),
            .I(N__47711));
    InMux I__11094 (
            .O(N__47720),
            .I(N__47708));
    LocalMux I__11093 (
            .O(N__47717),
            .I(N__47705));
    Span4Mux_h I__11092 (
            .O(N__47714),
            .I(N__47700));
    Span4Mux_v I__11091 (
            .O(N__47711),
            .I(N__47700));
    LocalMux I__11090 (
            .O(N__47708),
            .I(N__47697));
    Odrv12 I__11089 (
            .O(N__47705),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    Odrv4 I__11088 (
            .O(N__47700),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    Odrv4 I__11087 (
            .O(N__47697),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    CascadeMux I__11086 (
            .O(N__47690),
            .I(N__47687));
    InMux I__11085 (
            .O(N__47687),
            .I(N__47684));
    LocalMux I__11084 (
            .O(N__47684),
            .I(N__47681));
    Span4Mux_h I__11083 (
            .O(N__47681),
            .I(N__47678));
    Odrv4 I__11082 (
            .O(N__47678),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt22 ));
    InMux I__11081 (
            .O(N__47675),
            .I(N__47672));
    LocalMux I__11080 (
            .O(N__47672),
            .I(N__47669));
    Span12Mux_h I__11079 (
            .O(N__47669),
            .I(N__47665));
    InMux I__11078 (
            .O(N__47668),
            .I(N__47662));
    Odrv12 I__11077 (
            .O(N__47665),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    LocalMux I__11076 (
            .O(N__47662),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    InMux I__11075 (
            .O(N__47657),
            .I(N__47650));
    InMux I__11074 (
            .O(N__47656),
            .I(N__47650));
    InMux I__11073 (
            .O(N__47655),
            .I(N__47647));
    LocalMux I__11072 (
            .O(N__47650),
            .I(N__47644));
    LocalMux I__11071 (
            .O(N__47647),
            .I(N__47640));
    Span4Mux_v I__11070 (
            .O(N__47644),
            .I(N__47637));
    InMux I__11069 (
            .O(N__47643),
            .I(N__47634));
    Span4Mux_v I__11068 (
            .O(N__47640),
            .I(N__47629));
    Span4Mux_h I__11067 (
            .O(N__47637),
            .I(N__47629));
    LocalMux I__11066 (
            .O(N__47634),
            .I(N__47626));
    Odrv4 I__11065 (
            .O(N__47629),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv4 I__11064 (
            .O(N__47626),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    CascadeMux I__11063 (
            .O(N__47621),
            .I(elapsed_time_ns_1_RNI14DN9_0_23_cascade_));
    InMux I__11062 (
            .O(N__47618),
            .I(N__47612));
    InMux I__11061 (
            .O(N__47617),
            .I(N__47612));
    LocalMux I__11060 (
            .O(N__47612),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ));
    InMux I__11059 (
            .O(N__47609),
            .I(N__47603));
    InMux I__11058 (
            .O(N__47608),
            .I(N__47603));
    LocalMux I__11057 (
            .O(N__47603),
            .I(N__47599));
    InMux I__11056 (
            .O(N__47602),
            .I(N__47596));
    Span4Mux_h I__11055 (
            .O(N__47599),
            .I(N__47593));
    LocalMux I__11054 (
            .O(N__47596),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__11053 (
            .O(N__47593),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    CascadeMux I__11052 (
            .O(N__47588),
            .I(N__47584));
    CascadeMux I__11051 (
            .O(N__47587),
            .I(N__47581));
    InMux I__11050 (
            .O(N__47584),
            .I(N__47576));
    InMux I__11049 (
            .O(N__47581),
            .I(N__47576));
    LocalMux I__11048 (
            .O(N__47576),
            .I(N__47572));
    InMux I__11047 (
            .O(N__47575),
            .I(N__47569));
    Span4Mux_h I__11046 (
            .O(N__47572),
            .I(N__47566));
    LocalMux I__11045 (
            .O(N__47569),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__11044 (
            .O(N__47566),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__11043 (
            .O(N__47561),
            .I(N__47555));
    InMux I__11042 (
            .O(N__47560),
            .I(N__47555));
    LocalMux I__11041 (
            .O(N__47555),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ));
    InMux I__11040 (
            .O(N__47552),
            .I(N__47549));
    LocalMux I__11039 (
            .O(N__47549),
            .I(N__47546));
    Odrv12 I__11038 (
            .O(N__47546),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ));
    InMux I__11037 (
            .O(N__47543),
            .I(N__47540));
    LocalMux I__11036 (
            .O(N__47540),
            .I(N__47537));
    Span4Mux_h I__11035 (
            .O(N__47537),
            .I(N__47534));
    Span4Mux_h I__11034 (
            .O(N__47534),
            .I(N__47530));
    InMux I__11033 (
            .O(N__47533),
            .I(N__47527));
    Odrv4 I__11032 (
            .O(N__47530),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    LocalMux I__11031 (
            .O(N__47527),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    InMux I__11030 (
            .O(N__47522),
            .I(N__47515));
    InMux I__11029 (
            .O(N__47521),
            .I(N__47515));
    InMux I__11028 (
            .O(N__47520),
            .I(N__47512));
    LocalMux I__11027 (
            .O(N__47515),
            .I(N__47509));
    LocalMux I__11026 (
            .O(N__47512),
            .I(N__47505));
    Span12Mux_v I__11025 (
            .O(N__47509),
            .I(N__47502));
    InMux I__11024 (
            .O(N__47508),
            .I(N__47499));
    Odrv4 I__11023 (
            .O(N__47505),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv12 I__11022 (
            .O(N__47502),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    LocalMux I__11021 (
            .O(N__47499),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    CascadeMux I__11020 (
            .O(N__47492),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_));
    InMux I__11019 (
            .O(N__47489),
            .I(N__47486));
    LocalMux I__11018 (
            .O(N__47486),
            .I(N__47483));
    Span4Mux_h I__11017 (
            .O(N__47483),
            .I(N__47480));
    Odrv4 I__11016 (
            .O(N__47480),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__11015 (
            .O(N__47477),
            .I(N__47472));
    InMux I__11014 (
            .O(N__47476),
            .I(N__47469));
    InMux I__11013 (
            .O(N__47475),
            .I(N__47466));
    LocalMux I__11012 (
            .O(N__47472),
            .I(N__47461));
    LocalMux I__11011 (
            .O(N__47469),
            .I(N__47461));
    LocalMux I__11010 (
            .O(N__47466),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    Odrv12 I__11009 (
            .O(N__47461),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    InMux I__11008 (
            .O(N__47456),
            .I(N__47452));
    InMux I__11007 (
            .O(N__47455),
            .I(N__47449));
    LocalMux I__11006 (
            .O(N__47452),
            .I(N__47444));
    LocalMux I__11005 (
            .O(N__47449),
            .I(N__47441));
    InMux I__11004 (
            .O(N__47448),
            .I(N__47438));
    InMux I__11003 (
            .O(N__47447),
            .I(N__47435));
    Span4Mux_v I__11002 (
            .O(N__47444),
            .I(N__47430));
    Span4Mux_v I__11001 (
            .O(N__47441),
            .I(N__47430));
    LocalMux I__11000 (
            .O(N__47438),
            .I(N__47427));
    LocalMux I__10999 (
            .O(N__47435),
            .I(N__47424));
    Span4Mux_h I__10998 (
            .O(N__47430),
            .I(N__47419));
    Span4Mux_h I__10997 (
            .O(N__47427),
            .I(N__47419));
    Span4Mux_h I__10996 (
            .O(N__47424),
            .I(N__47416));
    Sp12to4 I__10995 (
            .O(N__47419),
            .I(N__47413));
    Odrv4 I__10994 (
            .O(N__47416),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    Odrv12 I__10993 (
            .O(N__47413),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__10992 (
            .O(N__47408),
            .I(N__47405));
    LocalMux I__10991 (
            .O(N__47405),
            .I(N__47402));
    Span4Mux_h I__10990 (
            .O(N__47402),
            .I(N__47399));
    Odrv4 I__10989 (
            .O(N__47399),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ));
    InMux I__10988 (
            .O(N__47396),
            .I(N__47389));
    InMux I__10987 (
            .O(N__47395),
            .I(N__47389));
    InMux I__10986 (
            .O(N__47394),
            .I(N__47386));
    LocalMux I__10985 (
            .O(N__47389),
            .I(N__47383));
    LocalMux I__10984 (
            .O(N__47386),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv4 I__10983 (
            .O(N__47383),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    CascadeMux I__10982 (
            .O(N__47378),
            .I(N__47375));
    InMux I__10981 (
            .O(N__47375),
            .I(N__47368));
    InMux I__10980 (
            .O(N__47374),
            .I(N__47368));
    InMux I__10979 (
            .O(N__47373),
            .I(N__47365));
    LocalMux I__10978 (
            .O(N__47368),
            .I(N__47362));
    LocalMux I__10977 (
            .O(N__47365),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv4 I__10976 (
            .O(N__47362),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    CascadeMux I__10975 (
            .O(N__47357),
            .I(N__47354));
    InMux I__10974 (
            .O(N__47354),
            .I(N__47348));
    InMux I__10973 (
            .O(N__47353),
            .I(N__47348));
    LocalMux I__10972 (
            .O(N__47348),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ));
    CascadeMux I__10971 (
            .O(N__47345),
            .I(N__47342));
    InMux I__10970 (
            .O(N__47342),
            .I(N__47339));
    LocalMux I__10969 (
            .O(N__47339),
            .I(N__47336));
    Span4Mux_h I__10968 (
            .O(N__47336),
            .I(N__47333));
    Odrv4 I__10967 (
            .O(N__47333),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt28 ));
    InMux I__10966 (
            .O(N__47330),
            .I(N__47327));
    LocalMux I__10965 (
            .O(N__47327),
            .I(N__47324));
    Span4Mux_h I__10964 (
            .O(N__47324),
            .I(N__47320));
    InMux I__10963 (
            .O(N__47323),
            .I(N__47317));
    Odrv4 I__10962 (
            .O(N__47320),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    LocalMux I__10961 (
            .O(N__47317),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    InMux I__10960 (
            .O(N__47312),
            .I(N__47306));
    InMux I__10959 (
            .O(N__47311),
            .I(N__47306));
    LocalMux I__10958 (
            .O(N__47306),
            .I(N__47302));
    InMux I__10957 (
            .O(N__47305),
            .I(N__47298));
    Span4Mux_v I__10956 (
            .O(N__47302),
            .I(N__47295));
    InMux I__10955 (
            .O(N__47301),
            .I(N__47292));
    LocalMux I__10954 (
            .O(N__47298),
            .I(N__47289));
    Span4Mux_v I__10953 (
            .O(N__47295),
            .I(N__47284));
    LocalMux I__10952 (
            .O(N__47292),
            .I(N__47284));
    Span4Mux_v I__10951 (
            .O(N__47289),
            .I(N__47281));
    Span4Mux_h I__10950 (
            .O(N__47284),
            .I(N__47278));
    Odrv4 I__10949 (
            .O(N__47281),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    Odrv4 I__10948 (
            .O(N__47278),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    CascadeMux I__10947 (
            .O(N__47273),
            .I(elapsed_time_ns_1_RNI69DN9_0_28_cascade_));
    InMux I__10946 (
            .O(N__47270),
            .I(N__47264));
    InMux I__10945 (
            .O(N__47269),
            .I(N__47264));
    LocalMux I__10944 (
            .O(N__47264),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ));
    InMux I__10943 (
            .O(N__47261),
            .I(N__47255));
    InMux I__10942 (
            .O(N__47260),
            .I(N__47255));
    LocalMux I__10941 (
            .O(N__47255),
            .I(N__47252));
    Odrv4 I__10940 (
            .O(N__47252),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    InMux I__10939 (
            .O(N__47249),
            .I(N__47245));
    InMux I__10938 (
            .O(N__47248),
            .I(N__47242));
    LocalMux I__10937 (
            .O(N__47245),
            .I(N__47237));
    LocalMux I__10936 (
            .O(N__47242),
            .I(N__47237));
    Odrv4 I__10935 (
            .O(N__47237),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    InMux I__10934 (
            .O(N__47234),
            .I(N__47231));
    LocalMux I__10933 (
            .O(N__47231),
            .I(N__47228));
    Span4Mux_h I__10932 (
            .O(N__47228),
            .I(N__47224));
    InMux I__10931 (
            .O(N__47227),
            .I(N__47221));
    Odrv4 I__10930 (
            .O(N__47224),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    LocalMux I__10929 (
            .O(N__47221),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    InMux I__10928 (
            .O(N__47216),
            .I(N__47210));
    InMux I__10927 (
            .O(N__47215),
            .I(N__47210));
    LocalMux I__10926 (
            .O(N__47210),
            .I(N__47206));
    InMux I__10925 (
            .O(N__47209),
            .I(N__47203));
    Span4Mux_h I__10924 (
            .O(N__47206),
            .I(N__47200));
    LocalMux I__10923 (
            .O(N__47203),
            .I(N__47196));
    Span4Mux_h I__10922 (
            .O(N__47200),
            .I(N__47193));
    InMux I__10921 (
            .O(N__47199),
            .I(N__47190));
    Odrv4 I__10920 (
            .O(N__47196),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv4 I__10919 (
            .O(N__47193),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    LocalMux I__10918 (
            .O(N__47190),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    CascadeMux I__10917 (
            .O(N__47183),
            .I(elapsed_time_ns_1_RNI46CN9_0_17_cascade_));
    InMux I__10916 (
            .O(N__47180),
            .I(N__47175));
    InMux I__10915 (
            .O(N__47179),
            .I(N__47170));
    InMux I__10914 (
            .O(N__47178),
            .I(N__47170));
    LocalMux I__10913 (
            .O(N__47175),
            .I(N__47165));
    LocalMux I__10912 (
            .O(N__47170),
            .I(N__47165));
    Odrv4 I__10911 (
            .O(N__47165),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__10910 (
            .O(N__47162),
            .I(N__47158));
    CascadeMux I__10909 (
            .O(N__47161),
            .I(N__47155));
    InMux I__10908 (
            .O(N__47158),
            .I(N__47150));
    InMux I__10907 (
            .O(N__47155),
            .I(N__47150));
    LocalMux I__10906 (
            .O(N__47150),
            .I(N__47146));
    InMux I__10905 (
            .O(N__47149),
            .I(N__47143));
    Span4Mux_v I__10904 (
            .O(N__47146),
            .I(N__47140));
    LocalMux I__10903 (
            .O(N__47143),
            .I(N__47135));
    Span4Mux_h I__10902 (
            .O(N__47140),
            .I(N__47135));
    Odrv4 I__10901 (
            .O(N__47135),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__10900 (
            .O(N__47132),
            .I(N__47126));
    InMux I__10899 (
            .O(N__47131),
            .I(N__47126));
    LocalMux I__10898 (
            .O(N__47126),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__10897 (
            .O(N__47123),
            .I(N__47120));
    LocalMux I__10896 (
            .O(N__47120),
            .I(N__47117));
    Span4Mux_h I__10895 (
            .O(N__47117),
            .I(N__47114));
    Odrv4 I__10894 (
            .O(N__47114),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    InMux I__10893 (
            .O(N__47111),
            .I(N__47108));
    LocalMux I__10892 (
            .O(N__47108),
            .I(N__47104));
    InMux I__10891 (
            .O(N__47107),
            .I(N__47101));
    Span4Mux_v I__10890 (
            .O(N__47104),
            .I(N__47098));
    LocalMux I__10889 (
            .O(N__47101),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    Odrv4 I__10888 (
            .O(N__47098),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    InMux I__10887 (
            .O(N__47093),
            .I(N__47086));
    InMux I__10886 (
            .O(N__47092),
            .I(N__47086));
    InMux I__10885 (
            .O(N__47091),
            .I(N__47083));
    LocalMux I__10884 (
            .O(N__47086),
            .I(N__47080));
    LocalMux I__10883 (
            .O(N__47083),
            .I(N__47076));
    Span4Mux_v I__10882 (
            .O(N__47080),
            .I(N__47073));
    InMux I__10881 (
            .O(N__47079),
            .I(N__47070));
    Odrv4 I__10880 (
            .O(N__47076),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    Odrv4 I__10879 (
            .O(N__47073),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    LocalMux I__10878 (
            .O(N__47070),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    CascadeMux I__10877 (
            .O(N__47063),
            .I(elapsed_time_ns_1_RNI13CN9_0_14_cascade_));
    InMux I__10876 (
            .O(N__47060),
            .I(N__47057));
    LocalMux I__10875 (
            .O(N__47057),
            .I(N__47054));
    Span4Mux_h I__10874 (
            .O(N__47054),
            .I(N__47051));
    Odrv4 I__10873 (
            .O(N__47051),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__10872 (
            .O(N__47048),
            .I(N__47042));
    InMux I__10871 (
            .O(N__47047),
            .I(N__47042));
    LocalMux I__10870 (
            .O(N__47042),
            .I(N__47039));
    Odrv12 I__10869 (
            .O(N__47039),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__10868 (
            .O(N__47036),
            .I(N__47033));
    InMux I__10867 (
            .O(N__47033),
            .I(N__47027));
    InMux I__10866 (
            .O(N__47032),
            .I(N__47027));
    LocalMux I__10865 (
            .O(N__47027),
            .I(N__47024));
    Span4Mux_h I__10864 (
            .O(N__47024),
            .I(N__47021));
    Odrv4 I__10863 (
            .O(N__47021),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ));
    InMux I__10862 (
            .O(N__47018),
            .I(N__47015));
    LocalMux I__10861 (
            .O(N__47015),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ));
    InMux I__10860 (
            .O(N__47012),
            .I(N__47009));
    LocalMux I__10859 (
            .O(N__47009),
            .I(N__47006));
    Odrv12 I__10858 (
            .O(N__47006),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    InMux I__10857 (
            .O(N__47003),
            .I(N__46999));
    InMux I__10856 (
            .O(N__47002),
            .I(N__46996));
    LocalMux I__10855 (
            .O(N__46999),
            .I(N__46993));
    LocalMux I__10854 (
            .O(N__46996),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    Odrv4 I__10853 (
            .O(N__46993),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    InMux I__10852 (
            .O(N__46988),
            .I(N__46982));
    InMux I__10851 (
            .O(N__46987),
            .I(N__46974));
    InMux I__10850 (
            .O(N__46986),
            .I(N__46974));
    InMux I__10849 (
            .O(N__46985),
            .I(N__46974));
    LocalMux I__10848 (
            .O(N__46982),
            .I(N__46971));
    InMux I__10847 (
            .O(N__46981),
            .I(N__46968));
    LocalMux I__10846 (
            .O(N__46974),
            .I(N__46965));
    Odrv12 I__10845 (
            .O(N__46971),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__10844 (
            .O(N__46968),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__10843 (
            .O(N__46965),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    InMux I__10842 (
            .O(N__46958),
            .I(N__46954));
    CascadeMux I__10841 (
            .O(N__46957),
            .I(N__46951));
    LocalMux I__10840 (
            .O(N__46954),
            .I(N__46947));
    InMux I__10839 (
            .O(N__46951),
            .I(N__46942));
    InMux I__10838 (
            .O(N__46950),
            .I(N__46942));
    Span4Mux_h I__10837 (
            .O(N__46947),
            .I(N__46939));
    LocalMux I__10836 (
            .O(N__46942),
            .I(N__46936));
    Odrv4 I__10835 (
            .O(N__46939),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv4 I__10834 (
            .O(N__46936),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    CascadeMux I__10833 (
            .O(N__46931),
            .I(N__46927));
    InMux I__10832 (
            .O(N__46930),
            .I(N__46923));
    InMux I__10831 (
            .O(N__46927),
            .I(N__46920));
    InMux I__10830 (
            .O(N__46926),
            .I(N__46917));
    LocalMux I__10829 (
            .O(N__46923),
            .I(N__46913));
    LocalMux I__10828 (
            .O(N__46920),
            .I(N__46910));
    LocalMux I__10827 (
            .O(N__46917),
            .I(N__46907));
    CascadeMux I__10826 (
            .O(N__46916),
            .I(N__46904));
    Span4Mux_h I__10825 (
            .O(N__46913),
            .I(N__46901));
    Span4Mux_v I__10824 (
            .O(N__46910),
            .I(N__46896));
    Span4Mux_h I__10823 (
            .O(N__46907),
            .I(N__46896));
    InMux I__10822 (
            .O(N__46904),
            .I(N__46891));
    Span4Mux_h I__10821 (
            .O(N__46901),
            .I(N__46888));
    Span4Mux_h I__10820 (
            .O(N__46896),
            .I(N__46885));
    InMux I__10819 (
            .O(N__46895),
            .I(N__46880));
    InMux I__10818 (
            .O(N__46894),
            .I(N__46880));
    LocalMux I__10817 (
            .O(N__46891),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__10816 (
            .O(N__46888),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__10815 (
            .O(N__46885),
            .I(phase_controller_inst1_state_4));
    LocalMux I__10814 (
            .O(N__46880),
            .I(phase_controller_inst1_state_4));
    InMux I__10813 (
            .O(N__46871),
            .I(N__46868));
    LocalMux I__10812 (
            .O(N__46868),
            .I(N__46865));
    Span4Mux_v I__10811 (
            .O(N__46865),
            .I(N__46862));
    Span4Mux_h I__10810 (
            .O(N__46862),
            .I(N__46859));
    Odrv4 I__10809 (
            .O(N__46859),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    CascadeMux I__10808 (
            .O(N__46856),
            .I(N__46853));
    InMux I__10807 (
            .O(N__46853),
            .I(N__46845));
    InMux I__10806 (
            .O(N__46852),
            .I(N__46845));
    InMux I__10805 (
            .O(N__46851),
            .I(N__46840));
    InMux I__10804 (
            .O(N__46850),
            .I(N__46840));
    LocalMux I__10803 (
            .O(N__46845),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__10802 (
            .O(N__46840),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__10801 (
            .O(N__46835),
            .I(N__46828));
    InMux I__10800 (
            .O(N__46834),
            .I(N__46828));
    CascadeMux I__10799 (
            .O(N__46833),
            .I(N__46825));
    LocalMux I__10798 (
            .O(N__46828),
            .I(N__46822));
    InMux I__10797 (
            .O(N__46825),
            .I(N__46817));
    Span4Mux_h I__10796 (
            .O(N__46822),
            .I(N__46814));
    InMux I__10795 (
            .O(N__46821),
            .I(N__46809));
    InMux I__10794 (
            .O(N__46820),
            .I(N__46809));
    LocalMux I__10793 (
            .O(N__46817),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__10792 (
            .O(N__46814),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    LocalMux I__10791 (
            .O(N__46809),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    CascadeMux I__10790 (
            .O(N__46802),
            .I(N__46799));
    InMux I__10789 (
            .O(N__46799),
            .I(N__46796));
    LocalMux I__10788 (
            .O(N__46796),
            .I(N__46793));
    Span4Mux_v I__10787 (
            .O(N__46793),
            .I(N__46790));
    Span4Mux_h I__10786 (
            .O(N__46790),
            .I(N__46787));
    Span4Mux_s3_h I__10785 (
            .O(N__46787),
            .I(N__46784));
    Odrv4 I__10784 (
            .O(N__46784),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    CascadeMux I__10783 (
            .O(N__46781),
            .I(N__46778));
    InMux I__10782 (
            .O(N__46778),
            .I(N__46773));
    InMux I__10781 (
            .O(N__46777),
            .I(N__46770));
    InMux I__10780 (
            .O(N__46776),
            .I(N__46767));
    LocalMux I__10779 (
            .O(N__46773),
            .I(N__46762));
    LocalMux I__10778 (
            .O(N__46770),
            .I(N__46762));
    LocalMux I__10777 (
            .O(N__46767),
            .I(N__46757));
    Span4Mux_v I__10776 (
            .O(N__46762),
            .I(N__46757));
    Odrv4 I__10775 (
            .O(N__46757),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__10774 (
            .O(N__46754),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    CascadeMux I__10773 (
            .O(N__46751),
            .I(N__46748));
    InMux I__10772 (
            .O(N__46748),
            .I(N__46744));
    InMux I__10771 (
            .O(N__46747),
            .I(N__46741));
    LocalMux I__10770 (
            .O(N__46744),
            .I(N__46735));
    LocalMux I__10769 (
            .O(N__46741),
            .I(N__46735));
    InMux I__10768 (
            .O(N__46740),
            .I(N__46732));
    Span4Mux_v I__10767 (
            .O(N__46735),
            .I(N__46729));
    LocalMux I__10766 (
            .O(N__46732),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__10765 (
            .O(N__46729),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__10764 (
            .O(N__46724),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__10763 (
            .O(N__46721),
            .I(N__46718));
    LocalMux I__10762 (
            .O(N__46718),
            .I(N__46714));
    InMux I__10761 (
            .O(N__46717),
            .I(N__46711));
    Span4Mux_h I__10760 (
            .O(N__46714),
            .I(N__46708));
    LocalMux I__10759 (
            .O(N__46711),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__10758 (
            .O(N__46708),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__10757 (
            .O(N__46703),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__10756 (
            .O(N__46700),
            .I(N__46684));
    InMux I__10755 (
            .O(N__46699),
            .I(N__46684));
    InMux I__10754 (
            .O(N__46698),
            .I(N__46684));
    InMux I__10753 (
            .O(N__46697),
            .I(N__46684));
    InMux I__10752 (
            .O(N__46696),
            .I(N__46675));
    InMux I__10751 (
            .O(N__46695),
            .I(N__46675));
    InMux I__10750 (
            .O(N__46694),
            .I(N__46675));
    InMux I__10749 (
            .O(N__46693),
            .I(N__46675));
    LocalMux I__10748 (
            .O(N__46684),
            .I(N__46648));
    LocalMux I__10747 (
            .O(N__46675),
            .I(N__46648));
    InMux I__10746 (
            .O(N__46674),
            .I(N__46639));
    InMux I__10745 (
            .O(N__46673),
            .I(N__46639));
    InMux I__10744 (
            .O(N__46672),
            .I(N__46639));
    InMux I__10743 (
            .O(N__46671),
            .I(N__46639));
    InMux I__10742 (
            .O(N__46670),
            .I(N__46634));
    InMux I__10741 (
            .O(N__46669),
            .I(N__46634));
    InMux I__10740 (
            .O(N__46668),
            .I(N__46625));
    InMux I__10739 (
            .O(N__46667),
            .I(N__46625));
    InMux I__10738 (
            .O(N__46666),
            .I(N__46625));
    InMux I__10737 (
            .O(N__46665),
            .I(N__46625));
    InMux I__10736 (
            .O(N__46664),
            .I(N__46616));
    InMux I__10735 (
            .O(N__46663),
            .I(N__46616));
    InMux I__10734 (
            .O(N__46662),
            .I(N__46616));
    InMux I__10733 (
            .O(N__46661),
            .I(N__46616));
    InMux I__10732 (
            .O(N__46660),
            .I(N__46607));
    InMux I__10731 (
            .O(N__46659),
            .I(N__46607));
    InMux I__10730 (
            .O(N__46658),
            .I(N__46607));
    InMux I__10729 (
            .O(N__46657),
            .I(N__46607));
    InMux I__10728 (
            .O(N__46656),
            .I(N__46598));
    InMux I__10727 (
            .O(N__46655),
            .I(N__46598));
    InMux I__10726 (
            .O(N__46654),
            .I(N__46598));
    InMux I__10725 (
            .O(N__46653),
            .I(N__46598));
    Span4Mux_h I__10724 (
            .O(N__46648),
            .I(N__46591));
    LocalMux I__10723 (
            .O(N__46639),
            .I(N__46591));
    LocalMux I__10722 (
            .O(N__46634),
            .I(N__46591));
    LocalMux I__10721 (
            .O(N__46625),
            .I(N__46582));
    LocalMux I__10720 (
            .O(N__46616),
            .I(N__46582));
    LocalMux I__10719 (
            .O(N__46607),
            .I(N__46582));
    LocalMux I__10718 (
            .O(N__46598),
            .I(N__46582));
    Span4Mux_v I__10717 (
            .O(N__46591),
            .I(N__46577));
    Span4Mux_v I__10716 (
            .O(N__46582),
            .I(N__46577));
    Odrv4 I__10715 (
            .O(N__46577),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__10714 (
            .O(N__46574),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__10713 (
            .O(N__46571),
            .I(N__46568));
    LocalMux I__10712 (
            .O(N__46568),
            .I(N__46564));
    InMux I__10711 (
            .O(N__46567),
            .I(N__46561));
    Span4Mux_h I__10710 (
            .O(N__46564),
            .I(N__46558));
    LocalMux I__10709 (
            .O(N__46561),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__10708 (
            .O(N__46558),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__10707 (
            .O(N__46553),
            .I(N__46548));
    CEMux I__10706 (
            .O(N__46552),
            .I(N__46545));
    CEMux I__10705 (
            .O(N__46551),
            .I(N__46541));
    LocalMux I__10704 (
            .O(N__46548),
            .I(N__46538));
    LocalMux I__10703 (
            .O(N__46545),
            .I(N__46535));
    CEMux I__10702 (
            .O(N__46544),
            .I(N__46532));
    LocalMux I__10701 (
            .O(N__46541),
            .I(N__46529));
    Span4Mux_v I__10700 (
            .O(N__46538),
            .I(N__46526));
    Span4Mux_v I__10699 (
            .O(N__46535),
            .I(N__46523));
    LocalMux I__10698 (
            .O(N__46532),
            .I(N__46520));
    Span4Mux_h I__10697 (
            .O(N__46529),
            .I(N__46517));
    Span4Mux_h I__10696 (
            .O(N__46526),
            .I(N__46514));
    Span4Mux_h I__10695 (
            .O(N__46523),
            .I(N__46509));
    Span4Mux_h I__10694 (
            .O(N__46520),
            .I(N__46509));
    Odrv4 I__10693 (
            .O(N__46517),
            .I(\current_shift_inst.timer_s1.N_163_i ));
    Odrv4 I__10692 (
            .O(N__46514),
            .I(\current_shift_inst.timer_s1.N_163_i ));
    Odrv4 I__10691 (
            .O(N__46509),
            .I(\current_shift_inst.timer_s1.N_163_i ));
    IoInMux I__10690 (
            .O(N__46502),
            .I(N__46499));
    LocalMux I__10689 (
            .O(N__46499),
            .I(N__46495));
    InMux I__10688 (
            .O(N__46498),
            .I(N__46492));
    Odrv12 I__10687 (
            .O(N__46495),
            .I(T12_c));
    LocalMux I__10686 (
            .O(N__46492),
            .I(T12_c));
    InMux I__10685 (
            .O(N__46487),
            .I(N__46484));
    LocalMux I__10684 (
            .O(N__46484),
            .I(N__46480));
    InMux I__10683 (
            .O(N__46483),
            .I(N__46477));
    Span4Mux_v I__10682 (
            .O(N__46480),
            .I(N__46471));
    LocalMux I__10681 (
            .O(N__46477),
            .I(N__46471));
    InMux I__10680 (
            .O(N__46476),
            .I(N__46468));
    Span4Mux_h I__10679 (
            .O(N__46471),
            .I(N__46465));
    LocalMux I__10678 (
            .O(N__46468),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__10677 (
            .O(N__46465),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    InMux I__10676 (
            .O(N__46460),
            .I(N__46455));
    InMux I__10675 (
            .O(N__46459),
            .I(N__46452));
    InMux I__10674 (
            .O(N__46458),
            .I(N__46449));
    LocalMux I__10673 (
            .O(N__46455),
            .I(N__46445));
    LocalMux I__10672 (
            .O(N__46452),
            .I(N__46442));
    LocalMux I__10671 (
            .O(N__46449),
            .I(N__46439));
    InMux I__10670 (
            .O(N__46448),
            .I(N__46436));
    Span4Mux_v I__10669 (
            .O(N__46445),
            .I(N__46431));
    Span4Mux_v I__10668 (
            .O(N__46442),
            .I(N__46431));
    Span4Mux_v I__10667 (
            .O(N__46439),
            .I(N__46428));
    LocalMux I__10666 (
            .O(N__46436),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    Odrv4 I__10665 (
            .O(N__46431),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    Odrv4 I__10664 (
            .O(N__46428),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__10663 (
            .O(N__46421),
            .I(N__46418));
    LocalMux I__10662 (
            .O(N__46418),
            .I(N__46415));
    Span4Mux_h I__10661 (
            .O(N__46415),
            .I(N__46410));
    InMux I__10660 (
            .O(N__46414),
            .I(N__46406));
    InMux I__10659 (
            .O(N__46413),
            .I(N__46403));
    Span4Mux_v I__10658 (
            .O(N__46410),
            .I(N__46400));
    InMux I__10657 (
            .O(N__46409),
            .I(N__46397));
    LocalMux I__10656 (
            .O(N__46406),
            .I(N__46394));
    LocalMux I__10655 (
            .O(N__46403),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    Odrv4 I__10654 (
            .O(N__46400),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__10653 (
            .O(N__46397),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    Odrv4 I__10652 (
            .O(N__46394),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    CascadeMux I__10651 (
            .O(N__46385),
            .I(N__46380));
    InMux I__10650 (
            .O(N__46384),
            .I(N__46376));
    InMux I__10649 (
            .O(N__46383),
            .I(N__46373));
    InMux I__10648 (
            .O(N__46380),
            .I(N__46370));
    InMux I__10647 (
            .O(N__46379),
            .I(N__46367));
    LocalMux I__10646 (
            .O(N__46376),
            .I(N__46364));
    LocalMux I__10645 (
            .O(N__46373),
            .I(N__46361));
    LocalMux I__10644 (
            .O(N__46370),
            .I(N__46358));
    LocalMux I__10643 (
            .O(N__46367),
            .I(N__46355));
    Span4Mux_v I__10642 (
            .O(N__46364),
            .I(N__46350));
    Span4Mux_v I__10641 (
            .O(N__46361),
            .I(N__46350));
    Span4Mux_v I__10640 (
            .O(N__46358),
            .I(N__46347));
    Odrv4 I__10639 (
            .O(N__46355),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv4 I__10638 (
            .O(N__46350),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv4 I__10637 (
            .O(N__46347),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__10636 (
            .O(N__46340),
            .I(N__46336));
    InMux I__10635 (
            .O(N__46339),
            .I(N__46332));
    LocalMux I__10634 (
            .O(N__46336),
            .I(N__46328));
    InMux I__10633 (
            .O(N__46335),
            .I(N__46325));
    LocalMux I__10632 (
            .O(N__46332),
            .I(N__46322));
    InMux I__10631 (
            .O(N__46331),
            .I(N__46319));
    Span4Mux_h I__10630 (
            .O(N__46328),
            .I(N__46316));
    LocalMux I__10629 (
            .O(N__46325),
            .I(N__46309));
    Span4Mux_v I__10628 (
            .O(N__46322),
            .I(N__46309));
    LocalMux I__10627 (
            .O(N__46319),
            .I(N__46309));
    Odrv4 I__10626 (
            .O(N__46316),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    Odrv4 I__10625 (
            .O(N__46309),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    InMux I__10624 (
            .O(N__46304),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    CascadeMux I__10623 (
            .O(N__46301),
            .I(N__46298));
    InMux I__10622 (
            .O(N__46298),
            .I(N__46293));
    InMux I__10621 (
            .O(N__46297),
            .I(N__46290));
    InMux I__10620 (
            .O(N__46296),
            .I(N__46287));
    LocalMux I__10619 (
            .O(N__46293),
            .I(N__46282));
    LocalMux I__10618 (
            .O(N__46290),
            .I(N__46282));
    LocalMux I__10617 (
            .O(N__46287),
            .I(N__46277));
    Span4Mux_v I__10616 (
            .O(N__46282),
            .I(N__46277));
    Odrv4 I__10615 (
            .O(N__46277),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__10614 (
            .O(N__46274),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__10613 (
            .O(N__46271),
            .I(N__46265));
    InMux I__10612 (
            .O(N__46270),
            .I(N__46265));
    LocalMux I__10611 (
            .O(N__46265),
            .I(N__46261));
    InMux I__10610 (
            .O(N__46264),
            .I(N__46258));
    Span4Mux_v I__10609 (
            .O(N__46261),
            .I(N__46255));
    LocalMux I__10608 (
            .O(N__46258),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__10607 (
            .O(N__46255),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__10606 (
            .O(N__46250),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__10605 (
            .O(N__46247),
            .I(N__46244));
    InMux I__10604 (
            .O(N__46244),
            .I(N__46240));
    InMux I__10603 (
            .O(N__46243),
            .I(N__46237));
    LocalMux I__10602 (
            .O(N__46240),
            .I(N__46231));
    LocalMux I__10601 (
            .O(N__46237),
            .I(N__46231));
    InMux I__10600 (
            .O(N__46236),
            .I(N__46228));
    Span4Mux_h I__10599 (
            .O(N__46231),
            .I(N__46225));
    LocalMux I__10598 (
            .O(N__46228),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__10597 (
            .O(N__46225),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__10596 (
            .O(N__46220),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__10595 (
            .O(N__46217),
            .I(N__46213));
    CascadeMux I__10594 (
            .O(N__46216),
            .I(N__46210));
    InMux I__10593 (
            .O(N__46213),
            .I(N__46205));
    InMux I__10592 (
            .O(N__46210),
            .I(N__46205));
    LocalMux I__10591 (
            .O(N__46205),
            .I(N__46201));
    InMux I__10590 (
            .O(N__46204),
            .I(N__46198));
    Span4Mux_h I__10589 (
            .O(N__46201),
            .I(N__46195));
    LocalMux I__10588 (
            .O(N__46198),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__10587 (
            .O(N__46195),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__10586 (
            .O(N__46190),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__10585 (
            .O(N__46187),
            .I(N__46181));
    InMux I__10584 (
            .O(N__46186),
            .I(N__46181));
    LocalMux I__10583 (
            .O(N__46181),
            .I(N__46177));
    InMux I__10582 (
            .O(N__46180),
            .I(N__46174));
    Span4Mux_h I__10581 (
            .O(N__46177),
            .I(N__46171));
    LocalMux I__10580 (
            .O(N__46174),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__10579 (
            .O(N__46171),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__10578 (
            .O(N__46166),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__10577 (
            .O(N__46163),
            .I(N__46157));
    InMux I__10576 (
            .O(N__46162),
            .I(N__46157));
    LocalMux I__10575 (
            .O(N__46157),
            .I(N__46153));
    InMux I__10574 (
            .O(N__46156),
            .I(N__46150));
    Span4Mux_h I__10573 (
            .O(N__46153),
            .I(N__46147));
    LocalMux I__10572 (
            .O(N__46150),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__10571 (
            .O(N__46147),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__10570 (
            .O(N__46142),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    CascadeMux I__10569 (
            .O(N__46139),
            .I(N__46135));
    CascadeMux I__10568 (
            .O(N__46138),
            .I(N__46132));
    InMux I__10567 (
            .O(N__46135),
            .I(N__46129));
    InMux I__10566 (
            .O(N__46132),
            .I(N__46126));
    LocalMux I__10565 (
            .O(N__46129),
            .I(N__46122));
    LocalMux I__10564 (
            .O(N__46126),
            .I(N__46119));
    InMux I__10563 (
            .O(N__46125),
            .I(N__46116));
    Span4Mux_h I__10562 (
            .O(N__46122),
            .I(N__46113));
    Span4Mux_h I__10561 (
            .O(N__46119),
            .I(N__46110));
    LocalMux I__10560 (
            .O(N__46116),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__10559 (
            .O(N__46113),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__10558 (
            .O(N__46110),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__10557 (
            .O(N__46103),
            .I(bfn_18_20_0_));
    CascadeMux I__10556 (
            .O(N__46100),
            .I(N__46096));
    CascadeMux I__10555 (
            .O(N__46099),
            .I(N__46093));
    InMux I__10554 (
            .O(N__46096),
            .I(N__46090));
    InMux I__10553 (
            .O(N__46093),
            .I(N__46087));
    LocalMux I__10552 (
            .O(N__46090),
            .I(N__46083));
    LocalMux I__10551 (
            .O(N__46087),
            .I(N__46080));
    InMux I__10550 (
            .O(N__46086),
            .I(N__46077));
    Span4Mux_h I__10549 (
            .O(N__46083),
            .I(N__46074));
    Span4Mux_h I__10548 (
            .O(N__46080),
            .I(N__46071));
    LocalMux I__10547 (
            .O(N__46077),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__10546 (
            .O(N__46074),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__10545 (
            .O(N__46071),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__10544 (
            .O(N__46064),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__10543 (
            .O(N__46061),
            .I(N__46058));
    InMux I__10542 (
            .O(N__46058),
            .I(N__46054));
    InMux I__10541 (
            .O(N__46057),
            .I(N__46051));
    LocalMux I__10540 (
            .O(N__46054),
            .I(N__46047));
    LocalMux I__10539 (
            .O(N__46051),
            .I(N__46044));
    InMux I__10538 (
            .O(N__46050),
            .I(N__46041));
    Span4Mux_h I__10537 (
            .O(N__46047),
            .I(N__46038));
    Span4Mux_h I__10536 (
            .O(N__46044),
            .I(N__46035));
    LocalMux I__10535 (
            .O(N__46041),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__10534 (
            .O(N__46038),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__10533 (
            .O(N__46035),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__10532 (
            .O(N__46028),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__10531 (
            .O(N__46025),
            .I(N__46018));
    InMux I__10530 (
            .O(N__46024),
            .I(N__46018));
    InMux I__10529 (
            .O(N__46023),
            .I(N__46015));
    LocalMux I__10528 (
            .O(N__46018),
            .I(N__46012));
    LocalMux I__10527 (
            .O(N__46015),
            .I(N__46007));
    Span4Mux_v I__10526 (
            .O(N__46012),
            .I(N__46007));
    Odrv4 I__10525 (
            .O(N__46007),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__10524 (
            .O(N__46004),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__10523 (
            .O(N__46001),
            .I(N__45995));
    InMux I__10522 (
            .O(N__46000),
            .I(N__45995));
    LocalMux I__10521 (
            .O(N__45995),
            .I(N__45991));
    InMux I__10520 (
            .O(N__45994),
            .I(N__45988));
    Span4Mux_v I__10519 (
            .O(N__45991),
            .I(N__45985));
    LocalMux I__10518 (
            .O(N__45988),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__10517 (
            .O(N__45985),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__10516 (
            .O(N__45980),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    CascadeMux I__10515 (
            .O(N__45977),
            .I(N__45973));
    CascadeMux I__10514 (
            .O(N__45976),
            .I(N__45970));
    InMux I__10513 (
            .O(N__45973),
            .I(N__45965));
    InMux I__10512 (
            .O(N__45970),
            .I(N__45965));
    LocalMux I__10511 (
            .O(N__45965),
            .I(N__45961));
    InMux I__10510 (
            .O(N__45964),
            .I(N__45958));
    Span4Mux_h I__10509 (
            .O(N__45961),
            .I(N__45955));
    LocalMux I__10508 (
            .O(N__45958),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__10507 (
            .O(N__45955),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__10506 (
            .O(N__45950),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__10505 (
            .O(N__45947),
            .I(N__45943));
    CascadeMux I__10504 (
            .O(N__45946),
            .I(N__45940));
    InMux I__10503 (
            .O(N__45943),
            .I(N__45935));
    InMux I__10502 (
            .O(N__45940),
            .I(N__45935));
    LocalMux I__10501 (
            .O(N__45935),
            .I(N__45931));
    InMux I__10500 (
            .O(N__45934),
            .I(N__45928));
    Span4Mux_h I__10499 (
            .O(N__45931),
            .I(N__45925));
    LocalMux I__10498 (
            .O(N__45928),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__10497 (
            .O(N__45925),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__10496 (
            .O(N__45920),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__10495 (
            .O(N__45917),
            .I(N__45911));
    InMux I__10494 (
            .O(N__45916),
            .I(N__45911));
    LocalMux I__10493 (
            .O(N__45911),
            .I(N__45907));
    InMux I__10492 (
            .O(N__45910),
            .I(N__45904));
    Span4Mux_h I__10491 (
            .O(N__45907),
            .I(N__45901));
    LocalMux I__10490 (
            .O(N__45904),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__10489 (
            .O(N__45901),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__10488 (
            .O(N__45896),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    CascadeMux I__10487 (
            .O(N__45893),
            .I(N__45890));
    InMux I__10486 (
            .O(N__45890),
            .I(N__45886));
    InMux I__10485 (
            .O(N__45889),
            .I(N__45883));
    LocalMux I__10484 (
            .O(N__45886),
            .I(N__45877));
    LocalMux I__10483 (
            .O(N__45883),
            .I(N__45877));
    InMux I__10482 (
            .O(N__45882),
            .I(N__45874));
    Span4Mux_h I__10481 (
            .O(N__45877),
            .I(N__45871));
    LocalMux I__10480 (
            .O(N__45874),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__10479 (
            .O(N__45871),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__10478 (
            .O(N__45866),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__10477 (
            .O(N__45863),
            .I(N__45859));
    CascadeMux I__10476 (
            .O(N__45862),
            .I(N__45856));
    InMux I__10475 (
            .O(N__45859),
            .I(N__45853));
    InMux I__10474 (
            .O(N__45856),
            .I(N__45850));
    LocalMux I__10473 (
            .O(N__45853),
            .I(N__45846));
    LocalMux I__10472 (
            .O(N__45850),
            .I(N__45843));
    InMux I__10471 (
            .O(N__45849),
            .I(N__45840));
    Span4Mux_h I__10470 (
            .O(N__45846),
            .I(N__45837));
    Span4Mux_h I__10469 (
            .O(N__45843),
            .I(N__45834));
    LocalMux I__10468 (
            .O(N__45840),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__10467 (
            .O(N__45837),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__10466 (
            .O(N__45834),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__10465 (
            .O(N__45827),
            .I(bfn_18_19_0_));
    CascadeMux I__10464 (
            .O(N__45824),
            .I(N__45821));
    InMux I__10463 (
            .O(N__45821),
            .I(N__45817));
    InMux I__10462 (
            .O(N__45820),
            .I(N__45814));
    LocalMux I__10461 (
            .O(N__45817),
            .I(N__45810));
    LocalMux I__10460 (
            .O(N__45814),
            .I(N__45807));
    InMux I__10459 (
            .O(N__45813),
            .I(N__45804));
    Span4Mux_h I__10458 (
            .O(N__45810),
            .I(N__45801));
    Span4Mux_h I__10457 (
            .O(N__45807),
            .I(N__45798));
    LocalMux I__10456 (
            .O(N__45804),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__10455 (
            .O(N__45801),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__10454 (
            .O(N__45798),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__10453 (
            .O(N__45791),
            .I(N__45787));
    InMux I__10452 (
            .O(N__45790),
            .I(N__45784));
    LocalMux I__10451 (
            .O(N__45787),
            .I(N__45780));
    LocalMux I__10450 (
            .O(N__45784),
            .I(N__45777));
    InMux I__10449 (
            .O(N__45783),
            .I(N__45774));
    Span4Mux_h I__10448 (
            .O(N__45780),
            .I(N__45771));
    Odrv4 I__10447 (
            .O(N__45777),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__10446 (
            .O(N__45774),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__10445 (
            .O(N__45771),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__10444 (
            .O(N__45764),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    CascadeMux I__10443 (
            .O(N__45761),
            .I(N__45757));
    CascadeMux I__10442 (
            .O(N__45760),
            .I(N__45754));
    InMux I__10441 (
            .O(N__45757),
            .I(N__45748));
    InMux I__10440 (
            .O(N__45754),
            .I(N__45748));
    InMux I__10439 (
            .O(N__45753),
            .I(N__45745));
    LocalMux I__10438 (
            .O(N__45748),
            .I(N__45742));
    LocalMux I__10437 (
            .O(N__45745),
            .I(N__45737));
    Span4Mux_v I__10436 (
            .O(N__45742),
            .I(N__45737));
    Odrv4 I__10435 (
            .O(N__45737),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__10434 (
            .O(N__45734),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    CascadeMux I__10433 (
            .O(N__45731),
            .I(N__45727));
    CascadeMux I__10432 (
            .O(N__45730),
            .I(N__45724));
    InMux I__10431 (
            .O(N__45727),
            .I(N__45719));
    InMux I__10430 (
            .O(N__45724),
            .I(N__45719));
    LocalMux I__10429 (
            .O(N__45719),
            .I(N__45715));
    InMux I__10428 (
            .O(N__45718),
            .I(N__45712));
    Span4Mux_v I__10427 (
            .O(N__45715),
            .I(N__45709));
    LocalMux I__10426 (
            .O(N__45712),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__10425 (
            .O(N__45709),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__10424 (
            .O(N__45704),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__10423 (
            .O(N__45701),
            .I(N__45698));
    InMux I__10422 (
            .O(N__45698),
            .I(N__45694));
    InMux I__10421 (
            .O(N__45697),
            .I(N__45691));
    LocalMux I__10420 (
            .O(N__45694),
            .I(N__45685));
    LocalMux I__10419 (
            .O(N__45691),
            .I(N__45685));
    InMux I__10418 (
            .O(N__45690),
            .I(N__45682));
    Span4Mux_h I__10417 (
            .O(N__45685),
            .I(N__45679));
    LocalMux I__10416 (
            .O(N__45682),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__10415 (
            .O(N__45679),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__10414 (
            .O(N__45674),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__10413 (
            .O(N__45671),
            .I(N__45668));
    InMux I__10412 (
            .O(N__45668),
            .I(N__45664));
    InMux I__10411 (
            .O(N__45667),
            .I(N__45661));
    LocalMux I__10410 (
            .O(N__45664),
            .I(N__45655));
    LocalMux I__10409 (
            .O(N__45661),
            .I(N__45655));
    InMux I__10408 (
            .O(N__45660),
            .I(N__45652));
    Span4Mux_h I__10407 (
            .O(N__45655),
            .I(N__45649));
    LocalMux I__10406 (
            .O(N__45652),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__10405 (
            .O(N__45649),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__10404 (
            .O(N__45644),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    CascadeMux I__10403 (
            .O(N__45641),
            .I(N__45638));
    InMux I__10402 (
            .O(N__45638),
            .I(N__45634));
    InMux I__10401 (
            .O(N__45637),
            .I(N__45631));
    LocalMux I__10400 (
            .O(N__45634),
            .I(N__45625));
    LocalMux I__10399 (
            .O(N__45631),
            .I(N__45625));
    InMux I__10398 (
            .O(N__45630),
            .I(N__45622));
    Span4Mux_h I__10397 (
            .O(N__45625),
            .I(N__45619));
    LocalMux I__10396 (
            .O(N__45622),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__10395 (
            .O(N__45619),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__10394 (
            .O(N__45614),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    CascadeMux I__10393 (
            .O(N__45611),
            .I(N__45608));
    InMux I__10392 (
            .O(N__45608),
            .I(N__45604));
    InMux I__10391 (
            .O(N__45607),
            .I(N__45601));
    LocalMux I__10390 (
            .O(N__45604),
            .I(N__45595));
    LocalMux I__10389 (
            .O(N__45601),
            .I(N__45595));
    InMux I__10388 (
            .O(N__45600),
            .I(N__45592));
    Span4Mux_h I__10387 (
            .O(N__45595),
            .I(N__45589));
    LocalMux I__10386 (
            .O(N__45592),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__10385 (
            .O(N__45589),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__10384 (
            .O(N__45584),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__10383 (
            .O(N__45581),
            .I(N__45578));
    InMux I__10382 (
            .O(N__45578),
            .I(N__45574));
    InMux I__10381 (
            .O(N__45577),
            .I(N__45571));
    LocalMux I__10380 (
            .O(N__45574),
            .I(N__45567));
    LocalMux I__10379 (
            .O(N__45571),
            .I(N__45564));
    InMux I__10378 (
            .O(N__45570),
            .I(N__45561));
    Span4Mux_h I__10377 (
            .O(N__45567),
            .I(N__45558));
    Span4Mux_h I__10376 (
            .O(N__45564),
            .I(N__45555));
    LocalMux I__10375 (
            .O(N__45561),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__10374 (
            .O(N__45558),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__10373 (
            .O(N__45555),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__10372 (
            .O(N__45548),
            .I(bfn_18_18_0_));
    InMux I__10371 (
            .O(N__45545),
            .I(N__45539));
    InMux I__10370 (
            .O(N__45544),
            .I(N__45539));
    LocalMux I__10369 (
            .O(N__45539),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ));
    CascadeMux I__10368 (
            .O(N__45536),
            .I(N__45533));
    InMux I__10367 (
            .O(N__45533),
            .I(N__45527));
    InMux I__10366 (
            .O(N__45532),
            .I(N__45527));
    LocalMux I__10365 (
            .O(N__45527),
            .I(N__45523));
    InMux I__10364 (
            .O(N__45526),
            .I(N__45520));
    Span4Mux_h I__10363 (
            .O(N__45523),
            .I(N__45517));
    LocalMux I__10362 (
            .O(N__45520),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv4 I__10361 (
            .O(N__45517),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__10360 (
            .O(N__45512),
            .I(N__45506));
    InMux I__10359 (
            .O(N__45511),
            .I(N__45506));
    LocalMux I__10358 (
            .O(N__45506),
            .I(N__45502));
    InMux I__10357 (
            .O(N__45505),
            .I(N__45499));
    Span12Mux_v I__10356 (
            .O(N__45502),
            .I(N__45496));
    LocalMux I__10355 (
            .O(N__45499),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv12 I__10354 (
            .O(N__45496),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__10353 (
            .O(N__45491),
            .I(N__45488));
    LocalMux I__10352 (
            .O(N__45488),
            .I(N__45485));
    Odrv4 I__10351 (
            .O(N__45485),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt28 ));
    CascadeMux I__10350 (
            .O(N__45482),
            .I(N__45477));
    InMux I__10349 (
            .O(N__45481),
            .I(N__45474));
    InMux I__10348 (
            .O(N__45480),
            .I(N__45471));
    InMux I__10347 (
            .O(N__45477),
            .I(N__45468));
    LocalMux I__10346 (
            .O(N__45474),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__10345 (
            .O(N__45471),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__10344 (
            .O(N__45468),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__10343 (
            .O(N__45461),
            .I(N__45458));
    LocalMux I__10342 (
            .O(N__45458),
            .I(\current_shift_inst.un4_control_input1_1 ));
    InMux I__10341 (
            .O(N__45455),
            .I(N__45426));
    InMux I__10340 (
            .O(N__45454),
            .I(N__45426));
    InMux I__10339 (
            .O(N__45453),
            .I(N__45419));
    InMux I__10338 (
            .O(N__45452),
            .I(N__45419));
    CascadeMux I__10337 (
            .O(N__45451),
            .I(N__45411));
    InMux I__10336 (
            .O(N__45450),
            .I(N__45401));
    CascadeMux I__10335 (
            .O(N__45449),
            .I(N__45393));
    CascadeMux I__10334 (
            .O(N__45448),
            .I(N__45387));
    CascadeMux I__10333 (
            .O(N__45447),
            .I(N__45379));
    InMux I__10332 (
            .O(N__45446),
            .I(N__45369));
    InMux I__10331 (
            .O(N__45445),
            .I(N__45369));
    InMux I__10330 (
            .O(N__45444),
            .I(N__45369));
    InMux I__10329 (
            .O(N__45443),
            .I(N__45362));
    InMux I__10328 (
            .O(N__45442),
            .I(N__45362));
    InMux I__10327 (
            .O(N__45441),
            .I(N__45362));
    InMux I__10326 (
            .O(N__45440),
            .I(N__45359));
    InMux I__10325 (
            .O(N__45439),
            .I(N__45352));
    InMux I__10324 (
            .O(N__45438),
            .I(N__45352));
    InMux I__10323 (
            .O(N__45437),
            .I(N__45352));
    InMux I__10322 (
            .O(N__45436),
            .I(N__45339));
    InMux I__10321 (
            .O(N__45435),
            .I(N__45339));
    InMux I__10320 (
            .O(N__45434),
            .I(N__45339));
    InMux I__10319 (
            .O(N__45433),
            .I(N__45339));
    InMux I__10318 (
            .O(N__45432),
            .I(N__45339));
    InMux I__10317 (
            .O(N__45431),
            .I(N__45339));
    LocalMux I__10316 (
            .O(N__45426),
            .I(N__45336));
    InMux I__10315 (
            .O(N__45425),
            .I(N__45330));
    InMux I__10314 (
            .O(N__45424),
            .I(N__45330));
    LocalMux I__10313 (
            .O(N__45419),
            .I(N__45327));
    InMux I__10312 (
            .O(N__45418),
            .I(N__45324));
    InMux I__10311 (
            .O(N__45417),
            .I(N__45319));
    InMux I__10310 (
            .O(N__45416),
            .I(N__45319));
    InMux I__10309 (
            .O(N__45415),
            .I(N__45304));
    InMux I__10308 (
            .O(N__45414),
            .I(N__45304));
    InMux I__10307 (
            .O(N__45411),
            .I(N__45304));
    InMux I__10306 (
            .O(N__45410),
            .I(N__45304));
    InMux I__10305 (
            .O(N__45409),
            .I(N__45304));
    InMux I__10304 (
            .O(N__45408),
            .I(N__45304));
    InMux I__10303 (
            .O(N__45407),
            .I(N__45304));
    InMux I__10302 (
            .O(N__45406),
            .I(N__45297));
    InMux I__10301 (
            .O(N__45405),
            .I(N__45297));
    InMux I__10300 (
            .O(N__45404),
            .I(N__45297));
    LocalMux I__10299 (
            .O(N__45401),
            .I(N__45294));
    InMux I__10298 (
            .O(N__45400),
            .I(N__45285));
    InMux I__10297 (
            .O(N__45399),
            .I(N__45285));
    InMux I__10296 (
            .O(N__45398),
            .I(N__45285));
    InMux I__10295 (
            .O(N__45397),
            .I(N__45285));
    InMux I__10294 (
            .O(N__45396),
            .I(N__45262));
    InMux I__10293 (
            .O(N__45393),
            .I(N__45262));
    InMux I__10292 (
            .O(N__45392),
            .I(N__45262));
    InMux I__10291 (
            .O(N__45391),
            .I(N__45262));
    InMux I__10290 (
            .O(N__45390),
            .I(N__45262));
    InMux I__10289 (
            .O(N__45387),
            .I(N__45262));
    InMux I__10288 (
            .O(N__45386),
            .I(N__45262));
    InMux I__10287 (
            .O(N__45385),
            .I(N__45247));
    InMux I__10286 (
            .O(N__45384),
            .I(N__45247));
    InMux I__10285 (
            .O(N__45383),
            .I(N__45247));
    InMux I__10284 (
            .O(N__45382),
            .I(N__45247));
    InMux I__10283 (
            .O(N__45379),
            .I(N__45247));
    InMux I__10282 (
            .O(N__45378),
            .I(N__45247));
    InMux I__10281 (
            .O(N__45377),
            .I(N__45247));
    InMux I__10280 (
            .O(N__45376),
            .I(N__45244));
    LocalMux I__10279 (
            .O(N__45369),
            .I(N__45241));
    LocalMux I__10278 (
            .O(N__45362),
            .I(N__45236));
    LocalMux I__10277 (
            .O(N__45359),
            .I(N__45236));
    LocalMux I__10276 (
            .O(N__45352),
            .I(N__45233));
    LocalMux I__10275 (
            .O(N__45339),
            .I(N__45228));
    Span4Mux_h I__10274 (
            .O(N__45336),
            .I(N__45228));
    InMux I__10273 (
            .O(N__45335),
            .I(N__45225));
    LocalMux I__10272 (
            .O(N__45330),
            .I(N__45209));
    Span4Mux_v I__10271 (
            .O(N__45327),
            .I(N__45209));
    LocalMux I__10270 (
            .O(N__45324),
            .I(N__45209));
    LocalMux I__10269 (
            .O(N__45319),
            .I(N__45209));
    LocalMux I__10268 (
            .O(N__45304),
            .I(N__45206));
    LocalMux I__10267 (
            .O(N__45297),
            .I(N__45203));
    Span4Mux_h I__10266 (
            .O(N__45294),
            .I(N__45198));
    LocalMux I__10265 (
            .O(N__45285),
            .I(N__45198));
    InMux I__10264 (
            .O(N__45284),
            .I(N__45195));
    InMux I__10263 (
            .O(N__45283),
            .I(N__45190));
    InMux I__10262 (
            .O(N__45282),
            .I(N__45190));
    InMux I__10261 (
            .O(N__45281),
            .I(N__45185));
    InMux I__10260 (
            .O(N__45280),
            .I(N__45185));
    InMux I__10259 (
            .O(N__45279),
            .I(N__45178));
    InMux I__10258 (
            .O(N__45278),
            .I(N__45178));
    InMux I__10257 (
            .O(N__45277),
            .I(N__45178));
    LocalMux I__10256 (
            .O(N__45262),
            .I(N__45173));
    LocalMux I__10255 (
            .O(N__45247),
            .I(N__45173));
    LocalMux I__10254 (
            .O(N__45244),
            .I(N__45170));
    Span4Mux_h I__10253 (
            .O(N__45241),
            .I(N__45165));
    Span4Mux_h I__10252 (
            .O(N__45236),
            .I(N__45165));
    Span4Mux_v I__10251 (
            .O(N__45233),
            .I(N__45158));
    Span4Mux_v I__10250 (
            .O(N__45228),
            .I(N__45158));
    LocalMux I__10249 (
            .O(N__45225),
            .I(N__45158));
    InMux I__10248 (
            .O(N__45224),
            .I(N__45151));
    InMux I__10247 (
            .O(N__45223),
            .I(N__45151));
    InMux I__10246 (
            .O(N__45222),
            .I(N__45151));
    InMux I__10245 (
            .O(N__45221),
            .I(N__45142));
    InMux I__10244 (
            .O(N__45220),
            .I(N__45142));
    InMux I__10243 (
            .O(N__45219),
            .I(N__45142));
    InMux I__10242 (
            .O(N__45218),
            .I(N__45142));
    Span4Mux_v I__10241 (
            .O(N__45209),
            .I(N__45139));
    Span4Mux_v I__10240 (
            .O(N__45206),
            .I(N__45132));
    Span4Mux_h I__10239 (
            .O(N__45203),
            .I(N__45132));
    Span4Mux_v I__10238 (
            .O(N__45198),
            .I(N__45132));
    LocalMux I__10237 (
            .O(N__45195),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10236 (
            .O(N__45190),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10235 (
            .O(N__45185),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10234 (
            .O(N__45178),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10233 (
            .O(N__45173),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10232 (
            .O(N__45170),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10231 (
            .O(N__45165),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10230 (
            .O(N__45158),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10229 (
            .O(N__45151),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10228 (
            .O(N__45142),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10227 (
            .O(N__45139),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10226 (
            .O(N__45132),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__10225 (
            .O(N__45107),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__10224 (
            .O(N__45104),
            .I(N__45098));
    InMux I__10223 (
            .O(N__45103),
            .I(N__45095));
    InMux I__10222 (
            .O(N__45102),
            .I(N__45090));
    InMux I__10221 (
            .O(N__45101),
            .I(N__45090));
    LocalMux I__10220 (
            .O(N__45098),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__10219 (
            .O(N__45095),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__10218 (
            .O(N__45090),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    InMux I__10217 (
            .O(N__45083),
            .I(N__45080));
    LocalMux I__10216 (
            .O(N__45080),
            .I(N__45077));
    Span4Mux_v I__10215 (
            .O(N__45077),
            .I(N__45073));
    InMux I__10214 (
            .O(N__45076),
            .I(N__45070));
    Span4Mux_h I__10213 (
            .O(N__45073),
            .I(N__45067));
    LocalMux I__10212 (
            .O(N__45070),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv4 I__10211 (
            .O(N__45067),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    CascadeMux I__10210 (
            .O(N__45062),
            .I(N__45059));
    InMux I__10209 (
            .O(N__45059),
            .I(N__45055));
    InMux I__10208 (
            .O(N__45058),
            .I(N__45052));
    LocalMux I__10207 (
            .O(N__45055),
            .I(N__45049));
    LocalMux I__10206 (
            .O(N__45052),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    Odrv12 I__10205 (
            .O(N__45049),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__10204 (
            .O(N__45044),
            .I(N__45038));
    InMux I__10203 (
            .O(N__45043),
            .I(N__45035));
    InMux I__10202 (
            .O(N__45042),
            .I(N__45028));
    InMux I__10201 (
            .O(N__45041),
            .I(N__45028));
    LocalMux I__10200 (
            .O(N__45038),
            .I(N__45023));
    LocalMux I__10199 (
            .O(N__45035),
            .I(N__45023));
    InMux I__10198 (
            .O(N__45034),
            .I(N__45020));
    InMux I__10197 (
            .O(N__45033),
            .I(N__45017));
    LocalMux I__10196 (
            .O(N__45028),
            .I(N__45014));
    Span4Mux_v I__10195 (
            .O(N__45023),
            .I(N__45011));
    LocalMux I__10194 (
            .O(N__45020),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__10193 (
            .O(N__45017),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv12 I__10192 (
            .O(N__45014),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__10191 (
            .O(N__45011),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    InMux I__10190 (
            .O(N__45002),
            .I(N__44998));
    InMux I__10189 (
            .O(N__45001),
            .I(N__44994));
    LocalMux I__10188 (
            .O(N__44998),
            .I(N__44991));
    InMux I__10187 (
            .O(N__44997),
            .I(N__44988));
    LocalMux I__10186 (
            .O(N__44994),
            .I(N__44985));
    Span4Mux_v I__10185 (
            .O(N__44991),
            .I(N__44982));
    LocalMux I__10184 (
            .O(N__44988),
            .I(N__44979));
    Span4Mux_v I__10183 (
            .O(N__44985),
            .I(N__44976));
    Span4Mux_v I__10182 (
            .O(N__44982),
            .I(N__44971));
    Span4Mux_v I__10181 (
            .O(N__44979),
            .I(N__44971));
    Odrv4 I__10180 (
            .O(N__44976),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__10179 (
            .O(N__44971),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__10178 (
            .O(N__44966),
            .I(N__44963));
    LocalMux I__10177 (
            .O(N__44963),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    CEMux I__10176 (
            .O(N__44960),
            .I(N__44936));
    CEMux I__10175 (
            .O(N__44959),
            .I(N__44936));
    CEMux I__10174 (
            .O(N__44958),
            .I(N__44936));
    CEMux I__10173 (
            .O(N__44957),
            .I(N__44936));
    CEMux I__10172 (
            .O(N__44956),
            .I(N__44936));
    CEMux I__10171 (
            .O(N__44955),
            .I(N__44936));
    CEMux I__10170 (
            .O(N__44954),
            .I(N__44936));
    CEMux I__10169 (
            .O(N__44953),
            .I(N__44936));
    GlobalMux I__10168 (
            .O(N__44936),
            .I(N__44933));
    gio2CtrlBuf I__10167 (
            .O(N__44933),
            .I(\current_shift_inst.timer_s1.N_162_i_g ));
    InMux I__10166 (
            .O(N__44930),
            .I(N__44923));
    InMux I__10165 (
            .O(N__44929),
            .I(N__44923));
    InMux I__10164 (
            .O(N__44928),
            .I(N__44920));
    LocalMux I__10163 (
            .O(N__44923),
            .I(N__44917));
    LocalMux I__10162 (
            .O(N__44920),
            .I(N__44893));
    Span4Mux_v I__10161 (
            .O(N__44917),
            .I(N__44893));
    InMux I__10160 (
            .O(N__44916),
            .I(N__44884));
    InMux I__10159 (
            .O(N__44915),
            .I(N__44884));
    InMux I__10158 (
            .O(N__44914),
            .I(N__44884));
    InMux I__10157 (
            .O(N__44913),
            .I(N__44884));
    InMux I__10156 (
            .O(N__44912),
            .I(N__44873));
    InMux I__10155 (
            .O(N__44911),
            .I(N__44873));
    InMux I__10154 (
            .O(N__44910),
            .I(N__44873));
    InMux I__10153 (
            .O(N__44909),
            .I(N__44873));
    InMux I__10152 (
            .O(N__44908),
            .I(N__44873));
    InMux I__10151 (
            .O(N__44907),
            .I(N__44866));
    InMux I__10150 (
            .O(N__44906),
            .I(N__44866));
    InMux I__10149 (
            .O(N__44905),
            .I(N__44866));
    InMux I__10148 (
            .O(N__44904),
            .I(N__44860));
    InMux I__10147 (
            .O(N__44903),
            .I(N__44849));
    InMux I__10146 (
            .O(N__44902),
            .I(N__44849));
    InMux I__10145 (
            .O(N__44901),
            .I(N__44849));
    InMux I__10144 (
            .O(N__44900),
            .I(N__44849));
    InMux I__10143 (
            .O(N__44899),
            .I(N__44849));
    InMux I__10142 (
            .O(N__44898),
            .I(N__44846));
    Sp12to4 I__10141 (
            .O(N__44893),
            .I(N__44837));
    LocalMux I__10140 (
            .O(N__44884),
            .I(N__44837));
    LocalMux I__10139 (
            .O(N__44873),
            .I(N__44837));
    LocalMux I__10138 (
            .O(N__44866),
            .I(N__44837));
    InMux I__10137 (
            .O(N__44865),
            .I(N__44834));
    InMux I__10136 (
            .O(N__44864),
            .I(N__44829));
    InMux I__10135 (
            .O(N__44863),
            .I(N__44829));
    LocalMux I__10134 (
            .O(N__44860),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10133 (
            .O(N__44849),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10132 (
            .O(N__44846),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv12 I__10131 (
            .O(N__44837),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10130 (
            .O(N__44834),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10129 (
            .O(N__44829),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__10128 (
            .O(N__44816),
            .I(N__44813));
    LocalMux I__10127 (
            .O(N__44813),
            .I(N__44808));
    InMux I__10126 (
            .O(N__44812),
            .I(N__44805));
    InMux I__10125 (
            .O(N__44811),
            .I(N__44802));
    Span4Mux_v I__10124 (
            .O(N__44808),
            .I(N__44799));
    LocalMux I__10123 (
            .O(N__44805),
            .I(N__44794));
    LocalMux I__10122 (
            .O(N__44802),
            .I(N__44794));
    Odrv4 I__10121 (
            .O(N__44799),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__10120 (
            .O(N__44794),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__10119 (
            .O(N__44789),
            .I(N__44786));
    LocalMux I__10118 (
            .O(N__44786),
            .I(N__44783));
    Span4Mux_v I__10117 (
            .O(N__44783),
            .I(N__44780));
    Odrv4 I__10116 (
            .O(N__44780),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__10115 (
            .O(N__44777),
            .I(N__44771));
    InMux I__10114 (
            .O(N__44776),
            .I(N__44768));
    InMux I__10113 (
            .O(N__44775),
            .I(N__44763));
    InMux I__10112 (
            .O(N__44774),
            .I(N__44763));
    LocalMux I__10111 (
            .O(N__44771),
            .I(N__44760));
    LocalMux I__10110 (
            .O(N__44768),
            .I(N__44757));
    LocalMux I__10109 (
            .O(N__44763),
            .I(N__44754));
    Span4Mux_h I__10108 (
            .O(N__44760),
            .I(N__44751));
    Span4Mux_v I__10107 (
            .O(N__44757),
            .I(N__44746));
    Span4Mux_h I__10106 (
            .O(N__44754),
            .I(N__44746));
    Odrv4 I__10105 (
            .O(N__44751),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__10104 (
            .O(N__44746),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__10103 (
            .O(N__44741),
            .I(N__44738));
    LocalMux I__10102 (
            .O(N__44738),
            .I(N__44735));
    Odrv4 I__10101 (
            .O(N__44735),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__10100 (
            .O(N__44732),
            .I(N__44728));
    InMux I__10099 (
            .O(N__44731),
            .I(N__44725));
    LocalMux I__10098 (
            .O(N__44728),
            .I(N__44721));
    LocalMux I__10097 (
            .O(N__44725),
            .I(N__44718));
    InMux I__10096 (
            .O(N__44724),
            .I(N__44715));
    Span4Mux_h I__10095 (
            .O(N__44721),
            .I(N__44712));
    Odrv4 I__10094 (
            .O(N__44718),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__10093 (
            .O(N__44715),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__10092 (
            .O(N__44712),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__10091 (
            .O(N__44705),
            .I(bfn_18_17_0_));
    InMux I__10090 (
            .O(N__44702),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__10089 (
            .O(N__44699),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__10088 (
            .O(N__44696),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    CascadeMux I__10087 (
            .O(N__44693),
            .I(N__44689));
    CascadeMux I__10086 (
            .O(N__44692),
            .I(N__44686));
    InMux I__10085 (
            .O(N__44689),
            .I(N__44681));
    InMux I__10084 (
            .O(N__44686),
            .I(N__44681));
    LocalMux I__10083 (
            .O(N__44681),
            .I(N__44677));
    InMux I__10082 (
            .O(N__44680),
            .I(N__44674));
    Span4Mux_v I__10081 (
            .O(N__44677),
            .I(N__44671));
    LocalMux I__10080 (
            .O(N__44674),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__10079 (
            .O(N__44671),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__10078 (
            .O(N__44666),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__10077 (
            .O(N__44663),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__10076 (
            .O(N__44660),
            .I(N__44654));
    InMux I__10075 (
            .O(N__44659),
            .I(N__44654));
    LocalMux I__10074 (
            .O(N__44654),
            .I(N__44650));
    InMux I__10073 (
            .O(N__44653),
            .I(N__44647));
    Span4Mux_v I__10072 (
            .O(N__44650),
            .I(N__44644));
    LocalMux I__10071 (
            .O(N__44647),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__10070 (
            .O(N__44644),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__10069 (
            .O(N__44639),
            .I(N__44636));
    InMux I__10068 (
            .O(N__44636),
            .I(N__44633));
    LocalMux I__10067 (
            .O(N__44633),
            .I(N__44630));
    Span4Mux_h I__10066 (
            .O(N__44630),
            .I(N__44627));
    Odrv4 I__10065 (
            .O(N__44627),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt26 ));
    CascadeMux I__10064 (
            .O(N__44624),
            .I(N__44620));
    InMux I__10063 (
            .O(N__44623),
            .I(N__44615));
    InMux I__10062 (
            .O(N__44620),
            .I(N__44615));
    LocalMux I__10061 (
            .O(N__44615),
            .I(N__44611));
    InMux I__10060 (
            .O(N__44614),
            .I(N__44608));
    Span4Mux_v I__10059 (
            .O(N__44611),
            .I(N__44605));
    LocalMux I__10058 (
            .O(N__44608),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    Odrv4 I__10057 (
            .O(N__44605),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    CascadeMux I__10056 (
            .O(N__44600),
            .I(N__44597));
    InMux I__10055 (
            .O(N__44597),
            .I(N__44593));
    InMux I__10054 (
            .O(N__44596),
            .I(N__44590));
    LocalMux I__10053 (
            .O(N__44593),
            .I(N__44584));
    LocalMux I__10052 (
            .O(N__44590),
            .I(N__44584));
    InMux I__10051 (
            .O(N__44589),
            .I(N__44581));
    Span4Mux_v I__10050 (
            .O(N__44584),
            .I(N__44578));
    LocalMux I__10049 (
            .O(N__44581),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    Odrv4 I__10048 (
            .O(N__44578),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__10047 (
            .O(N__44573),
            .I(N__44570));
    LocalMux I__10046 (
            .O(N__44570),
            .I(N__44567));
    Odrv12 I__10045 (
            .O(N__44567),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ));
    CascadeMux I__10044 (
            .O(N__44564),
            .I(N__44561));
    InMux I__10043 (
            .O(N__44561),
            .I(N__44558));
    LocalMux I__10042 (
            .O(N__44558),
            .I(N__44555));
    Odrv4 I__10041 (
            .O(N__44555),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ));
    CascadeMux I__10040 (
            .O(N__44552),
            .I(N__44549));
    InMux I__10039 (
            .O(N__44549),
            .I(N__44542));
    InMux I__10038 (
            .O(N__44548),
            .I(N__44542));
    InMux I__10037 (
            .O(N__44547),
            .I(N__44539));
    LocalMux I__10036 (
            .O(N__44542),
            .I(N__44536));
    LocalMux I__10035 (
            .O(N__44539),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv12 I__10034 (
            .O(N__44536),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__10033 (
            .O(N__44531),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__10032 (
            .O(N__44528),
            .I(N__44521));
    InMux I__10031 (
            .O(N__44527),
            .I(N__44521));
    InMux I__10030 (
            .O(N__44526),
            .I(N__44518));
    LocalMux I__10029 (
            .O(N__44521),
            .I(N__44515));
    LocalMux I__10028 (
            .O(N__44518),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv12 I__10027 (
            .O(N__44515),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__10026 (
            .O(N__44510),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    CascadeMux I__10025 (
            .O(N__44507),
            .I(N__44503));
    InMux I__10024 (
            .O(N__44506),
            .I(N__44497));
    InMux I__10023 (
            .O(N__44503),
            .I(N__44497));
    InMux I__10022 (
            .O(N__44502),
            .I(N__44494));
    LocalMux I__10021 (
            .O(N__44497),
            .I(N__44491));
    LocalMux I__10020 (
            .O(N__44494),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv12 I__10019 (
            .O(N__44491),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__10018 (
            .O(N__44486),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    CascadeMux I__10017 (
            .O(N__44483),
            .I(N__44480));
    InMux I__10016 (
            .O(N__44480),
            .I(N__44475));
    InMux I__10015 (
            .O(N__44479),
            .I(N__44472));
    InMux I__10014 (
            .O(N__44478),
            .I(N__44469));
    LocalMux I__10013 (
            .O(N__44475),
            .I(N__44464));
    LocalMux I__10012 (
            .O(N__44472),
            .I(N__44464));
    LocalMux I__10011 (
            .O(N__44469),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv12 I__10010 (
            .O(N__44464),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__10009 (
            .O(N__44459),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__10008 (
            .O(N__44456),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__10007 (
            .O(N__44453),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__10006 (
            .O(N__44450),
            .I(N__44445));
    InMux I__10005 (
            .O(N__44449),
            .I(N__44440));
    InMux I__10004 (
            .O(N__44448),
            .I(N__44440));
    LocalMux I__10003 (
            .O(N__44445),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    LocalMux I__10002 (
            .O(N__44440),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__10001 (
            .O(N__44435),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    CascadeMux I__10000 (
            .O(N__44432),
            .I(N__44427));
    InMux I__9999 (
            .O(N__44431),
            .I(N__44424));
    InMux I__9998 (
            .O(N__44430),
            .I(N__44419));
    InMux I__9997 (
            .O(N__44427),
            .I(N__44419));
    LocalMux I__9996 (
            .O(N__44424),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__9995 (
            .O(N__44419),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__9994 (
            .O(N__44414),
            .I(bfn_18_14_0_));
    InMux I__9993 (
            .O(N__44411),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__9992 (
            .O(N__44408),
            .I(N__44404));
    InMux I__9991 (
            .O(N__44407),
            .I(N__44401));
    LocalMux I__9990 (
            .O(N__44404),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__9989 (
            .O(N__44401),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__9988 (
            .O(N__44396),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__9987 (
            .O(N__44393),
            .I(N__44389));
    InMux I__9986 (
            .O(N__44392),
            .I(N__44386));
    LocalMux I__9985 (
            .O(N__44389),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__9984 (
            .O(N__44386),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__9983 (
            .O(N__44381),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__9982 (
            .O(N__44378),
            .I(N__44375));
    LocalMux I__9981 (
            .O(N__44375),
            .I(N__44371));
    InMux I__9980 (
            .O(N__44374),
            .I(N__44368));
    Span4Mux_h I__9979 (
            .O(N__44371),
            .I(N__44365));
    LocalMux I__9978 (
            .O(N__44368),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__9977 (
            .O(N__44365),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__9976 (
            .O(N__44360),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__9975 (
            .O(N__44357),
            .I(N__44353));
    InMux I__9974 (
            .O(N__44356),
            .I(N__44350));
    LocalMux I__9973 (
            .O(N__44353),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__9972 (
            .O(N__44350),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__9971 (
            .O(N__44345),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__9970 (
            .O(N__44342),
            .I(N__44338));
    InMux I__9969 (
            .O(N__44341),
            .I(N__44335));
    LocalMux I__9968 (
            .O(N__44338),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__9967 (
            .O(N__44335),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__9966 (
            .O(N__44330),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__9965 (
            .O(N__44327),
            .I(N__44323));
    InMux I__9964 (
            .O(N__44326),
            .I(N__44320));
    LocalMux I__9963 (
            .O(N__44323),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__9962 (
            .O(N__44320),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__9961 (
            .O(N__44315),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__9960 (
            .O(N__44312),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__9959 (
            .O(N__44309),
            .I(bfn_18_13_0_));
    InMux I__9958 (
            .O(N__44306),
            .I(N__44303));
    LocalMux I__9957 (
            .O(N__44303),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    CascadeMux I__9956 (
            .O(N__44300),
            .I(N__44297));
    InMux I__9955 (
            .O(N__44297),
            .I(N__44293));
    CascadeMux I__9954 (
            .O(N__44296),
            .I(N__44289));
    LocalMux I__9953 (
            .O(N__44293),
            .I(N__44286));
    InMux I__9952 (
            .O(N__44292),
            .I(N__44283));
    InMux I__9951 (
            .O(N__44289),
            .I(N__44280));
    Span12Mux_h I__9950 (
            .O(N__44286),
            .I(N__44277));
    LocalMux I__9949 (
            .O(N__44283),
            .I(N__44274));
    LocalMux I__9948 (
            .O(N__44280),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv12 I__9947 (
            .O(N__44277),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv12 I__9946 (
            .O(N__44274),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__9945 (
            .O(N__44267),
            .I(N__44263));
    InMux I__9944 (
            .O(N__44266),
            .I(N__44260));
    LocalMux I__9943 (
            .O(N__44263),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__9942 (
            .O(N__44260),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__9941 (
            .O(N__44255),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__9940 (
            .O(N__44252),
            .I(N__44249));
    InMux I__9939 (
            .O(N__44249),
            .I(N__44246));
    LocalMux I__9938 (
            .O(N__44246),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ));
    InMux I__9937 (
            .O(N__44243),
            .I(N__44239));
    InMux I__9936 (
            .O(N__44242),
            .I(N__44236));
    LocalMux I__9935 (
            .O(N__44239),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__9934 (
            .O(N__44236),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__9933 (
            .O(N__44231),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__9932 (
            .O(N__44228),
            .I(N__44224));
    InMux I__9931 (
            .O(N__44227),
            .I(N__44221));
    LocalMux I__9930 (
            .O(N__44224),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__9929 (
            .O(N__44221),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__9928 (
            .O(N__44216),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__9927 (
            .O(N__44213),
            .I(N__44209));
    InMux I__9926 (
            .O(N__44212),
            .I(N__44206));
    LocalMux I__9925 (
            .O(N__44209),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__9924 (
            .O(N__44206),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__9923 (
            .O(N__44201),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__9922 (
            .O(N__44198),
            .I(N__44194));
    InMux I__9921 (
            .O(N__44197),
            .I(N__44191));
    LocalMux I__9920 (
            .O(N__44194),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__9919 (
            .O(N__44191),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__9918 (
            .O(N__44186),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__9917 (
            .O(N__44183),
            .I(N__44179));
    InMux I__9916 (
            .O(N__44182),
            .I(N__44176));
    LocalMux I__9915 (
            .O(N__44179),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__9914 (
            .O(N__44176),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__9913 (
            .O(N__44171),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__9912 (
            .O(N__44168),
            .I(N__44164));
    InMux I__9911 (
            .O(N__44167),
            .I(N__44161));
    LocalMux I__9910 (
            .O(N__44164),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__9909 (
            .O(N__44161),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__9908 (
            .O(N__44156),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__9907 (
            .O(N__44153),
            .I(N__44149));
    InMux I__9906 (
            .O(N__44152),
            .I(N__44146));
    LocalMux I__9905 (
            .O(N__44149),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__9904 (
            .O(N__44146),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__9903 (
            .O(N__44141),
            .I(bfn_18_12_0_));
    InMux I__9902 (
            .O(N__44138),
            .I(N__44135));
    LocalMux I__9901 (
            .O(N__44135),
            .I(N__44132));
    Span4Mux_v I__9900 (
            .O(N__44132),
            .I(N__44129));
    Odrv4 I__9899 (
            .O(N__44129),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    InMux I__9898 (
            .O(N__44126),
            .I(N__44123));
    LocalMux I__9897 (
            .O(N__44123),
            .I(N__44120));
    Span4Mux_h I__9896 (
            .O(N__44120),
            .I(N__44116));
    InMux I__9895 (
            .O(N__44119),
            .I(N__44113));
    Odrv4 I__9894 (
            .O(N__44116),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    LocalMux I__9893 (
            .O(N__44113),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    CascadeMux I__9892 (
            .O(N__44108),
            .I(elapsed_time_ns_1_RNI68CN9_0_19_cascade_));
    InMux I__9891 (
            .O(N__44105),
            .I(N__44100));
    InMux I__9890 (
            .O(N__44104),
            .I(N__44095));
    InMux I__9889 (
            .O(N__44103),
            .I(N__44095));
    LocalMux I__9888 (
            .O(N__44100),
            .I(N__44091));
    LocalMux I__9887 (
            .O(N__44095),
            .I(N__44088));
    InMux I__9886 (
            .O(N__44094),
            .I(N__44085));
    Span4Mux_v I__9885 (
            .O(N__44091),
            .I(N__44080));
    Span4Mux_h I__9884 (
            .O(N__44088),
            .I(N__44080));
    LocalMux I__9883 (
            .O(N__44085),
            .I(N__44077));
    Odrv4 I__9882 (
            .O(N__44080),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    Odrv4 I__9881 (
            .O(N__44077),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    CascadeMux I__9880 (
            .O(N__44072),
            .I(N__44068));
    InMux I__9879 (
            .O(N__44071),
            .I(N__44063));
    InMux I__9878 (
            .O(N__44068),
            .I(N__44063));
    LocalMux I__9877 (
            .O(N__44063),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__9876 (
            .O(N__44060),
            .I(N__44056));
    InMux I__9875 (
            .O(N__44059),
            .I(N__44052));
    LocalMux I__9874 (
            .O(N__44056),
            .I(N__44049));
    InMux I__9873 (
            .O(N__44055),
            .I(N__44046));
    LocalMux I__9872 (
            .O(N__44052),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    Odrv12 I__9871 (
            .O(N__44049),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    LocalMux I__9870 (
            .O(N__44046),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    InMux I__9869 (
            .O(N__44039),
            .I(N__44036));
    LocalMux I__9868 (
            .O(N__44036),
            .I(N__44032));
    InMux I__9867 (
            .O(N__44035),
            .I(N__44029));
    Span4Mux_v I__9866 (
            .O(N__44032),
            .I(N__44022));
    LocalMux I__9865 (
            .O(N__44029),
            .I(N__44022));
    InMux I__9864 (
            .O(N__44028),
            .I(N__44017));
    InMux I__9863 (
            .O(N__44027),
            .I(N__44017));
    Odrv4 I__9862 (
            .O(N__44022),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    LocalMux I__9861 (
            .O(N__44017),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    InMux I__9860 (
            .O(N__44012),
            .I(N__44009));
    LocalMux I__9859 (
            .O(N__44009),
            .I(N__44006));
    Odrv4 I__9858 (
            .O(N__44006),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__9857 (
            .O(N__44003),
            .I(N__43997));
    InMux I__9856 (
            .O(N__44002),
            .I(N__43997));
    LocalMux I__9855 (
            .O(N__43997),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__9854 (
            .O(N__43994),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    InMux I__9853 (
            .O(N__43991),
            .I(N__43988));
    LocalMux I__9852 (
            .O(N__43988),
            .I(N__43985));
    Span4Mux_h I__9851 (
            .O(N__43985),
            .I(N__43981));
    InMux I__9850 (
            .O(N__43984),
            .I(N__43978));
    Odrv4 I__9849 (
            .O(N__43981),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__9848 (
            .O(N__43978),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    InMux I__9847 (
            .O(N__43973),
            .I(N__43967));
    InMux I__9846 (
            .O(N__43972),
            .I(N__43967));
    LocalMux I__9845 (
            .O(N__43967),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ));
    InMux I__9844 (
            .O(N__43964),
            .I(N__43960));
    InMux I__9843 (
            .O(N__43963),
            .I(N__43957));
    LocalMux I__9842 (
            .O(N__43960),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ));
    LocalMux I__9841 (
            .O(N__43957),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ));
    InMux I__9840 (
            .O(N__43952),
            .I(N__43949));
    LocalMux I__9839 (
            .O(N__43949),
            .I(N__43946));
    Span4Mux_v I__9838 (
            .O(N__43946),
            .I(N__43943));
    Odrv4 I__9837 (
            .O(N__43943),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ));
    InMux I__9836 (
            .O(N__43940),
            .I(N__43935));
    InMux I__9835 (
            .O(N__43939),
            .I(N__43932));
    CascadeMux I__9834 (
            .O(N__43938),
            .I(N__43929));
    LocalMux I__9833 (
            .O(N__43935),
            .I(N__43926));
    LocalMux I__9832 (
            .O(N__43932),
            .I(N__43923));
    InMux I__9831 (
            .O(N__43929),
            .I(N__43920));
    Span4Mux_v I__9830 (
            .O(N__43926),
            .I(N__43916));
    Span4Mux_h I__9829 (
            .O(N__43923),
            .I(N__43913));
    LocalMux I__9828 (
            .O(N__43920),
            .I(N__43910));
    InMux I__9827 (
            .O(N__43919),
            .I(N__43907));
    Span4Mux_v I__9826 (
            .O(N__43916),
            .I(N__43904));
    Span4Mux_v I__9825 (
            .O(N__43913),
            .I(N__43901));
    Span4Mux_h I__9824 (
            .O(N__43910),
            .I(N__43898));
    LocalMux I__9823 (
            .O(N__43907),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    Odrv4 I__9822 (
            .O(N__43904),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    Odrv4 I__9821 (
            .O(N__43901),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    Odrv4 I__9820 (
            .O(N__43898),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__9819 (
            .O(N__43889),
            .I(N__43886));
    LocalMux I__9818 (
            .O(N__43886),
            .I(N__43882));
    InMux I__9817 (
            .O(N__43885),
            .I(N__43878));
    Span4Mux_v I__9816 (
            .O(N__43882),
            .I(N__43875));
    InMux I__9815 (
            .O(N__43881),
            .I(N__43872));
    LocalMux I__9814 (
            .O(N__43878),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    Odrv4 I__9813 (
            .O(N__43875),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    LocalMux I__9812 (
            .O(N__43872),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    InMux I__9811 (
            .O(N__43865),
            .I(N__43862));
    LocalMux I__9810 (
            .O(N__43862),
            .I(N__43858));
    InMux I__9809 (
            .O(N__43861),
            .I(N__43855));
    Span4Mux_v I__9808 (
            .O(N__43858),
            .I(N__43851));
    LocalMux I__9807 (
            .O(N__43855),
            .I(N__43848));
    InMux I__9806 (
            .O(N__43854),
            .I(N__43845));
    Odrv4 I__9805 (
            .O(N__43851),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv12 I__9804 (
            .O(N__43848),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__9803 (
            .O(N__43845),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    CascadeMux I__9802 (
            .O(N__43838),
            .I(N__43834));
    InMux I__9801 (
            .O(N__43837),
            .I(N__43831));
    InMux I__9800 (
            .O(N__43834),
            .I(N__43828));
    LocalMux I__9799 (
            .O(N__43831),
            .I(N__43825));
    LocalMux I__9798 (
            .O(N__43828),
            .I(N__43821));
    Span4Mux_v I__9797 (
            .O(N__43825),
            .I(N__43818));
    InMux I__9796 (
            .O(N__43824),
            .I(N__43815));
    Span4Mux_v I__9795 (
            .O(N__43821),
            .I(N__43812));
    Odrv4 I__9794 (
            .O(N__43818),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__9793 (
            .O(N__43815),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__9792 (
            .O(N__43812),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    CEMux I__9791 (
            .O(N__43805),
            .I(N__43802));
    LocalMux I__9790 (
            .O(N__43802),
            .I(N__43797));
    CEMux I__9789 (
            .O(N__43801),
            .I(N__43794));
    CEMux I__9788 (
            .O(N__43800),
            .I(N__43789));
    Span4Mux_h I__9787 (
            .O(N__43797),
            .I(N__43784));
    LocalMux I__9786 (
            .O(N__43794),
            .I(N__43784));
    CEMux I__9785 (
            .O(N__43793),
            .I(N__43781));
    CEMux I__9784 (
            .O(N__43792),
            .I(N__43778));
    LocalMux I__9783 (
            .O(N__43789),
            .I(N__43775));
    Span4Mux_v I__9782 (
            .O(N__43784),
            .I(N__43772));
    LocalMux I__9781 (
            .O(N__43781),
            .I(N__43769));
    LocalMux I__9780 (
            .O(N__43778),
            .I(N__43766));
    Span4Mux_h I__9779 (
            .O(N__43775),
            .I(N__43763));
    Span4Mux_h I__9778 (
            .O(N__43772),
            .I(N__43758));
    Span4Mux_h I__9777 (
            .O(N__43769),
            .I(N__43758));
    Span4Mux_h I__9776 (
            .O(N__43766),
            .I(N__43755));
    Odrv4 I__9775 (
            .O(N__43763),
            .I(\delay_measurement_inst.delay_hc_timer.N_198_i ));
    Odrv4 I__9774 (
            .O(N__43758),
            .I(\delay_measurement_inst.delay_hc_timer.N_198_i ));
    Odrv4 I__9773 (
            .O(N__43755),
            .I(\delay_measurement_inst.delay_hc_timer.N_198_i ));
    InMux I__9772 (
            .O(N__43748),
            .I(N__43745));
    LocalMux I__9771 (
            .O(N__43745),
            .I(N__43741));
    InMux I__9770 (
            .O(N__43744),
            .I(N__43737));
    Span12Mux_h I__9769 (
            .O(N__43741),
            .I(N__43734));
    InMux I__9768 (
            .O(N__43740),
            .I(N__43731));
    LocalMux I__9767 (
            .O(N__43737),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv12 I__9766 (
            .O(N__43734),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    LocalMux I__9765 (
            .O(N__43731),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    InMux I__9764 (
            .O(N__43724),
            .I(N__43721));
    LocalMux I__9763 (
            .O(N__43721),
            .I(N__43717));
    InMux I__9762 (
            .O(N__43720),
            .I(N__43713));
    Span4Mux_v I__9761 (
            .O(N__43717),
            .I(N__43710));
    InMux I__9760 (
            .O(N__43716),
            .I(N__43707));
    LocalMux I__9759 (
            .O(N__43713),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    Odrv4 I__9758 (
            .O(N__43710),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    LocalMux I__9757 (
            .O(N__43707),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    InMux I__9756 (
            .O(N__43700),
            .I(N__43697));
    LocalMux I__9755 (
            .O(N__43697),
            .I(N__43693));
    InMux I__9754 (
            .O(N__43696),
            .I(N__43689));
    Span4Mux_v I__9753 (
            .O(N__43693),
            .I(N__43686));
    InMux I__9752 (
            .O(N__43692),
            .I(N__43683));
    LocalMux I__9751 (
            .O(N__43689),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    Odrv4 I__9750 (
            .O(N__43686),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    LocalMux I__9749 (
            .O(N__43683),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    CascadeMux I__9748 (
            .O(N__43676),
            .I(N__43673));
    InMux I__9747 (
            .O(N__43673),
            .I(N__43670));
    LocalMux I__9746 (
            .O(N__43670),
            .I(N__43667));
    Span4Mux_v I__9745 (
            .O(N__43667),
            .I(N__43664));
    Odrv4 I__9744 (
            .O(N__43664),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    InMux I__9743 (
            .O(N__43661),
            .I(N__43658));
    LocalMux I__9742 (
            .O(N__43658),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__9741 (
            .O(N__43655),
            .I(N__43652));
    InMux I__9740 (
            .O(N__43652),
            .I(N__43649));
    LocalMux I__9739 (
            .O(N__43649),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__9738 (
            .O(N__43646),
            .I(N__43643));
    LocalMux I__9737 (
            .O(N__43643),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    CascadeMux I__9736 (
            .O(N__43640),
            .I(N__43637));
    InMux I__9735 (
            .O(N__43637),
            .I(N__43634));
    LocalMux I__9734 (
            .O(N__43634),
            .I(N__43631));
    Span4Mux_h I__9733 (
            .O(N__43631),
            .I(N__43628));
    Span4Mux_v I__9732 (
            .O(N__43628),
            .I(N__43625));
    Odrv4 I__9731 (
            .O(N__43625),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__9730 (
            .O(N__43622),
            .I(N__43619));
    LocalMux I__9729 (
            .O(N__43619),
            .I(N__43616));
    Span4Mux_v I__9728 (
            .O(N__43616),
            .I(N__43613));
    Odrv4 I__9727 (
            .O(N__43613),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__9726 (
            .O(N__43610),
            .I(N__43607));
    InMux I__9725 (
            .O(N__43607),
            .I(N__43604));
    LocalMux I__9724 (
            .O(N__43604),
            .I(N__43601));
    Span12Mux_s11_v I__9723 (
            .O(N__43601),
            .I(N__43598));
    Odrv12 I__9722 (
            .O(N__43598),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__9721 (
            .O(N__43595),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__9720 (
            .O(N__43592),
            .I(N__43586));
    InMux I__9719 (
            .O(N__43591),
            .I(N__43583));
    CascadeMux I__9718 (
            .O(N__43590),
            .I(N__43568));
    CascadeMux I__9717 (
            .O(N__43589),
            .I(N__43563));
    LocalMux I__9716 (
            .O(N__43586),
            .I(N__43546));
    LocalMux I__9715 (
            .O(N__43583),
            .I(N__43546));
    InMux I__9714 (
            .O(N__43582),
            .I(N__43543));
    InMux I__9713 (
            .O(N__43581),
            .I(N__43532));
    InMux I__9712 (
            .O(N__43580),
            .I(N__43532));
    InMux I__9711 (
            .O(N__43579),
            .I(N__43532));
    InMux I__9710 (
            .O(N__43578),
            .I(N__43532));
    InMux I__9709 (
            .O(N__43577),
            .I(N__43532));
    InMux I__9708 (
            .O(N__43576),
            .I(N__43529));
    InMux I__9707 (
            .O(N__43575),
            .I(N__43520));
    InMux I__9706 (
            .O(N__43574),
            .I(N__43520));
    InMux I__9705 (
            .O(N__43573),
            .I(N__43520));
    InMux I__9704 (
            .O(N__43572),
            .I(N__43520));
    InMux I__9703 (
            .O(N__43571),
            .I(N__43517));
    InMux I__9702 (
            .O(N__43568),
            .I(N__43512));
    InMux I__9701 (
            .O(N__43567),
            .I(N__43501));
    InMux I__9700 (
            .O(N__43566),
            .I(N__43501));
    InMux I__9699 (
            .O(N__43563),
            .I(N__43501));
    InMux I__9698 (
            .O(N__43562),
            .I(N__43501));
    InMux I__9697 (
            .O(N__43561),
            .I(N__43501));
    InMux I__9696 (
            .O(N__43560),
            .I(N__43496));
    InMux I__9695 (
            .O(N__43559),
            .I(N__43496));
    InMux I__9694 (
            .O(N__43558),
            .I(N__43491));
    InMux I__9693 (
            .O(N__43557),
            .I(N__43491));
    InMux I__9692 (
            .O(N__43556),
            .I(N__43488));
    InMux I__9691 (
            .O(N__43555),
            .I(N__43477));
    InMux I__9690 (
            .O(N__43554),
            .I(N__43477));
    InMux I__9689 (
            .O(N__43553),
            .I(N__43477));
    InMux I__9688 (
            .O(N__43552),
            .I(N__43477));
    InMux I__9687 (
            .O(N__43551),
            .I(N__43477));
    Span4Mux_v I__9686 (
            .O(N__43546),
            .I(N__43466));
    LocalMux I__9685 (
            .O(N__43543),
            .I(N__43466));
    LocalMux I__9684 (
            .O(N__43532),
            .I(N__43466));
    LocalMux I__9683 (
            .O(N__43529),
            .I(N__43466));
    LocalMux I__9682 (
            .O(N__43520),
            .I(N__43466));
    LocalMux I__9681 (
            .O(N__43517),
            .I(N__43463));
    InMux I__9680 (
            .O(N__43516),
            .I(N__43458));
    InMux I__9679 (
            .O(N__43515),
            .I(N__43458));
    LocalMux I__9678 (
            .O(N__43512),
            .I(N__43451));
    LocalMux I__9677 (
            .O(N__43501),
            .I(N__43451));
    LocalMux I__9676 (
            .O(N__43496),
            .I(N__43451));
    LocalMux I__9675 (
            .O(N__43491),
            .I(N__43442));
    LocalMux I__9674 (
            .O(N__43488),
            .I(N__43442));
    LocalMux I__9673 (
            .O(N__43477),
            .I(N__43442));
    Span4Mux_h I__9672 (
            .O(N__43466),
            .I(N__43442));
    Span4Mux_h I__9671 (
            .O(N__43463),
            .I(N__43439));
    LocalMux I__9670 (
            .O(N__43458),
            .I(N__43436));
    Span4Mux_h I__9669 (
            .O(N__43451),
            .I(N__43433));
    Span4Mux_v I__9668 (
            .O(N__43442),
            .I(N__43430));
    Span4Mux_h I__9667 (
            .O(N__43439),
            .I(N__43427));
    Span12Mux_h I__9666 (
            .O(N__43436),
            .I(N__43424));
    Span4Mux_v I__9665 (
            .O(N__43433),
            .I(N__43419));
    Span4Mux_v I__9664 (
            .O(N__43430),
            .I(N__43419));
    Odrv4 I__9663 (
            .O(N__43427),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv12 I__9662 (
            .O(N__43424),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__9661 (
            .O(N__43419),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    CascadeMux I__9660 (
            .O(N__43412),
            .I(N__43409));
    InMux I__9659 (
            .O(N__43409),
            .I(N__43406));
    LocalMux I__9658 (
            .O(N__43406),
            .I(N__43403));
    Span4Mux_v I__9657 (
            .O(N__43403),
            .I(N__43400));
    Odrv4 I__9656 (
            .O(N__43400),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt20 ));
    InMux I__9655 (
            .O(N__43397),
            .I(N__43394));
    LocalMux I__9654 (
            .O(N__43394),
            .I(N__43391));
    Odrv12 I__9653 (
            .O(N__43391),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__9652 (
            .O(N__43388),
            .I(N__43385));
    InMux I__9651 (
            .O(N__43385),
            .I(N__43382));
    LocalMux I__9650 (
            .O(N__43382),
            .I(N__43379));
    Span4Mux_v I__9649 (
            .O(N__43379),
            .I(N__43376));
    Odrv4 I__9648 (
            .O(N__43376),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__9647 (
            .O(N__43373),
            .I(N__43370));
    LocalMux I__9646 (
            .O(N__43370),
            .I(N__43367));
    Span4Mux_v I__9645 (
            .O(N__43367),
            .I(N__43364));
    Odrv4 I__9644 (
            .O(N__43364),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    CascadeMux I__9643 (
            .O(N__43361),
            .I(N__43358));
    InMux I__9642 (
            .O(N__43358),
            .I(N__43355));
    LocalMux I__9641 (
            .O(N__43355),
            .I(N__43352));
    Span4Mux_v I__9640 (
            .O(N__43352),
            .I(N__43349));
    Odrv4 I__9639 (
            .O(N__43349),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__9638 (
            .O(N__43346),
            .I(N__43343));
    LocalMux I__9637 (
            .O(N__43343),
            .I(N__43340));
    Odrv12 I__9636 (
            .O(N__43340),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    CascadeMux I__9635 (
            .O(N__43337),
            .I(N__43334));
    InMux I__9634 (
            .O(N__43334),
            .I(N__43331));
    LocalMux I__9633 (
            .O(N__43331),
            .I(N__43328));
    Odrv4 I__9632 (
            .O(N__43328),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__9631 (
            .O(N__43325),
            .I(N__43322));
    LocalMux I__9630 (
            .O(N__43322),
            .I(N__43319));
    Odrv12 I__9629 (
            .O(N__43319),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    CascadeMux I__9628 (
            .O(N__43316),
            .I(N__43313));
    InMux I__9627 (
            .O(N__43313),
            .I(N__43310));
    LocalMux I__9626 (
            .O(N__43310),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    CascadeMux I__9625 (
            .O(N__43307),
            .I(N__43304));
    InMux I__9624 (
            .O(N__43304),
            .I(N__43301));
    LocalMux I__9623 (
            .O(N__43301),
            .I(N__43298));
    Span4Mux_v I__9622 (
            .O(N__43298),
            .I(N__43295));
    Odrv4 I__9621 (
            .O(N__43295),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__9620 (
            .O(N__43292),
            .I(N__43289));
    LocalMux I__9619 (
            .O(N__43289),
            .I(N__43286));
    Odrv12 I__9618 (
            .O(N__43286),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    CascadeMux I__9617 (
            .O(N__43283),
            .I(N__43280));
    InMux I__9616 (
            .O(N__43280),
            .I(N__43277));
    LocalMux I__9615 (
            .O(N__43277),
            .I(N__43274));
    Span4Mux_v I__9614 (
            .O(N__43274),
            .I(N__43271));
    Odrv4 I__9613 (
            .O(N__43271),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    CascadeMux I__9612 (
            .O(N__43268),
            .I(N__43265));
    InMux I__9611 (
            .O(N__43265),
            .I(N__43262));
    LocalMux I__9610 (
            .O(N__43262),
            .I(N__43259));
    Span4Mux_v I__9609 (
            .O(N__43259),
            .I(N__43256));
    Odrv4 I__9608 (
            .O(N__43256),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__9607 (
            .O(N__43253),
            .I(N__43250));
    LocalMux I__9606 (
            .O(N__43250),
            .I(N__43247));
    Odrv12 I__9605 (
            .O(N__43247),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__9604 (
            .O(N__43244),
            .I(N__43241));
    InMux I__9603 (
            .O(N__43241),
            .I(N__43238));
    LocalMux I__9602 (
            .O(N__43238),
            .I(N__43235));
    Odrv12 I__9601 (
            .O(N__43235),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__9600 (
            .O(N__43232),
            .I(N__43229));
    LocalMux I__9599 (
            .O(N__43229),
            .I(N__43226));
    Odrv12 I__9598 (
            .O(N__43226),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__9597 (
            .O(N__43223),
            .I(N__43220));
    InMux I__9596 (
            .O(N__43220),
            .I(N__43217));
    LocalMux I__9595 (
            .O(N__43217),
            .I(N__43214));
    Odrv12 I__9594 (
            .O(N__43214),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__9593 (
            .O(N__43211),
            .I(N__43208));
    InMux I__9592 (
            .O(N__43208),
            .I(N__43205));
    LocalMux I__9591 (
            .O(N__43205),
            .I(N__43202));
    Span4Mux_v I__9590 (
            .O(N__43202),
            .I(N__43199));
    Odrv4 I__9589 (
            .O(N__43199),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__9588 (
            .O(N__43196),
            .I(N__43193));
    LocalMux I__9587 (
            .O(N__43193),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__9586 (
            .O(N__43190),
            .I(N__43187));
    InMux I__9585 (
            .O(N__43187),
            .I(N__43184));
    LocalMux I__9584 (
            .O(N__43184),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__9583 (
            .O(N__43181),
            .I(N__43178));
    LocalMux I__9582 (
            .O(N__43178),
            .I(N__43175));
    Span4Mux_v I__9581 (
            .O(N__43175),
            .I(N__43172));
    Odrv4 I__9580 (
            .O(N__43172),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__9579 (
            .O(N__43169),
            .I(N__43166));
    InMux I__9578 (
            .O(N__43166),
            .I(N__43163));
    LocalMux I__9577 (
            .O(N__43163),
            .I(N__43160));
    Odrv12 I__9576 (
            .O(N__43160),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__9575 (
            .O(N__43157),
            .I(N__43154));
    LocalMux I__9574 (
            .O(N__43154),
            .I(N__43151));
    Odrv12 I__9573 (
            .O(N__43151),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__9572 (
            .O(N__43148),
            .I(N__43145));
    InMux I__9571 (
            .O(N__43145),
            .I(N__43142));
    LocalMux I__9570 (
            .O(N__43142),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__9569 (
            .O(N__43139),
            .I(N__43133));
    InMux I__9568 (
            .O(N__43138),
            .I(N__43130));
    InMux I__9567 (
            .O(N__43137),
            .I(N__43125));
    InMux I__9566 (
            .O(N__43136),
            .I(N__43125));
    InMux I__9565 (
            .O(N__43133),
            .I(N__43122));
    LocalMux I__9564 (
            .O(N__43130),
            .I(N__43119));
    LocalMux I__9563 (
            .O(N__43125),
            .I(N__43116));
    LocalMux I__9562 (
            .O(N__43122),
            .I(N__43113));
    Span4Mux_v I__9561 (
            .O(N__43119),
            .I(N__43108));
    Span4Mux_v I__9560 (
            .O(N__43116),
            .I(N__43108));
    Span4Mux_h I__9559 (
            .O(N__43113),
            .I(N__43105));
    Span4Mux_h I__9558 (
            .O(N__43108),
            .I(N__43102));
    Odrv4 I__9557 (
            .O(N__43105),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__9556 (
            .O(N__43102),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__9555 (
            .O(N__43097),
            .I(N__43094));
    LocalMux I__9554 (
            .O(N__43094),
            .I(N__43091));
    Span4Mux_h I__9553 (
            .O(N__43091),
            .I(N__43086));
    InMux I__9552 (
            .O(N__43090),
            .I(N__43083));
    InMux I__9551 (
            .O(N__43089),
            .I(N__43080));
    Odrv4 I__9550 (
            .O(N__43086),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__9549 (
            .O(N__43083),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__9548 (
            .O(N__43080),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__9547 (
            .O(N__43073),
            .I(N__43070));
    LocalMux I__9546 (
            .O(N__43070),
            .I(N__43065));
    InMux I__9545 (
            .O(N__43069),
            .I(N__43062));
    InMux I__9544 (
            .O(N__43068),
            .I(N__43059));
    Span4Mux_h I__9543 (
            .O(N__43065),
            .I(N__43056));
    LocalMux I__9542 (
            .O(N__43062),
            .I(N__43050));
    LocalMux I__9541 (
            .O(N__43059),
            .I(N__43050));
    Span4Mux_h I__9540 (
            .O(N__43056),
            .I(N__43047));
    InMux I__9539 (
            .O(N__43055),
            .I(N__43044));
    Span4Mux_v I__9538 (
            .O(N__43050),
            .I(N__43041));
    Odrv4 I__9537 (
            .O(N__43047),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    LocalMux I__9536 (
            .O(N__43044),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__9535 (
            .O(N__43041),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    CascadeMux I__9534 (
            .O(N__43034),
            .I(N__43030));
    InMux I__9533 (
            .O(N__43033),
            .I(N__43026));
    InMux I__9532 (
            .O(N__43030),
            .I(N__43023));
    CascadeMux I__9531 (
            .O(N__43029),
            .I(N__43020));
    LocalMux I__9530 (
            .O(N__43026),
            .I(N__43017));
    LocalMux I__9529 (
            .O(N__43023),
            .I(N__43014));
    InMux I__9528 (
            .O(N__43020),
            .I(N__43011));
    Span4Mux_v I__9527 (
            .O(N__43017),
            .I(N__43008));
    Odrv4 I__9526 (
            .O(N__43014),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__9525 (
            .O(N__43011),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__9524 (
            .O(N__43008),
            .I(\current_shift_inst.un4_control_input1_8 ));
    CascadeMux I__9523 (
            .O(N__43001),
            .I(N__42997));
    InMux I__9522 (
            .O(N__43000),
            .I(N__42993));
    InMux I__9521 (
            .O(N__42997),
            .I(N__42990));
    CascadeMux I__9520 (
            .O(N__42996),
            .I(N__42987));
    LocalMux I__9519 (
            .O(N__42993),
            .I(N__42984));
    LocalMux I__9518 (
            .O(N__42990),
            .I(N__42981));
    InMux I__9517 (
            .O(N__42987),
            .I(N__42978));
    Span4Mux_h I__9516 (
            .O(N__42984),
            .I(N__42975));
    Odrv4 I__9515 (
            .O(N__42981),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    LocalMux I__9514 (
            .O(N__42978),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    Odrv4 I__9513 (
            .O(N__42975),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__9512 (
            .O(N__42968),
            .I(N__42965));
    InMux I__9511 (
            .O(N__42965),
            .I(N__42962));
    LocalMux I__9510 (
            .O(N__42962),
            .I(N__42959));
    Span4Mux_v I__9509 (
            .O(N__42959),
            .I(N__42956));
    Odrv4 I__9508 (
            .O(N__42956),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    CascadeMux I__9507 (
            .O(N__42953),
            .I(N__42949));
    InMux I__9506 (
            .O(N__42952),
            .I(N__42945));
    InMux I__9505 (
            .O(N__42949),
            .I(N__42940));
    InMux I__9504 (
            .O(N__42948),
            .I(N__42940));
    LocalMux I__9503 (
            .O(N__42945),
            .I(N__42935));
    LocalMux I__9502 (
            .O(N__42940),
            .I(N__42935));
    Span4Mux_v I__9501 (
            .O(N__42935),
            .I(N__42931));
    InMux I__9500 (
            .O(N__42934),
            .I(N__42928));
    Odrv4 I__9499 (
            .O(N__42931),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__9498 (
            .O(N__42928),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    CascadeMux I__9497 (
            .O(N__42923),
            .I(N__42920));
    InMux I__9496 (
            .O(N__42920),
            .I(N__42917));
    LocalMux I__9495 (
            .O(N__42917),
            .I(N__42914));
    Odrv4 I__9494 (
            .O(N__42914),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    CascadeMux I__9493 (
            .O(N__42911),
            .I(N__42903));
    CascadeMux I__9492 (
            .O(N__42910),
            .I(N__42899));
    CascadeMux I__9491 (
            .O(N__42909),
            .I(N__42884));
    InMux I__9490 (
            .O(N__42908),
            .I(N__42871));
    InMux I__9489 (
            .O(N__42907),
            .I(N__42871));
    InMux I__9488 (
            .O(N__42906),
            .I(N__42866));
    InMux I__9487 (
            .O(N__42903),
            .I(N__42866));
    CascadeMux I__9486 (
            .O(N__42902),
            .I(N__42851));
    InMux I__9485 (
            .O(N__42899),
            .I(N__42848));
    CascadeMux I__9484 (
            .O(N__42898),
            .I(N__42843));
    CascadeMux I__9483 (
            .O(N__42897),
            .I(N__42834));
    CascadeMux I__9482 (
            .O(N__42896),
            .I(N__42828));
    CascadeMux I__9481 (
            .O(N__42895),
            .I(N__42820));
    CascadeMux I__9480 (
            .O(N__42894),
            .I(N__42816));
    CascadeMux I__9479 (
            .O(N__42893),
            .I(N__42812));
    CascadeMux I__9478 (
            .O(N__42892),
            .I(N__42809));
    CascadeMux I__9477 (
            .O(N__42891),
            .I(N__42805));
    CascadeMux I__9476 (
            .O(N__42890),
            .I(N__42801));
    CascadeMux I__9475 (
            .O(N__42889),
            .I(N__42797));
    InMux I__9474 (
            .O(N__42888),
            .I(N__42789));
    InMux I__9473 (
            .O(N__42887),
            .I(N__42773));
    InMux I__9472 (
            .O(N__42884),
            .I(N__42773));
    CascadeMux I__9471 (
            .O(N__42883),
            .I(N__42768));
    CascadeMux I__9470 (
            .O(N__42882),
            .I(N__42765));
    InMux I__9469 (
            .O(N__42881),
            .I(N__42762));
    InMux I__9468 (
            .O(N__42880),
            .I(N__42757));
    InMux I__9467 (
            .O(N__42879),
            .I(N__42757));
    CascadeMux I__9466 (
            .O(N__42878),
            .I(N__42754));
    CascadeMux I__9465 (
            .O(N__42877),
            .I(N__42750));
    CascadeMux I__9464 (
            .O(N__42876),
            .I(N__42746));
    LocalMux I__9463 (
            .O(N__42871),
            .I(N__42740));
    LocalMux I__9462 (
            .O(N__42866),
            .I(N__42740));
    CascadeMux I__9461 (
            .O(N__42865),
            .I(N__42737));
    CascadeMux I__9460 (
            .O(N__42864),
            .I(N__42734));
    CascadeMux I__9459 (
            .O(N__42863),
            .I(N__42731));
    CascadeMux I__9458 (
            .O(N__42862),
            .I(N__42727));
    CascadeMux I__9457 (
            .O(N__42861),
            .I(N__42724));
    InMux I__9456 (
            .O(N__42860),
            .I(N__42713));
    InMux I__9455 (
            .O(N__42859),
            .I(N__42710));
    InMux I__9454 (
            .O(N__42858),
            .I(N__42697));
    InMux I__9453 (
            .O(N__42857),
            .I(N__42697));
    InMux I__9452 (
            .O(N__42856),
            .I(N__42697));
    InMux I__9451 (
            .O(N__42855),
            .I(N__42697));
    InMux I__9450 (
            .O(N__42854),
            .I(N__42697));
    InMux I__9449 (
            .O(N__42851),
            .I(N__42697));
    LocalMux I__9448 (
            .O(N__42848),
            .I(N__42694));
    InMux I__9447 (
            .O(N__42847),
            .I(N__42689));
    InMux I__9446 (
            .O(N__42846),
            .I(N__42689));
    InMux I__9445 (
            .O(N__42843),
            .I(N__42674));
    InMux I__9444 (
            .O(N__42842),
            .I(N__42674));
    InMux I__9443 (
            .O(N__42841),
            .I(N__42674));
    InMux I__9442 (
            .O(N__42840),
            .I(N__42674));
    InMux I__9441 (
            .O(N__42839),
            .I(N__42674));
    InMux I__9440 (
            .O(N__42838),
            .I(N__42674));
    InMux I__9439 (
            .O(N__42837),
            .I(N__42674));
    InMux I__9438 (
            .O(N__42834),
            .I(N__42659));
    InMux I__9437 (
            .O(N__42833),
            .I(N__42659));
    InMux I__9436 (
            .O(N__42832),
            .I(N__42659));
    InMux I__9435 (
            .O(N__42831),
            .I(N__42659));
    InMux I__9434 (
            .O(N__42828),
            .I(N__42659));
    InMux I__9433 (
            .O(N__42827),
            .I(N__42659));
    InMux I__9432 (
            .O(N__42826),
            .I(N__42659));
    InMux I__9431 (
            .O(N__42825),
            .I(N__42656));
    InMux I__9430 (
            .O(N__42824),
            .I(N__42641));
    InMux I__9429 (
            .O(N__42823),
            .I(N__42641));
    InMux I__9428 (
            .O(N__42820),
            .I(N__42641));
    InMux I__9427 (
            .O(N__42819),
            .I(N__42641));
    InMux I__9426 (
            .O(N__42816),
            .I(N__42641));
    InMux I__9425 (
            .O(N__42815),
            .I(N__42641));
    InMux I__9424 (
            .O(N__42812),
            .I(N__42641));
    InMux I__9423 (
            .O(N__42809),
            .I(N__42624));
    InMux I__9422 (
            .O(N__42808),
            .I(N__42624));
    InMux I__9421 (
            .O(N__42805),
            .I(N__42624));
    InMux I__9420 (
            .O(N__42804),
            .I(N__42624));
    InMux I__9419 (
            .O(N__42801),
            .I(N__42624));
    InMux I__9418 (
            .O(N__42800),
            .I(N__42624));
    InMux I__9417 (
            .O(N__42797),
            .I(N__42624));
    InMux I__9416 (
            .O(N__42796),
            .I(N__42624));
    CascadeMux I__9415 (
            .O(N__42795),
            .I(N__42621));
    CascadeMux I__9414 (
            .O(N__42794),
            .I(N__42617));
    CascadeMux I__9413 (
            .O(N__42793),
            .I(N__42613));
    CascadeMux I__9412 (
            .O(N__42792),
            .I(N__42609));
    LocalMux I__9411 (
            .O(N__42789),
            .I(N__42602));
    InMux I__9410 (
            .O(N__42788),
            .I(N__42595));
    InMux I__9409 (
            .O(N__42787),
            .I(N__42595));
    InMux I__9408 (
            .O(N__42786),
            .I(N__42595));
    CascadeMux I__9407 (
            .O(N__42785),
            .I(N__42592));
    CascadeMux I__9406 (
            .O(N__42784),
            .I(N__42588));
    CascadeMux I__9405 (
            .O(N__42783),
            .I(N__42584));
    CascadeMux I__9404 (
            .O(N__42782),
            .I(N__42580));
    CascadeMux I__9403 (
            .O(N__42781),
            .I(N__42576));
    CascadeMux I__9402 (
            .O(N__42780),
            .I(N__42572));
    CascadeMux I__9401 (
            .O(N__42779),
            .I(N__42568));
    CascadeMux I__9400 (
            .O(N__42778),
            .I(N__42564));
    LocalMux I__9399 (
            .O(N__42773),
            .I(N__42560));
    InMux I__9398 (
            .O(N__42772),
            .I(N__42553));
    InMux I__9397 (
            .O(N__42771),
            .I(N__42553));
    InMux I__9396 (
            .O(N__42768),
            .I(N__42553));
    InMux I__9395 (
            .O(N__42765),
            .I(N__42550));
    LocalMux I__9394 (
            .O(N__42762),
            .I(N__42545));
    LocalMux I__9393 (
            .O(N__42757),
            .I(N__42545));
    InMux I__9392 (
            .O(N__42754),
            .I(N__42532));
    InMux I__9391 (
            .O(N__42753),
            .I(N__42532));
    InMux I__9390 (
            .O(N__42750),
            .I(N__42532));
    InMux I__9389 (
            .O(N__42749),
            .I(N__42532));
    InMux I__9388 (
            .O(N__42746),
            .I(N__42532));
    InMux I__9387 (
            .O(N__42745),
            .I(N__42532));
    Span4Mux_v I__9386 (
            .O(N__42740),
            .I(N__42529));
    InMux I__9385 (
            .O(N__42737),
            .I(N__42524));
    InMux I__9384 (
            .O(N__42734),
            .I(N__42524));
    InMux I__9383 (
            .O(N__42731),
            .I(N__42513));
    InMux I__9382 (
            .O(N__42730),
            .I(N__42513));
    InMux I__9381 (
            .O(N__42727),
            .I(N__42513));
    InMux I__9380 (
            .O(N__42724),
            .I(N__42513));
    InMux I__9379 (
            .O(N__42723),
            .I(N__42513));
    CascadeMux I__9378 (
            .O(N__42722),
            .I(N__42508));
    CascadeMux I__9377 (
            .O(N__42721),
            .I(N__42505));
    CascadeMux I__9376 (
            .O(N__42720),
            .I(N__42499));
    CascadeMux I__9375 (
            .O(N__42719),
            .I(N__42495));
    CascadeMux I__9374 (
            .O(N__42718),
            .I(N__42491));
    CascadeMux I__9373 (
            .O(N__42717),
            .I(N__42487));
    CascadeMux I__9372 (
            .O(N__42716),
            .I(N__42483));
    LocalMux I__9371 (
            .O(N__42713),
            .I(N__42475));
    LocalMux I__9370 (
            .O(N__42710),
            .I(N__42475));
    LocalMux I__9369 (
            .O(N__42697),
            .I(N__42475));
    Span4Mux_v I__9368 (
            .O(N__42694),
            .I(N__42460));
    LocalMux I__9367 (
            .O(N__42689),
            .I(N__42460));
    LocalMux I__9366 (
            .O(N__42674),
            .I(N__42460));
    LocalMux I__9365 (
            .O(N__42659),
            .I(N__42460));
    LocalMux I__9364 (
            .O(N__42656),
            .I(N__42460));
    LocalMux I__9363 (
            .O(N__42641),
            .I(N__42460));
    LocalMux I__9362 (
            .O(N__42624),
            .I(N__42460));
    InMux I__9361 (
            .O(N__42621),
            .I(N__42443));
    InMux I__9360 (
            .O(N__42620),
            .I(N__42443));
    InMux I__9359 (
            .O(N__42617),
            .I(N__42443));
    InMux I__9358 (
            .O(N__42616),
            .I(N__42443));
    InMux I__9357 (
            .O(N__42613),
            .I(N__42443));
    InMux I__9356 (
            .O(N__42612),
            .I(N__42443));
    InMux I__9355 (
            .O(N__42609),
            .I(N__42443));
    InMux I__9354 (
            .O(N__42608),
            .I(N__42443));
    CascadeMux I__9353 (
            .O(N__42607),
            .I(N__42440));
    CascadeMux I__9352 (
            .O(N__42606),
            .I(N__42436));
    CascadeMux I__9351 (
            .O(N__42605),
            .I(N__42432));
    Span4Mux_v I__9350 (
            .O(N__42602),
            .I(N__42426));
    LocalMux I__9349 (
            .O(N__42595),
            .I(N__42426));
    InMux I__9348 (
            .O(N__42592),
            .I(N__42423));
    InMux I__9347 (
            .O(N__42591),
            .I(N__42408));
    InMux I__9346 (
            .O(N__42588),
            .I(N__42408));
    InMux I__9345 (
            .O(N__42587),
            .I(N__42408));
    InMux I__9344 (
            .O(N__42584),
            .I(N__42408));
    InMux I__9343 (
            .O(N__42583),
            .I(N__42408));
    InMux I__9342 (
            .O(N__42580),
            .I(N__42408));
    InMux I__9341 (
            .O(N__42579),
            .I(N__42408));
    InMux I__9340 (
            .O(N__42576),
            .I(N__42391));
    InMux I__9339 (
            .O(N__42575),
            .I(N__42391));
    InMux I__9338 (
            .O(N__42572),
            .I(N__42391));
    InMux I__9337 (
            .O(N__42571),
            .I(N__42391));
    InMux I__9336 (
            .O(N__42568),
            .I(N__42391));
    InMux I__9335 (
            .O(N__42567),
            .I(N__42391));
    InMux I__9334 (
            .O(N__42564),
            .I(N__42391));
    InMux I__9333 (
            .O(N__42563),
            .I(N__42391));
    Span4Mux_v I__9332 (
            .O(N__42560),
            .I(N__42380));
    LocalMux I__9331 (
            .O(N__42553),
            .I(N__42380));
    LocalMux I__9330 (
            .O(N__42550),
            .I(N__42380));
    Span4Mux_h I__9329 (
            .O(N__42545),
            .I(N__42380));
    LocalMux I__9328 (
            .O(N__42532),
            .I(N__42380));
    Span4Mux_h I__9327 (
            .O(N__42529),
            .I(N__42377));
    LocalMux I__9326 (
            .O(N__42524),
            .I(N__42372));
    LocalMux I__9325 (
            .O(N__42513),
            .I(N__42372));
    InMux I__9324 (
            .O(N__42512),
            .I(N__42359));
    InMux I__9323 (
            .O(N__42511),
            .I(N__42359));
    InMux I__9322 (
            .O(N__42508),
            .I(N__42359));
    InMux I__9321 (
            .O(N__42505),
            .I(N__42359));
    InMux I__9320 (
            .O(N__42504),
            .I(N__42359));
    InMux I__9319 (
            .O(N__42503),
            .I(N__42359));
    InMux I__9318 (
            .O(N__42502),
            .I(N__42352));
    InMux I__9317 (
            .O(N__42499),
            .I(N__42352));
    InMux I__9316 (
            .O(N__42498),
            .I(N__42352));
    InMux I__9315 (
            .O(N__42495),
            .I(N__42335));
    InMux I__9314 (
            .O(N__42494),
            .I(N__42335));
    InMux I__9313 (
            .O(N__42491),
            .I(N__42335));
    InMux I__9312 (
            .O(N__42490),
            .I(N__42335));
    InMux I__9311 (
            .O(N__42487),
            .I(N__42335));
    InMux I__9310 (
            .O(N__42486),
            .I(N__42335));
    InMux I__9309 (
            .O(N__42483),
            .I(N__42335));
    InMux I__9308 (
            .O(N__42482),
            .I(N__42335));
    Span4Mux_h I__9307 (
            .O(N__42475),
            .I(N__42328));
    Span4Mux_v I__9306 (
            .O(N__42460),
            .I(N__42328));
    LocalMux I__9305 (
            .O(N__42443),
            .I(N__42328));
    InMux I__9304 (
            .O(N__42440),
            .I(N__42315));
    InMux I__9303 (
            .O(N__42439),
            .I(N__42315));
    InMux I__9302 (
            .O(N__42436),
            .I(N__42315));
    InMux I__9301 (
            .O(N__42435),
            .I(N__42315));
    InMux I__9300 (
            .O(N__42432),
            .I(N__42315));
    InMux I__9299 (
            .O(N__42431),
            .I(N__42315));
    Span4Mux_h I__9298 (
            .O(N__42426),
            .I(N__42304));
    LocalMux I__9297 (
            .O(N__42423),
            .I(N__42304));
    LocalMux I__9296 (
            .O(N__42408),
            .I(N__42304));
    LocalMux I__9295 (
            .O(N__42391),
            .I(N__42304));
    Span4Mux_h I__9294 (
            .O(N__42380),
            .I(N__42304));
    Odrv4 I__9293 (
            .O(N__42377),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__9292 (
            .O(N__42372),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9291 (
            .O(N__42359),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9290 (
            .O(N__42352),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9289 (
            .O(N__42335),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__9288 (
            .O(N__42328),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__9287 (
            .O(N__42315),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__9286 (
            .O(N__42304),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    CascadeMux I__9285 (
            .O(N__42287),
            .I(N__42282));
    InMux I__9284 (
            .O(N__42286),
            .I(N__42279));
    InMux I__9283 (
            .O(N__42285),
            .I(N__42276));
    InMux I__9282 (
            .O(N__42282),
            .I(N__42273));
    LocalMux I__9281 (
            .O(N__42279),
            .I(N__42270));
    LocalMux I__9280 (
            .O(N__42276),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__9279 (
            .O(N__42273),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv12 I__9278 (
            .O(N__42270),
            .I(\current_shift_inst.un4_control_input1_26 ));
    CascadeMux I__9277 (
            .O(N__42263),
            .I(N__42260));
    InMux I__9276 (
            .O(N__42260),
            .I(N__42257));
    LocalMux I__9275 (
            .O(N__42257),
            .I(N__42252));
    InMux I__9274 (
            .O(N__42256),
            .I(N__42249));
    InMux I__9273 (
            .O(N__42255),
            .I(N__42246));
    Span4Mux_h I__9272 (
            .O(N__42252),
            .I(N__42242));
    LocalMux I__9271 (
            .O(N__42249),
            .I(N__42239));
    LocalMux I__9270 (
            .O(N__42246),
            .I(N__42236));
    InMux I__9269 (
            .O(N__42245),
            .I(N__42233));
    Odrv4 I__9268 (
            .O(N__42242),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__9267 (
            .O(N__42239),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__9266 (
            .O(N__42236),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__9265 (
            .O(N__42233),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__9264 (
            .O(N__42224),
            .I(N__42221));
    LocalMux I__9263 (
            .O(N__42221),
            .I(N__42218));
    Span4Mux_h I__9262 (
            .O(N__42218),
            .I(N__42215));
    Span4Mux_h I__9261 (
            .O(N__42215),
            .I(N__42212));
    Odrv4 I__9260 (
            .O(N__42212),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    CascadeMux I__9259 (
            .O(N__42209),
            .I(N__42205));
    InMux I__9258 (
            .O(N__42208),
            .I(N__42202));
    InMux I__9257 (
            .O(N__42205),
            .I(N__42199));
    LocalMux I__9256 (
            .O(N__42202),
            .I(N__42195));
    LocalMux I__9255 (
            .O(N__42199),
            .I(N__42192));
    InMux I__9254 (
            .O(N__42198),
            .I(N__42189));
    Span4Mux_v I__9253 (
            .O(N__42195),
            .I(N__42185));
    Span4Mux_h I__9252 (
            .O(N__42192),
            .I(N__42180));
    LocalMux I__9251 (
            .O(N__42189),
            .I(N__42180));
    InMux I__9250 (
            .O(N__42188),
            .I(N__42177));
    Odrv4 I__9249 (
            .O(N__42185),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__9248 (
            .O(N__42180),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__9247 (
            .O(N__42177),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__9246 (
            .O(N__42170),
            .I(N__42166));
    CascadeMux I__9245 (
            .O(N__42169),
            .I(N__42163));
    LocalMux I__9244 (
            .O(N__42166),
            .I(N__42159));
    InMux I__9243 (
            .O(N__42163),
            .I(N__42156));
    InMux I__9242 (
            .O(N__42162),
            .I(N__42153));
    Odrv4 I__9241 (
            .O(N__42159),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__9240 (
            .O(N__42156),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__9239 (
            .O(N__42153),
            .I(\current_shift_inst.un4_control_input1_30 ));
    CascadeMux I__9238 (
            .O(N__42146),
            .I(N__42142));
    InMux I__9237 (
            .O(N__42145),
            .I(N__42139));
    InMux I__9236 (
            .O(N__42142),
            .I(N__42136));
    LocalMux I__9235 (
            .O(N__42139),
            .I(N__42133));
    LocalMux I__9234 (
            .O(N__42136),
            .I(N__42126));
    Span4Mux_v I__9233 (
            .O(N__42133),
            .I(N__42126));
    InMux I__9232 (
            .O(N__42132),
            .I(N__42123));
    InMux I__9231 (
            .O(N__42131),
            .I(N__42120));
    Odrv4 I__9230 (
            .O(N__42126),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__9229 (
            .O(N__42123),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__9228 (
            .O(N__42120),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__9227 (
            .O(N__42113),
            .I(N__42110));
    LocalMux I__9226 (
            .O(N__42110),
            .I(N__42105));
    InMux I__9225 (
            .O(N__42109),
            .I(N__42102));
    InMux I__9224 (
            .O(N__42108),
            .I(N__42099));
    Span4Mux_v I__9223 (
            .O(N__42105),
            .I(N__42094));
    LocalMux I__9222 (
            .O(N__42102),
            .I(N__42094));
    LocalMux I__9221 (
            .O(N__42099),
            .I(N__42091));
    Span4Mux_v I__9220 (
            .O(N__42094),
            .I(N__42086));
    Span4Mux_v I__9219 (
            .O(N__42091),
            .I(N__42086));
    Odrv4 I__9218 (
            .O(N__42086),
            .I(\current_shift_inst.un4_control_input1_3 ));
    CascadeMux I__9217 (
            .O(N__42083),
            .I(N__42080));
    InMux I__9216 (
            .O(N__42080),
            .I(N__42077));
    LocalMux I__9215 (
            .O(N__42077),
            .I(N__42072));
    InMux I__9214 (
            .O(N__42076),
            .I(N__42069));
    InMux I__9213 (
            .O(N__42075),
            .I(N__42066));
    Span4Mux_h I__9212 (
            .O(N__42072),
            .I(N__42060));
    LocalMux I__9211 (
            .O(N__42069),
            .I(N__42060));
    LocalMux I__9210 (
            .O(N__42066),
            .I(N__42057));
    InMux I__9209 (
            .O(N__42065),
            .I(N__42054));
    Odrv4 I__9208 (
            .O(N__42060),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__9207 (
            .O(N__42057),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__9206 (
            .O(N__42054),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__9205 (
            .O(N__42047),
            .I(N__42044));
    LocalMux I__9204 (
            .O(N__42044),
            .I(N__42041));
    Span4Mux_h I__9203 (
            .O(N__42041),
            .I(N__42038));
    Odrv4 I__9202 (
            .O(N__42038),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    CascadeMux I__9201 (
            .O(N__42035),
            .I(N__42031));
    CascadeMux I__9200 (
            .O(N__42034),
            .I(N__42028));
    InMux I__9199 (
            .O(N__42031),
            .I(N__42023));
    InMux I__9198 (
            .O(N__42028),
            .I(N__42023));
    LocalMux I__9197 (
            .O(N__42023),
            .I(N__42018));
    InMux I__9196 (
            .O(N__42022),
            .I(N__42015));
    InMux I__9195 (
            .O(N__42021),
            .I(N__42012));
    Span4Mux_h I__9194 (
            .O(N__42018),
            .I(N__42007));
    LocalMux I__9193 (
            .O(N__42015),
            .I(N__42007));
    LocalMux I__9192 (
            .O(N__42012),
            .I(N__42004));
    Odrv4 I__9191 (
            .O(N__42007),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv12 I__9190 (
            .O(N__42004),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__9189 (
            .O(N__41999),
            .I(N__41993));
    InMux I__9188 (
            .O(N__41998),
            .I(N__41993));
    LocalMux I__9187 (
            .O(N__41993),
            .I(N__41989));
    InMux I__9186 (
            .O(N__41992),
            .I(N__41986));
    Span4Mux_h I__9185 (
            .O(N__41989),
            .I(N__41981));
    LocalMux I__9184 (
            .O(N__41986),
            .I(N__41981));
    Span4Mux_v I__9183 (
            .O(N__41981),
            .I(N__41978));
    Odrv4 I__9182 (
            .O(N__41978),
            .I(\current_shift_inst.un4_control_input1_4 ));
    CascadeMux I__9181 (
            .O(N__41975),
            .I(N__41971));
    CascadeMux I__9180 (
            .O(N__41974),
            .I(N__41968));
    InMux I__9179 (
            .O(N__41971),
            .I(N__41965));
    InMux I__9178 (
            .O(N__41968),
            .I(N__41962));
    LocalMux I__9177 (
            .O(N__41965),
            .I(N__41959));
    LocalMux I__9176 (
            .O(N__41962),
            .I(N__41955));
    Sp12to4 I__9175 (
            .O(N__41959),
            .I(N__41952));
    InMux I__9174 (
            .O(N__41958),
            .I(N__41949));
    Span4Mux_v I__9173 (
            .O(N__41955),
            .I(N__41945));
    Span12Mux_v I__9172 (
            .O(N__41952),
            .I(N__41942));
    LocalMux I__9171 (
            .O(N__41949),
            .I(N__41939));
    InMux I__9170 (
            .O(N__41948),
            .I(N__41936));
    Odrv4 I__9169 (
            .O(N__41945),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv12 I__9168 (
            .O(N__41942),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__9167 (
            .O(N__41939),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__9166 (
            .O(N__41936),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__9165 (
            .O(N__41927),
            .I(N__41923));
    InMux I__9164 (
            .O(N__41926),
            .I(N__41920));
    LocalMux I__9163 (
            .O(N__41923),
            .I(N__41917));
    LocalMux I__9162 (
            .O(N__41920),
            .I(N__41911));
    Span4Mux_v I__9161 (
            .O(N__41917),
            .I(N__41911));
    InMux I__9160 (
            .O(N__41916),
            .I(N__41908));
    Odrv4 I__9159 (
            .O(N__41911),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__9158 (
            .O(N__41908),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__9157 (
            .O(N__41903),
            .I(N__41900));
    LocalMux I__9156 (
            .O(N__41900),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__9155 (
            .O(N__41897),
            .I(N__41892));
    InMux I__9154 (
            .O(N__41896),
            .I(N__41889));
    InMux I__9153 (
            .O(N__41895),
            .I(N__41886));
    LocalMux I__9152 (
            .O(N__41892),
            .I(N__41880));
    LocalMux I__9151 (
            .O(N__41889),
            .I(N__41880));
    LocalMux I__9150 (
            .O(N__41886),
            .I(N__41877));
    InMux I__9149 (
            .O(N__41885),
            .I(N__41874));
    Span4Mux_h I__9148 (
            .O(N__41880),
            .I(N__41867));
    Span4Mux_v I__9147 (
            .O(N__41877),
            .I(N__41867));
    LocalMux I__9146 (
            .O(N__41874),
            .I(N__41867));
    Odrv4 I__9145 (
            .O(N__41867),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__9144 (
            .O(N__41864),
            .I(N__41861));
    LocalMux I__9143 (
            .O(N__41861),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    CascadeMux I__9142 (
            .O(N__41858),
            .I(N__41853));
    InMux I__9141 (
            .O(N__41857),
            .I(N__41850));
    InMux I__9140 (
            .O(N__41856),
            .I(N__41847));
    InMux I__9139 (
            .O(N__41853),
            .I(N__41844));
    LocalMux I__9138 (
            .O(N__41850),
            .I(N__41840));
    LocalMux I__9137 (
            .O(N__41847),
            .I(N__41837));
    LocalMux I__9136 (
            .O(N__41844),
            .I(N__41834));
    InMux I__9135 (
            .O(N__41843),
            .I(N__41831));
    Span4Mux_h I__9134 (
            .O(N__41840),
            .I(N__41828));
    Span4Mux_h I__9133 (
            .O(N__41837),
            .I(N__41825));
    Span4Mux_v I__9132 (
            .O(N__41834),
            .I(N__41820));
    LocalMux I__9131 (
            .O(N__41831),
            .I(N__41820));
    Odrv4 I__9130 (
            .O(N__41828),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__9129 (
            .O(N__41825),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__9128 (
            .O(N__41820),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__9127 (
            .O(N__41813),
            .I(N__41810));
    LocalMux I__9126 (
            .O(N__41810),
            .I(N__41805));
    InMux I__9125 (
            .O(N__41809),
            .I(N__41802));
    InMux I__9124 (
            .O(N__41808),
            .I(N__41799));
    Odrv4 I__9123 (
            .O(N__41805),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__9122 (
            .O(N__41802),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__9121 (
            .O(N__41799),
            .I(\current_shift_inst.un4_control_input1_20 ));
    CascadeMux I__9120 (
            .O(N__41792),
            .I(N__41788));
    InMux I__9119 (
            .O(N__41791),
            .I(N__41785));
    InMux I__9118 (
            .O(N__41788),
            .I(N__41782));
    LocalMux I__9117 (
            .O(N__41785),
            .I(N__41778));
    LocalMux I__9116 (
            .O(N__41782),
            .I(N__41775));
    InMux I__9115 (
            .O(N__41781),
            .I(N__41772));
    Span4Mux_v I__9114 (
            .O(N__41778),
            .I(N__41766));
    Span4Mux_h I__9113 (
            .O(N__41775),
            .I(N__41766));
    LocalMux I__9112 (
            .O(N__41772),
            .I(N__41763));
    InMux I__9111 (
            .O(N__41771),
            .I(N__41760));
    Odrv4 I__9110 (
            .O(N__41766),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__9109 (
            .O(N__41763),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__9108 (
            .O(N__41760),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__9107 (
            .O(N__41753),
            .I(N__41749));
    CascadeMux I__9106 (
            .O(N__41752),
            .I(N__41746));
    LocalMux I__9105 (
            .O(N__41749),
            .I(N__41743));
    InMux I__9104 (
            .O(N__41746),
            .I(N__41739));
    Span4Mux_h I__9103 (
            .O(N__41743),
            .I(N__41736));
    InMux I__9102 (
            .O(N__41742),
            .I(N__41733));
    LocalMux I__9101 (
            .O(N__41739),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv4 I__9100 (
            .O(N__41736),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__9099 (
            .O(N__41733),
            .I(\current_shift_inst.un4_control_input1_19 ));
    CascadeMux I__9098 (
            .O(N__41726),
            .I(N__41722));
    InMux I__9097 (
            .O(N__41725),
            .I(N__41716));
    InMux I__9096 (
            .O(N__41722),
            .I(N__41716));
    InMux I__9095 (
            .O(N__41721),
            .I(N__41713));
    LocalMux I__9094 (
            .O(N__41716),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__9093 (
            .O(N__41713),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__9092 (
            .O(N__41708),
            .I(N__41700));
    InMux I__9091 (
            .O(N__41707),
            .I(N__41700));
    InMux I__9090 (
            .O(N__41706),
            .I(N__41695));
    InMux I__9089 (
            .O(N__41705),
            .I(N__41695));
    LocalMux I__9088 (
            .O(N__41700),
            .I(N__41692));
    LocalMux I__9087 (
            .O(N__41695),
            .I(N__41689));
    Odrv4 I__9086 (
            .O(N__41692),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__9085 (
            .O(N__41689),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    CascadeMux I__9084 (
            .O(N__41684),
            .I(N__41681));
    InMux I__9083 (
            .O(N__41681),
            .I(N__41678));
    LocalMux I__9082 (
            .O(N__41678),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__9081 (
            .O(N__41675),
            .I(N__41672));
    LocalMux I__9080 (
            .O(N__41672),
            .I(N__41667));
    InMux I__9079 (
            .O(N__41671),
            .I(N__41664));
    InMux I__9078 (
            .O(N__41670),
            .I(N__41661));
    Span4Mux_v I__9077 (
            .O(N__41667),
            .I(N__41657));
    LocalMux I__9076 (
            .O(N__41664),
            .I(N__41654));
    LocalMux I__9075 (
            .O(N__41661),
            .I(N__41651));
    InMux I__9074 (
            .O(N__41660),
            .I(N__41648));
    Odrv4 I__9073 (
            .O(N__41657),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv4 I__9072 (
            .O(N__41654),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv4 I__9071 (
            .O(N__41651),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__9070 (
            .O(N__41648),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    CascadeMux I__9069 (
            .O(N__41639),
            .I(N__41635));
    InMux I__9068 (
            .O(N__41638),
            .I(N__41632));
    InMux I__9067 (
            .O(N__41635),
            .I(N__41628));
    LocalMux I__9066 (
            .O(N__41632),
            .I(N__41625));
    InMux I__9065 (
            .O(N__41631),
            .I(N__41622));
    LocalMux I__9064 (
            .O(N__41628),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv4 I__9063 (
            .O(N__41625),
            .I(\current_shift_inst.un4_control_input1_22 ));
    LocalMux I__9062 (
            .O(N__41622),
            .I(\current_shift_inst.un4_control_input1_22 ));
    CascadeMux I__9061 (
            .O(N__41615),
            .I(N__41611));
    CascadeMux I__9060 (
            .O(N__41614),
            .I(N__41608));
    InMux I__9059 (
            .O(N__41611),
            .I(N__41604));
    InMux I__9058 (
            .O(N__41608),
            .I(N__41599));
    InMux I__9057 (
            .O(N__41607),
            .I(N__41599));
    LocalMux I__9056 (
            .O(N__41604),
            .I(N__41595));
    LocalMux I__9055 (
            .O(N__41599),
            .I(N__41592));
    InMux I__9054 (
            .O(N__41598),
            .I(N__41589));
    Span4Mux_v I__9053 (
            .O(N__41595),
            .I(N__41586));
    Span4Mux_h I__9052 (
            .O(N__41592),
            .I(N__41583));
    LocalMux I__9051 (
            .O(N__41589),
            .I(N__41580));
    Odrv4 I__9050 (
            .O(N__41586),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__9049 (
            .O(N__41583),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv12 I__9048 (
            .O(N__41580),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__9047 (
            .O(N__41573),
            .I(N__41570));
    LocalMux I__9046 (
            .O(N__41570),
            .I(N__41567));
    Span4Mux_h I__9045 (
            .O(N__41567),
            .I(N__41562));
    InMux I__9044 (
            .O(N__41566),
            .I(N__41557));
    InMux I__9043 (
            .O(N__41565),
            .I(N__41557));
    Odrv4 I__9042 (
            .O(N__41562),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__9041 (
            .O(N__41557),
            .I(\current_shift_inst.un4_control_input1_9 ));
    CascadeMux I__9040 (
            .O(N__41552),
            .I(N__41549));
    InMux I__9039 (
            .O(N__41549),
            .I(N__41546));
    LocalMux I__9038 (
            .O(N__41546),
            .I(N__41543));
    Span4Mux_h I__9037 (
            .O(N__41543),
            .I(N__41540));
    Odrv4 I__9036 (
            .O(N__41540),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    InMux I__9035 (
            .O(N__41537),
            .I(N__41532));
    InMux I__9034 (
            .O(N__41536),
            .I(N__41529));
    InMux I__9033 (
            .O(N__41535),
            .I(N__41526));
    LocalMux I__9032 (
            .O(N__41532),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__9031 (
            .O(N__41529),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__9030 (
            .O(N__41526),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__9029 (
            .O(N__41519),
            .I(N__41514));
    InMux I__9028 (
            .O(N__41518),
            .I(N__41508));
    InMux I__9027 (
            .O(N__41517),
            .I(N__41508));
    LocalMux I__9026 (
            .O(N__41514),
            .I(N__41505));
    InMux I__9025 (
            .O(N__41513),
            .I(N__41502));
    LocalMux I__9024 (
            .O(N__41508),
            .I(N__41499));
    Span4Mux_h I__9023 (
            .O(N__41505),
            .I(N__41496));
    LocalMux I__9022 (
            .O(N__41502),
            .I(N__41493));
    Span4Mux_v I__9021 (
            .O(N__41499),
            .I(N__41490));
    Odrv4 I__9020 (
            .O(N__41496),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__9019 (
            .O(N__41493),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__9018 (
            .O(N__41490),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__9017 (
            .O(N__41483),
            .I(N__41480));
    LocalMux I__9016 (
            .O(N__41480),
            .I(N__41476));
    InMux I__9015 (
            .O(N__41479),
            .I(N__41473));
    Span4Mux_h I__9014 (
            .O(N__41476),
            .I(N__41469));
    LocalMux I__9013 (
            .O(N__41473),
            .I(N__41466));
    InMux I__9012 (
            .O(N__41472),
            .I(N__41463));
    Odrv4 I__9011 (
            .O(N__41469),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__9010 (
            .O(N__41466),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__9009 (
            .O(N__41463),
            .I(\current_shift_inst.un4_control_input1_5 ));
    CascadeMux I__9008 (
            .O(N__41456),
            .I(N__41453));
    InMux I__9007 (
            .O(N__41453),
            .I(N__41450));
    LocalMux I__9006 (
            .O(N__41450),
            .I(N__41447));
    Span4Mux_h I__9005 (
            .O(N__41447),
            .I(N__41444));
    Odrv4 I__9004 (
            .O(N__41444),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ));
    CascadeMux I__9003 (
            .O(N__41441),
            .I(N__41437));
    CascadeMux I__9002 (
            .O(N__41440),
            .I(N__41434));
    InMux I__9001 (
            .O(N__41437),
            .I(N__41431));
    InMux I__9000 (
            .O(N__41434),
            .I(N__41428));
    LocalMux I__8999 (
            .O(N__41431),
            .I(N__41422));
    LocalMux I__8998 (
            .O(N__41428),
            .I(N__41422));
    InMux I__8997 (
            .O(N__41427),
            .I(N__41419));
    Span4Mux_h I__8996 (
            .O(N__41422),
            .I(N__41413));
    LocalMux I__8995 (
            .O(N__41419),
            .I(N__41413));
    InMux I__8994 (
            .O(N__41418),
            .I(N__41410));
    Odrv4 I__8993 (
            .O(N__41413),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__8992 (
            .O(N__41410),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__8991 (
            .O(N__41405),
            .I(N__41402));
    LocalMux I__8990 (
            .O(N__41402),
            .I(N__41398));
    InMux I__8989 (
            .O(N__41401),
            .I(N__41394));
    Span4Mux_h I__8988 (
            .O(N__41398),
            .I(N__41391));
    InMux I__8987 (
            .O(N__41397),
            .I(N__41388));
    LocalMux I__8986 (
            .O(N__41394),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__8985 (
            .O(N__41391),
            .I(\current_shift_inst.un4_control_input1_16 ));
    LocalMux I__8984 (
            .O(N__41388),
            .I(\current_shift_inst.un4_control_input1_16 ));
    CascadeMux I__8983 (
            .O(N__41381),
            .I(N__41378));
    InMux I__8982 (
            .O(N__41378),
            .I(N__41373));
    InMux I__8981 (
            .O(N__41377),
            .I(N__41370));
    InMux I__8980 (
            .O(N__41376),
            .I(N__41366));
    LocalMux I__8979 (
            .O(N__41373),
            .I(N__41361));
    LocalMux I__8978 (
            .O(N__41370),
            .I(N__41361));
    InMux I__8977 (
            .O(N__41369),
            .I(N__41358));
    LocalMux I__8976 (
            .O(N__41366),
            .I(N__41355));
    Span4Mux_h I__8975 (
            .O(N__41361),
            .I(N__41350));
    LocalMux I__8974 (
            .O(N__41358),
            .I(N__41350));
    Odrv4 I__8973 (
            .O(N__41355),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__8972 (
            .O(N__41350),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__8971 (
            .O(N__41345),
            .I(N__41341));
    InMux I__8970 (
            .O(N__41344),
            .I(N__41338));
    LocalMux I__8969 (
            .O(N__41341),
            .I(N__41334));
    LocalMux I__8968 (
            .O(N__41338),
            .I(N__41331));
    InMux I__8967 (
            .O(N__41337),
            .I(N__41328));
    Odrv4 I__8966 (
            .O(N__41334),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv12 I__8965 (
            .O(N__41331),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__8964 (
            .O(N__41328),
            .I(\current_shift_inst.un4_control_input1_13 ));
    CascadeMux I__8963 (
            .O(N__41321),
            .I(N__41318));
    InMux I__8962 (
            .O(N__41318),
            .I(N__41315));
    LocalMux I__8961 (
            .O(N__41315),
            .I(N__41312));
    Span4Mux_h I__8960 (
            .O(N__41312),
            .I(N__41309));
    Span4Mux_h I__8959 (
            .O(N__41309),
            .I(N__41306));
    Odrv4 I__8958 (
            .O(N__41306),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    InMux I__8957 (
            .O(N__41303),
            .I(N__41298));
    InMux I__8956 (
            .O(N__41302),
            .I(N__41295));
    InMux I__8955 (
            .O(N__41301),
            .I(N__41292));
    LocalMux I__8954 (
            .O(N__41298),
            .I(N__41289));
    LocalMux I__8953 (
            .O(N__41295),
            .I(N__41286));
    LocalMux I__8952 (
            .O(N__41292),
            .I(N__41283));
    Span4Mux_v I__8951 (
            .O(N__41289),
            .I(N__41280));
    Span4Mux_h I__8950 (
            .O(N__41286),
            .I(N__41275));
    Span4Mux_v I__8949 (
            .O(N__41283),
            .I(N__41275));
    Span4Mux_h I__8948 (
            .O(N__41280),
            .I(N__41269));
    Span4Mux_v I__8947 (
            .O(N__41275),
            .I(N__41269));
    InMux I__8946 (
            .O(N__41274),
            .I(N__41266));
    Sp12to4 I__8945 (
            .O(N__41269),
            .I(N__41263));
    LocalMux I__8944 (
            .O(N__41266),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv12 I__8943 (
            .O(N__41263),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__8942 (
            .O(N__41258),
            .I(N__41255));
    LocalMux I__8941 (
            .O(N__41255),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__8940 (
            .O(N__41252),
            .I(N__41247));
    CascadeMux I__8939 (
            .O(N__41251),
            .I(N__41244));
    InMux I__8938 (
            .O(N__41250),
            .I(N__41241));
    LocalMux I__8937 (
            .O(N__41247),
            .I(N__41238));
    InMux I__8936 (
            .O(N__41244),
            .I(N__41235));
    LocalMux I__8935 (
            .O(N__41241),
            .I(N__41232));
    Span4Mux_v I__8934 (
            .O(N__41238),
            .I(N__41228));
    LocalMux I__8933 (
            .O(N__41235),
            .I(N__41225));
    Span4Mux_h I__8932 (
            .O(N__41232),
            .I(N__41222));
    InMux I__8931 (
            .O(N__41231),
            .I(N__41219));
    Odrv4 I__8930 (
            .O(N__41228),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__8929 (
            .O(N__41225),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__8928 (
            .O(N__41222),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__8927 (
            .O(N__41219),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__8926 (
            .O(N__41210),
            .I(N__41206));
    InMux I__8925 (
            .O(N__41209),
            .I(N__41203));
    LocalMux I__8924 (
            .O(N__41206),
            .I(N__41200));
    LocalMux I__8923 (
            .O(N__41203),
            .I(N__41196));
    Span4Mux_h I__8922 (
            .O(N__41200),
            .I(N__41193));
    InMux I__8921 (
            .O(N__41199),
            .I(N__41190));
    Odrv12 I__8920 (
            .O(N__41196),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__8919 (
            .O(N__41193),
            .I(\current_shift_inst.un4_control_input1_17 ));
    LocalMux I__8918 (
            .O(N__41190),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CascadeMux I__8917 (
            .O(N__41183),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    CascadeMux I__8916 (
            .O(N__41180),
            .I(N__41176));
    InMux I__8915 (
            .O(N__41179),
            .I(N__41173));
    InMux I__8914 (
            .O(N__41176),
            .I(N__41170));
    LocalMux I__8913 (
            .O(N__41173),
            .I(N__41167));
    LocalMux I__8912 (
            .O(N__41170),
            .I(N__41164));
    Span4Mux_h I__8911 (
            .O(N__41167),
            .I(N__41159));
    Span4Mux_v I__8910 (
            .O(N__41164),
            .I(N__41159));
    Odrv4 I__8909 (
            .O(N__41159),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    CascadeMux I__8908 (
            .O(N__41156),
            .I(N__41153));
    InMux I__8907 (
            .O(N__41153),
            .I(N__41150));
    LocalMux I__8906 (
            .O(N__41150),
            .I(N__41147));
    Span4Mux_h I__8905 (
            .O(N__41147),
            .I(N__41144));
    Odrv4 I__8904 (
            .O(N__41144),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ));
    InMux I__8903 (
            .O(N__41141),
            .I(N__41138));
    LocalMux I__8902 (
            .O(N__41138),
            .I(N__41135));
    Span4Mux_h I__8901 (
            .O(N__41135),
            .I(N__41129));
    InMux I__8900 (
            .O(N__41134),
            .I(N__41126));
    InMux I__8899 (
            .O(N__41133),
            .I(N__41121));
    InMux I__8898 (
            .O(N__41132),
            .I(N__41121));
    Span4Mux_h I__8897 (
            .O(N__41129),
            .I(N__41116));
    LocalMux I__8896 (
            .O(N__41126),
            .I(N__41116));
    LocalMux I__8895 (
            .O(N__41121),
            .I(N__41113));
    Odrv4 I__8894 (
            .O(N__41116),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv12 I__8893 (
            .O(N__41113),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__8892 (
            .O(N__41108),
            .I(N__41105));
    LocalMux I__8891 (
            .O(N__41105),
            .I(N__41100));
    InMux I__8890 (
            .O(N__41104),
            .I(N__41097));
    InMux I__8889 (
            .O(N__41103),
            .I(N__41094));
    Odrv4 I__8888 (
            .O(N__41100),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__8887 (
            .O(N__41097),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__8886 (
            .O(N__41094),
            .I(\current_shift_inst.un4_control_input1_6 ));
    CascadeMux I__8885 (
            .O(N__41087),
            .I(N__41084));
    InMux I__8884 (
            .O(N__41084),
            .I(N__41081));
    LocalMux I__8883 (
            .O(N__41081),
            .I(N__41076));
    InMux I__8882 (
            .O(N__41080),
            .I(N__41073));
    InMux I__8881 (
            .O(N__41079),
            .I(N__41070));
    Span4Mux_h I__8880 (
            .O(N__41076),
            .I(N__41065));
    LocalMux I__8879 (
            .O(N__41073),
            .I(N__41065));
    LocalMux I__8878 (
            .O(N__41070),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__8877 (
            .O(N__41065),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__8876 (
            .O(N__41060),
            .I(N__41056));
    CascadeMux I__8875 (
            .O(N__41059),
            .I(N__41052));
    LocalMux I__8874 (
            .O(N__41056),
            .I(N__41049));
    InMux I__8873 (
            .O(N__41055),
            .I(N__41045));
    InMux I__8872 (
            .O(N__41052),
            .I(N__41042));
    Span4Mux_h I__8871 (
            .O(N__41049),
            .I(N__41039));
    InMux I__8870 (
            .O(N__41048),
            .I(N__41036));
    LocalMux I__8869 (
            .O(N__41045),
            .I(N__41033));
    LocalMux I__8868 (
            .O(N__41042),
            .I(N__41030));
    Span4Mux_v I__8867 (
            .O(N__41039),
            .I(N__41025));
    LocalMux I__8866 (
            .O(N__41036),
            .I(N__41025));
    Odrv12 I__8865 (
            .O(N__41033),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__8864 (
            .O(N__41030),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__8863 (
            .O(N__41025),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    CascadeMux I__8862 (
            .O(N__41018),
            .I(N__41014));
    InMux I__8861 (
            .O(N__41017),
            .I(N__41011));
    InMux I__8860 (
            .O(N__41014),
            .I(N__41008));
    LocalMux I__8859 (
            .O(N__41011),
            .I(N__41005));
    LocalMux I__8858 (
            .O(N__41008),
            .I(N__41002));
    Span4Mux_h I__8857 (
            .O(N__41005),
            .I(N__40999));
    Span4Mux_h I__8856 (
            .O(N__41002),
            .I(N__40993));
    Span4Mux_v I__8855 (
            .O(N__40999),
            .I(N__40993));
    InMux I__8854 (
            .O(N__40998),
            .I(N__40990));
    Odrv4 I__8853 (
            .O(N__40993),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__8852 (
            .O(N__40990),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__8851 (
            .O(N__40985),
            .I(N__40980));
    InMux I__8850 (
            .O(N__40984),
            .I(N__40977));
    InMux I__8849 (
            .O(N__40983),
            .I(N__40974));
    LocalMux I__8848 (
            .O(N__40980),
            .I(N__40971));
    LocalMux I__8847 (
            .O(N__40977),
            .I(N__40968));
    LocalMux I__8846 (
            .O(N__40974),
            .I(N__40965));
    Span4Mux_v I__8845 (
            .O(N__40971),
            .I(N__40957));
    Span4Mux_h I__8844 (
            .O(N__40968),
            .I(N__40957));
    Span4Mux_h I__8843 (
            .O(N__40965),
            .I(N__40957));
    InMux I__8842 (
            .O(N__40964),
            .I(N__40954));
    Odrv4 I__8841 (
            .O(N__40957),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__8840 (
            .O(N__40954),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    CascadeMux I__8839 (
            .O(N__40949),
            .I(N__40945));
    InMux I__8838 (
            .O(N__40948),
            .I(N__40942));
    InMux I__8837 (
            .O(N__40945),
            .I(N__40939));
    LocalMux I__8836 (
            .O(N__40942),
            .I(N__40936));
    LocalMux I__8835 (
            .O(N__40939),
            .I(N__40933));
    Span4Mux_h I__8834 (
            .O(N__40936),
            .I(N__40929));
    Span4Mux_h I__8833 (
            .O(N__40933),
            .I(N__40926));
    InMux I__8832 (
            .O(N__40932),
            .I(N__40923));
    Odrv4 I__8831 (
            .O(N__40929),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__8830 (
            .O(N__40926),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__8829 (
            .O(N__40923),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__8828 (
            .O(N__40916),
            .I(N__40913));
    LocalMux I__8827 (
            .O(N__40913),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__8826 (
            .O(N__40910),
            .I(N__40906));
    CascadeMux I__8825 (
            .O(N__40909),
            .I(N__40903));
    InMux I__8824 (
            .O(N__40906),
            .I(N__40900));
    InMux I__8823 (
            .O(N__40903),
            .I(N__40896));
    LocalMux I__8822 (
            .O(N__40900),
            .I(N__40893));
    InMux I__8821 (
            .O(N__40899),
            .I(N__40890));
    LocalMux I__8820 (
            .O(N__40896),
            .I(N__40887));
    Span4Mux_v I__8819 (
            .O(N__40893),
            .I(N__40883));
    LocalMux I__8818 (
            .O(N__40890),
            .I(N__40880));
    Span4Mux_v I__8817 (
            .O(N__40887),
            .I(N__40877));
    InMux I__8816 (
            .O(N__40886),
            .I(N__40874));
    Span4Mux_h I__8815 (
            .O(N__40883),
            .I(N__40869));
    Span4Mux_v I__8814 (
            .O(N__40880),
            .I(N__40869));
    Odrv4 I__8813 (
            .O(N__40877),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__8812 (
            .O(N__40874),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__8811 (
            .O(N__40869),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__8810 (
            .O(N__40862),
            .I(N__40859));
    InMux I__8809 (
            .O(N__40859),
            .I(N__40856));
    LocalMux I__8808 (
            .O(N__40856),
            .I(N__40853));
    Span4Mux_v I__8807 (
            .O(N__40853),
            .I(N__40850));
    Odrv4 I__8806 (
            .O(N__40850),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    InMux I__8805 (
            .O(N__40847),
            .I(N__40844));
    LocalMux I__8804 (
            .O(N__40844),
            .I(N__40841));
    Span4Mux_h I__8803 (
            .O(N__40841),
            .I(N__40838));
    Span4Mux_v I__8802 (
            .O(N__40838),
            .I(N__40832));
    InMux I__8801 (
            .O(N__40837),
            .I(N__40829));
    InMux I__8800 (
            .O(N__40836),
            .I(N__40824));
    InMux I__8799 (
            .O(N__40835),
            .I(N__40824));
    Odrv4 I__8798 (
            .O(N__40832),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__8797 (
            .O(N__40829),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__8796 (
            .O(N__40824),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    InMux I__8795 (
            .O(N__40817),
            .I(N__40814));
    LocalMux I__8794 (
            .O(N__40814),
            .I(N__40811));
    Span4Mux_v I__8793 (
            .O(N__40811),
            .I(N__40806));
    InMux I__8792 (
            .O(N__40810),
            .I(N__40803));
    InMux I__8791 (
            .O(N__40809),
            .I(N__40800));
    Odrv4 I__8790 (
            .O(N__40806),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__8789 (
            .O(N__40803),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__8788 (
            .O(N__40800),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__8787 (
            .O(N__40793),
            .I(N__40790));
    LocalMux I__8786 (
            .O(N__40790),
            .I(N__40787));
    Span4Mux_h I__8785 (
            .O(N__40787),
            .I(N__40784));
    Span4Mux_h I__8784 (
            .O(N__40784),
            .I(N__40781));
    Odrv4 I__8783 (
            .O(N__40781),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ));
    InMux I__8782 (
            .O(N__40778),
            .I(N__40775));
    LocalMux I__8781 (
            .O(N__40775),
            .I(N__40772));
    Span4Mux_h I__8780 (
            .O(N__40772),
            .I(N__40769));
    Odrv4 I__8779 (
            .O(N__40769),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ));
    InMux I__8778 (
            .O(N__40766),
            .I(N__40763));
    LocalMux I__8777 (
            .O(N__40763),
            .I(N__40760));
    Span4Mux_h I__8776 (
            .O(N__40760),
            .I(N__40757));
    Span4Mux_v I__8775 (
            .O(N__40757),
            .I(N__40754));
    Odrv4 I__8774 (
            .O(N__40754),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    CascadeMux I__8773 (
            .O(N__40751),
            .I(N__40747));
    InMux I__8772 (
            .O(N__40750),
            .I(N__40739));
    InMux I__8771 (
            .O(N__40747),
            .I(N__40739));
    InMux I__8770 (
            .O(N__40746),
            .I(N__40739));
    LocalMux I__8769 (
            .O(N__40739),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__8768 (
            .O(N__40736),
            .I(N__40733));
    LocalMux I__8767 (
            .O(N__40733),
            .I(N__40730));
    Odrv4 I__8766 (
            .O(N__40730),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    CascadeMux I__8765 (
            .O(N__40727),
            .I(N__40724));
    InMux I__8764 (
            .O(N__40724),
            .I(N__40721));
    LocalMux I__8763 (
            .O(N__40721),
            .I(N__40718));
    Odrv12 I__8762 (
            .O(N__40718),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    InMux I__8761 (
            .O(N__40715),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    InMux I__8760 (
            .O(N__40712),
            .I(N__40709));
    LocalMux I__8759 (
            .O(N__40709),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt24 ));
    CascadeMux I__8758 (
            .O(N__40706),
            .I(N__40703));
    InMux I__8757 (
            .O(N__40703),
            .I(N__40700));
    LocalMux I__8756 (
            .O(N__40700),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ));
    InMux I__8755 (
            .O(N__40697),
            .I(N__40694));
    LocalMux I__8754 (
            .O(N__40694),
            .I(N__40691));
    Span4Mux_h I__8753 (
            .O(N__40691),
            .I(N__40687));
    InMux I__8752 (
            .O(N__40690),
            .I(N__40684));
    Odrv4 I__8751 (
            .O(N__40687),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    LocalMux I__8750 (
            .O(N__40684),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    CascadeMux I__8749 (
            .O(N__40679),
            .I(N__40675));
    InMux I__8748 (
            .O(N__40678),
            .I(N__40672));
    InMux I__8747 (
            .O(N__40675),
            .I(N__40667));
    LocalMux I__8746 (
            .O(N__40672),
            .I(N__40664));
    InMux I__8745 (
            .O(N__40671),
            .I(N__40659));
    InMux I__8744 (
            .O(N__40670),
            .I(N__40659));
    LocalMux I__8743 (
            .O(N__40667),
            .I(N__40656));
    Span4Mux_h I__8742 (
            .O(N__40664),
            .I(N__40651));
    LocalMux I__8741 (
            .O(N__40659),
            .I(N__40651));
    Span4Mux_h I__8740 (
            .O(N__40656),
            .I(N__40648));
    Odrv4 I__8739 (
            .O(N__40651),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv4 I__8738 (
            .O(N__40648),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    CascadeMux I__8737 (
            .O(N__40643),
            .I(elapsed_time_ns_1_RNI36DN9_0_25_cascade_));
    CascadeMux I__8736 (
            .O(N__40640),
            .I(N__40636));
    InMux I__8735 (
            .O(N__40639),
            .I(N__40631));
    InMux I__8734 (
            .O(N__40636),
            .I(N__40631));
    LocalMux I__8733 (
            .O(N__40631),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    InMux I__8732 (
            .O(N__40628),
            .I(N__40623));
    CascadeMux I__8731 (
            .O(N__40627),
            .I(N__40619));
    InMux I__8730 (
            .O(N__40626),
            .I(N__40616));
    LocalMux I__8729 (
            .O(N__40623),
            .I(N__40613));
    InMux I__8728 (
            .O(N__40622),
            .I(N__40610));
    InMux I__8727 (
            .O(N__40619),
            .I(N__40607));
    LocalMux I__8726 (
            .O(N__40616),
            .I(N__40604));
    Span4Mux_h I__8725 (
            .O(N__40613),
            .I(N__40601));
    LocalMux I__8724 (
            .O(N__40610),
            .I(N__40598));
    LocalMux I__8723 (
            .O(N__40607),
            .I(N__40595));
    Odrv4 I__8722 (
            .O(N__40604),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    Odrv4 I__8721 (
            .O(N__40601),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    Odrv4 I__8720 (
            .O(N__40598),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    Odrv4 I__8719 (
            .O(N__40595),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__8718 (
            .O(N__40586),
            .I(N__40583));
    LocalMux I__8717 (
            .O(N__40583),
            .I(N__40579));
    InMux I__8716 (
            .O(N__40582),
            .I(N__40575));
    Span4Mux_v I__8715 (
            .O(N__40579),
            .I(N__40572));
    InMux I__8714 (
            .O(N__40578),
            .I(N__40569));
    LocalMux I__8713 (
            .O(N__40575),
            .I(N__40566));
    Span4Mux_h I__8712 (
            .O(N__40572),
            .I(N__40563));
    LocalMux I__8711 (
            .O(N__40569),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    Odrv12 I__8710 (
            .O(N__40566),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    Odrv4 I__8709 (
            .O(N__40563),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    InMux I__8708 (
            .O(N__40556),
            .I(N__40550));
    InMux I__8707 (
            .O(N__40555),
            .I(N__40550));
    LocalMux I__8706 (
            .O(N__40550),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    CascadeMux I__8705 (
            .O(N__40547),
            .I(N__40544));
    InMux I__8704 (
            .O(N__40544),
            .I(N__40541));
    LocalMux I__8703 (
            .O(N__40541),
            .I(N__40538));
    Span4Mux_h I__8702 (
            .O(N__40538),
            .I(N__40535));
    Odrv4 I__8701 (
            .O(N__40535),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__8700 (
            .O(N__40532),
            .I(N__40529));
    LocalMux I__8699 (
            .O(N__40529),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__8698 (
            .O(N__40526),
            .I(N__40523));
    InMux I__8697 (
            .O(N__40523),
            .I(N__40520));
    LocalMux I__8696 (
            .O(N__40520),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__8695 (
            .O(N__40517),
            .I(N__40514));
    InMux I__8694 (
            .O(N__40514),
            .I(N__40511));
    LocalMux I__8693 (
            .O(N__40511),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__8692 (
            .O(N__40508),
            .I(N__40505));
    InMux I__8691 (
            .O(N__40505),
            .I(N__40502));
    LocalMux I__8690 (
            .O(N__40502),
            .I(N__40499));
    Odrv4 I__8689 (
            .O(N__40499),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__8688 (
            .O(N__40496),
            .I(N__40493));
    LocalMux I__8687 (
            .O(N__40493),
            .I(N__40490));
    Span4Mux_v I__8686 (
            .O(N__40490),
            .I(N__40487));
    Odrv4 I__8685 (
            .O(N__40487),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__8684 (
            .O(N__40484),
            .I(N__40481));
    InMux I__8683 (
            .O(N__40481),
            .I(N__40478));
    LocalMux I__8682 (
            .O(N__40478),
            .I(N__40475));
    Odrv4 I__8681 (
            .O(N__40475),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__8680 (
            .O(N__40472),
            .I(N__40469));
    InMux I__8679 (
            .O(N__40469),
            .I(N__40466));
    LocalMux I__8678 (
            .O(N__40466),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__8677 (
            .O(N__40463),
            .I(N__40460));
    LocalMux I__8676 (
            .O(N__40460),
            .I(N__40457));
    Span4Mux_h I__8675 (
            .O(N__40457),
            .I(N__40454));
    Odrv4 I__8674 (
            .O(N__40454),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__8673 (
            .O(N__40451),
            .I(N__40448));
    InMux I__8672 (
            .O(N__40448),
            .I(N__40445));
    LocalMux I__8671 (
            .O(N__40445),
            .I(N__40442));
    Odrv12 I__8670 (
            .O(N__40442),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__8669 (
            .O(N__40439),
            .I(N__40436));
    LocalMux I__8668 (
            .O(N__40436),
            .I(N__40433));
    Span4Mux_h I__8667 (
            .O(N__40433),
            .I(N__40430));
    Odrv4 I__8666 (
            .O(N__40430),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__8665 (
            .O(N__40427),
            .I(N__40424));
    InMux I__8664 (
            .O(N__40424),
            .I(N__40421));
    LocalMux I__8663 (
            .O(N__40421),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__8662 (
            .O(N__40418),
            .I(N__40415));
    LocalMux I__8661 (
            .O(N__40415),
            .I(N__40412));
    Span4Mux_v I__8660 (
            .O(N__40412),
            .I(N__40409));
    Odrv4 I__8659 (
            .O(N__40409),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__8658 (
            .O(N__40406),
            .I(N__40403));
    InMux I__8657 (
            .O(N__40403),
            .I(N__40400));
    LocalMux I__8656 (
            .O(N__40400),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__8655 (
            .O(N__40397),
            .I(N__40394));
    LocalMux I__8654 (
            .O(N__40394),
            .I(N__40391));
    Span4Mux_h I__8653 (
            .O(N__40391),
            .I(N__40388));
    Odrv4 I__8652 (
            .O(N__40388),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__8651 (
            .O(N__40385),
            .I(N__40382));
    InMux I__8650 (
            .O(N__40382),
            .I(N__40379));
    LocalMux I__8649 (
            .O(N__40379),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__8648 (
            .O(N__40376),
            .I(N__40373));
    LocalMux I__8647 (
            .O(N__40373),
            .I(N__40370));
    Odrv12 I__8646 (
            .O(N__40370),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__8645 (
            .O(N__40367),
            .I(N__40364));
    InMux I__8644 (
            .O(N__40364),
            .I(N__40361));
    LocalMux I__8643 (
            .O(N__40361),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__8642 (
            .O(N__40358),
            .I(N__40352));
    InMux I__8641 (
            .O(N__40357),
            .I(N__40352));
    LocalMux I__8640 (
            .O(N__40352),
            .I(N__40349));
    Span4Mux_v I__8639 (
            .O(N__40349),
            .I(N__40346));
    Odrv4 I__8638 (
            .O(N__40346),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ));
    InMux I__8637 (
            .O(N__40343),
            .I(N__40337));
    InMux I__8636 (
            .O(N__40342),
            .I(N__40337));
    LocalMux I__8635 (
            .O(N__40337),
            .I(N__40334));
    Odrv12 I__8634 (
            .O(N__40334),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ));
    InMux I__8633 (
            .O(N__40331),
            .I(N__40328));
    LocalMux I__8632 (
            .O(N__40328),
            .I(N__40325));
    Span4Mux_h I__8631 (
            .O(N__40325),
            .I(N__40319));
    InMux I__8630 (
            .O(N__40324),
            .I(N__40316));
    InMux I__8629 (
            .O(N__40323),
            .I(N__40313));
    InMux I__8628 (
            .O(N__40322),
            .I(N__40310));
    Odrv4 I__8627 (
            .O(N__40319),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    LocalMux I__8626 (
            .O(N__40316),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    LocalMux I__8625 (
            .O(N__40313),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    LocalMux I__8624 (
            .O(N__40310),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__8623 (
            .O(N__40301),
            .I(N__40298));
    LocalMux I__8622 (
            .O(N__40298),
            .I(N__40294));
    InMux I__8621 (
            .O(N__40297),
            .I(N__40290));
    Span4Mux_v I__8620 (
            .O(N__40294),
            .I(N__40287));
    InMux I__8619 (
            .O(N__40293),
            .I(N__40284));
    LocalMux I__8618 (
            .O(N__40290),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    Odrv4 I__8617 (
            .O(N__40287),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    LocalMux I__8616 (
            .O(N__40284),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    InMux I__8615 (
            .O(N__40277),
            .I(N__40272));
    InMux I__8614 (
            .O(N__40276),
            .I(N__40269));
    InMux I__8613 (
            .O(N__40275),
            .I(N__40266));
    LocalMux I__8612 (
            .O(N__40272),
            .I(N__40262));
    LocalMux I__8611 (
            .O(N__40269),
            .I(N__40259));
    LocalMux I__8610 (
            .O(N__40266),
            .I(N__40256));
    InMux I__8609 (
            .O(N__40265),
            .I(N__40253));
    Span4Mux_v I__8608 (
            .O(N__40262),
            .I(N__40250));
    Span4Mux_h I__8607 (
            .O(N__40259),
            .I(N__40247));
    Span4Mux_v I__8606 (
            .O(N__40256),
            .I(N__40244));
    LocalMux I__8605 (
            .O(N__40253),
            .I(N__40241));
    Odrv4 I__8604 (
            .O(N__40250),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__8603 (
            .O(N__40247),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__8602 (
            .O(N__40244),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__8601 (
            .O(N__40241),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__8600 (
            .O(N__40232),
            .I(N__40229));
    LocalMux I__8599 (
            .O(N__40229),
            .I(N__40226));
    Span4Mux_v I__8598 (
            .O(N__40226),
            .I(N__40223));
    Odrv4 I__8597 (
            .O(N__40223),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    CascadeMux I__8596 (
            .O(N__40220),
            .I(N__40217));
    InMux I__8595 (
            .O(N__40217),
            .I(N__40214));
    LocalMux I__8594 (
            .O(N__40214),
            .I(N__40211));
    Odrv4 I__8593 (
            .O(N__40211),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    CascadeMux I__8592 (
            .O(N__40208),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    CascadeMux I__8591 (
            .O(N__40205),
            .I(N__40202));
    InMux I__8590 (
            .O(N__40202),
            .I(N__40199));
    LocalMux I__8589 (
            .O(N__40199),
            .I(N__40196));
    Odrv4 I__8588 (
            .O(N__40196),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__8587 (
            .O(N__40193),
            .I(N__40190));
    LocalMux I__8586 (
            .O(N__40190),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__8585 (
            .O(N__40187),
            .I(N__40184));
    LocalMux I__8584 (
            .O(N__40184),
            .I(N__40181));
    Odrv4 I__8583 (
            .O(N__40181),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__8582 (
            .O(N__40178),
            .I(N__40175));
    InMux I__8581 (
            .O(N__40175),
            .I(N__40172));
    LocalMux I__8580 (
            .O(N__40172),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__8579 (
            .O(N__40169),
            .I(N__40166));
    LocalMux I__8578 (
            .O(N__40166),
            .I(N__40163));
    Odrv4 I__8577 (
            .O(N__40163),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__8576 (
            .O(N__40160),
            .I(N__40157));
    InMux I__8575 (
            .O(N__40157),
            .I(N__40154));
    LocalMux I__8574 (
            .O(N__40154),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__8573 (
            .O(N__40151),
            .I(N__40148));
    InMux I__8572 (
            .O(N__40148),
            .I(N__40145));
    LocalMux I__8571 (
            .O(N__40145),
            .I(N__40142));
    Odrv4 I__8570 (
            .O(N__40142),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__8569 (
            .O(N__40139),
            .I(N__40136));
    LocalMux I__8568 (
            .O(N__40136),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__8567 (
            .O(N__40133),
            .I(N__40130));
    LocalMux I__8566 (
            .O(N__40130),
            .I(N__40127));
    Odrv4 I__8565 (
            .O(N__40127),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__8564 (
            .O(N__40124),
            .I(N__40121));
    LocalMux I__8563 (
            .O(N__40121),
            .I(N__40115));
    InMux I__8562 (
            .O(N__40120),
            .I(N__40112));
    InMux I__8561 (
            .O(N__40119),
            .I(N__40109));
    InMux I__8560 (
            .O(N__40118),
            .I(N__40106));
    Odrv4 I__8559 (
            .O(N__40115),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__8558 (
            .O(N__40112),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__8557 (
            .O(N__40109),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__8556 (
            .O(N__40106),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__8555 (
            .O(N__40097),
            .I(N__40094));
    LocalMux I__8554 (
            .O(N__40094),
            .I(N__40090));
    InMux I__8553 (
            .O(N__40093),
            .I(N__40086));
    Span4Mux_h I__8552 (
            .O(N__40090),
            .I(N__40083));
    InMux I__8551 (
            .O(N__40089),
            .I(N__40080));
    LocalMux I__8550 (
            .O(N__40086),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    Odrv4 I__8549 (
            .O(N__40083),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    LocalMux I__8548 (
            .O(N__40080),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    InMux I__8547 (
            .O(N__40073),
            .I(N__40069));
    InMux I__8546 (
            .O(N__40072),
            .I(N__40066));
    LocalMux I__8545 (
            .O(N__40069),
            .I(N__40061));
    LocalMux I__8544 (
            .O(N__40066),
            .I(N__40058));
    InMux I__8543 (
            .O(N__40065),
            .I(N__40055));
    InMux I__8542 (
            .O(N__40064),
            .I(N__40052));
    Odrv4 I__8541 (
            .O(N__40061),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__8540 (
            .O(N__40058),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    LocalMux I__8539 (
            .O(N__40055),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    LocalMux I__8538 (
            .O(N__40052),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__8537 (
            .O(N__40043),
            .I(N__40040));
    LocalMux I__8536 (
            .O(N__40040),
            .I(N__40036));
    InMux I__8535 (
            .O(N__40039),
            .I(N__40032));
    Span4Mux_h I__8534 (
            .O(N__40036),
            .I(N__40029));
    InMux I__8533 (
            .O(N__40035),
            .I(N__40026));
    LocalMux I__8532 (
            .O(N__40032),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    Odrv4 I__8531 (
            .O(N__40029),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    LocalMux I__8530 (
            .O(N__40026),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    InMux I__8529 (
            .O(N__40019),
            .I(N__40016));
    LocalMux I__8528 (
            .O(N__40016),
            .I(N__40013));
    Odrv12 I__8527 (
            .O(N__40013),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__8526 (
            .O(N__40010),
            .I(N__40003));
    InMux I__8525 (
            .O(N__40009),
            .I(N__40003));
    InMux I__8524 (
            .O(N__40008),
            .I(N__39999));
    LocalMux I__8523 (
            .O(N__40003),
            .I(N__39996));
    InMux I__8522 (
            .O(N__40002),
            .I(N__39993));
    LocalMux I__8521 (
            .O(N__39999),
            .I(N__39990));
    Span4Mux_h I__8520 (
            .O(N__39996),
            .I(N__39985));
    LocalMux I__8519 (
            .O(N__39993),
            .I(N__39985));
    Odrv4 I__8518 (
            .O(N__39990),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__8517 (
            .O(N__39985),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    CascadeMux I__8516 (
            .O(N__39980),
            .I(N__39975));
    InMux I__8515 (
            .O(N__39979),
            .I(N__39972));
    InMux I__8514 (
            .O(N__39978),
            .I(N__39967));
    InMux I__8513 (
            .O(N__39975),
            .I(N__39967));
    LocalMux I__8512 (
            .O(N__39972),
            .I(N__39964));
    LocalMux I__8511 (
            .O(N__39967),
            .I(N__39961));
    Span4Mux_v I__8510 (
            .O(N__39964),
            .I(N__39958));
    Odrv4 I__8509 (
            .O(N__39961),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__8508 (
            .O(N__39958),
            .I(\current_shift_inst.un4_control_input1_23 ));
    CascadeMux I__8507 (
            .O(N__39953),
            .I(N__39950));
    InMux I__8506 (
            .O(N__39950),
            .I(N__39946));
    InMux I__8505 (
            .O(N__39949),
            .I(N__39943));
    LocalMux I__8504 (
            .O(N__39946),
            .I(N__39940));
    LocalMux I__8503 (
            .O(N__39943),
            .I(N__39935));
    Span4Mux_h I__8502 (
            .O(N__39940),
            .I(N__39932));
    InMux I__8501 (
            .O(N__39939),
            .I(N__39929));
    InMux I__8500 (
            .O(N__39938),
            .I(N__39926));
    Span4Mux_h I__8499 (
            .O(N__39935),
            .I(N__39923));
    Span4Mux_v I__8498 (
            .O(N__39932),
            .I(N__39920));
    LocalMux I__8497 (
            .O(N__39929),
            .I(N__39915));
    LocalMux I__8496 (
            .O(N__39926),
            .I(N__39915));
    Odrv4 I__8495 (
            .O(N__39923),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__8494 (
            .O(N__39920),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv12 I__8493 (
            .O(N__39915),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__8492 (
            .O(N__39908),
            .I(N__39905));
    LocalMux I__8491 (
            .O(N__39905),
            .I(N__39900));
    InMux I__8490 (
            .O(N__39904),
            .I(N__39897));
    InMux I__8489 (
            .O(N__39903),
            .I(N__39894));
    Span4Mux_v I__8488 (
            .O(N__39900),
            .I(N__39891));
    LocalMux I__8487 (
            .O(N__39897),
            .I(N__39886));
    LocalMux I__8486 (
            .O(N__39894),
            .I(N__39886));
    Odrv4 I__8485 (
            .O(N__39891),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv12 I__8484 (
            .O(N__39886),
            .I(\current_shift_inst.un4_control_input1_25 ));
    CascadeMux I__8483 (
            .O(N__39881),
            .I(N__39878));
    InMux I__8482 (
            .O(N__39878),
            .I(N__39875));
    LocalMux I__8481 (
            .O(N__39875),
            .I(N__39872));
    Span4Mux_h I__8480 (
            .O(N__39872),
            .I(N__39869));
    Span4Mux_v I__8479 (
            .O(N__39869),
            .I(N__39866));
    Odrv4 I__8478 (
            .O(N__39866),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ));
    InMux I__8477 (
            .O(N__39863),
            .I(N__39860));
    LocalMux I__8476 (
            .O(N__39860),
            .I(N__39857));
    Span4Mux_s1_v I__8475 (
            .O(N__39857),
            .I(N__39853));
    InMux I__8474 (
            .O(N__39856),
            .I(N__39850));
    Span4Mux_h I__8473 (
            .O(N__39853),
            .I(N__39847));
    LocalMux I__8472 (
            .O(N__39850),
            .I(N__39840));
    Sp12to4 I__8471 (
            .O(N__39847),
            .I(N__39840));
    InMux I__8470 (
            .O(N__39846),
            .I(N__39836));
    InMux I__8469 (
            .O(N__39845),
            .I(N__39833));
    Span12Mux_s10_v I__8468 (
            .O(N__39840),
            .I(N__39830));
    InMux I__8467 (
            .O(N__39839),
            .I(N__39827));
    LocalMux I__8466 (
            .O(N__39836),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__8465 (
            .O(N__39833),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__8464 (
            .O(N__39830),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__8463 (
            .O(N__39827),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__8462 (
            .O(N__39818),
            .I(N__39815));
    LocalMux I__8461 (
            .O(N__39815),
            .I(N__39812));
    Span4Mux_s0_v I__8460 (
            .O(N__39812),
            .I(N__39808));
    InMux I__8459 (
            .O(N__39811),
            .I(N__39805));
    Odrv4 I__8458 (
            .O(N__39808),
            .I(T23_c));
    LocalMux I__8457 (
            .O(N__39805),
            .I(T23_c));
    InMux I__8456 (
            .O(N__39800),
            .I(N__39796));
    InMux I__8455 (
            .O(N__39799),
            .I(N__39793));
    LocalMux I__8454 (
            .O(N__39796),
            .I(N__39789));
    LocalMux I__8453 (
            .O(N__39793),
            .I(N__39786));
    InMux I__8452 (
            .O(N__39792),
            .I(N__39783));
    Span4Mux_h I__8451 (
            .O(N__39789),
            .I(N__39780));
    Span4Mux_v I__8450 (
            .O(N__39786),
            .I(N__39777));
    LocalMux I__8449 (
            .O(N__39783),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv4 I__8448 (
            .O(N__39780),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv4 I__8447 (
            .O(N__39777),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    InMux I__8446 (
            .O(N__39770),
            .I(N__39764));
    InMux I__8445 (
            .O(N__39769),
            .I(N__39761));
    InMux I__8444 (
            .O(N__39768),
            .I(N__39758));
    InMux I__8443 (
            .O(N__39767),
            .I(N__39755));
    LocalMux I__8442 (
            .O(N__39764),
            .I(N__39752));
    LocalMux I__8441 (
            .O(N__39761),
            .I(N__39747));
    LocalMux I__8440 (
            .O(N__39758),
            .I(N__39747));
    LocalMux I__8439 (
            .O(N__39755),
            .I(N__39744));
    Span4Mux_h I__8438 (
            .O(N__39752),
            .I(N__39739));
    Span4Mux_v I__8437 (
            .O(N__39747),
            .I(N__39739));
    Span4Mux_v I__8436 (
            .O(N__39744),
            .I(N__39736));
    Odrv4 I__8435 (
            .O(N__39739),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    Odrv4 I__8434 (
            .O(N__39736),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__8433 (
            .O(N__39731),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__8432 (
            .O(N__39728),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__8431 (
            .O(N__39725),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__8430 (
            .O(N__39722),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__8429 (
            .O(N__39719),
            .I(N__39716));
    LocalMux I__8428 (
            .O(N__39716),
            .I(N__39713));
    Odrv12 I__8427 (
            .O(N__39713),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    CascadeMux I__8426 (
            .O(N__39710),
            .I(N__39707));
    InMux I__8425 (
            .O(N__39707),
            .I(N__39704));
    LocalMux I__8424 (
            .O(N__39704),
            .I(N__39701));
    Span4Mux_h I__8423 (
            .O(N__39701),
            .I(N__39696));
    InMux I__8422 (
            .O(N__39700),
            .I(N__39691));
    InMux I__8421 (
            .O(N__39699),
            .I(N__39691));
    Span4Mux_v I__8420 (
            .O(N__39696),
            .I(N__39687));
    LocalMux I__8419 (
            .O(N__39691),
            .I(N__39684));
    InMux I__8418 (
            .O(N__39690),
            .I(N__39681));
    Odrv4 I__8417 (
            .O(N__39687),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__8416 (
            .O(N__39684),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__8415 (
            .O(N__39681),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__8414 (
            .O(N__39674),
            .I(N__39671));
    LocalMux I__8413 (
            .O(N__39671),
            .I(N__39668));
    Odrv12 I__8412 (
            .O(N__39668),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__8411 (
            .O(N__39665),
            .I(N__39662));
    LocalMux I__8410 (
            .O(N__39662),
            .I(N__39659));
    Odrv12 I__8409 (
            .O(N__39659),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__8408 (
            .O(N__39656),
            .I(N__39652));
    CascadeMux I__8407 (
            .O(N__39655),
            .I(N__39649));
    LocalMux I__8406 (
            .O(N__39652),
            .I(N__39646));
    InMux I__8405 (
            .O(N__39649),
            .I(N__39643));
    Span4Mux_h I__8404 (
            .O(N__39646),
            .I(N__39636));
    LocalMux I__8403 (
            .O(N__39643),
            .I(N__39636));
    InMux I__8402 (
            .O(N__39642),
            .I(N__39633));
    InMux I__8401 (
            .O(N__39641),
            .I(N__39630));
    Odrv4 I__8400 (
            .O(N__39636),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__8399 (
            .O(N__39633),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__8398 (
            .O(N__39630),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__8397 (
            .O(N__39623),
            .I(N__39620));
    LocalMux I__8396 (
            .O(N__39620),
            .I(N__39615));
    InMux I__8395 (
            .O(N__39619),
            .I(N__39612));
    InMux I__8394 (
            .O(N__39618),
            .I(N__39609));
    Span4Mux_v I__8393 (
            .O(N__39615),
            .I(N__39606));
    LocalMux I__8392 (
            .O(N__39612),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__8391 (
            .O(N__39609),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv4 I__8390 (
            .O(N__39606),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__8389 (
            .O(N__39599),
            .I(N__39594));
    InMux I__8388 (
            .O(N__39598),
            .I(N__39591));
    InMux I__8387 (
            .O(N__39597),
            .I(N__39588));
    LocalMux I__8386 (
            .O(N__39594),
            .I(N__39585));
    LocalMux I__8385 (
            .O(N__39591),
            .I(N__39582));
    LocalMux I__8384 (
            .O(N__39588),
            .I(N__39579));
    Span4Mux_h I__8383 (
            .O(N__39585),
            .I(N__39576));
    Span4Mux_v I__8382 (
            .O(N__39582),
            .I(N__39573));
    Odrv4 I__8381 (
            .O(N__39579),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__8380 (
            .O(N__39576),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__8379 (
            .O(N__39573),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__8378 (
            .O(N__39566),
            .I(bfn_16_21_0_));
    InMux I__8377 (
            .O(N__39563),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__8376 (
            .O(N__39560),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__8375 (
            .O(N__39557),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__8374 (
            .O(N__39554),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__8373 (
            .O(N__39551),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__8372 (
            .O(N__39548),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__8371 (
            .O(N__39545),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__8370 (
            .O(N__39542),
            .I(bfn_16_22_0_));
    InMux I__8369 (
            .O(N__39539),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__8368 (
            .O(N__39536),
            .I(bfn_16_20_0_));
    InMux I__8367 (
            .O(N__39533),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__8366 (
            .O(N__39530),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__8365 (
            .O(N__39527),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__8364 (
            .O(N__39524),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__8363 (
            .O(N__39521),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__8362 (
            .O(N__39518),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__8361 (
            .O(N__39515),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__8360 (
            .O(N__39512),
            .I(\current_shift_inst.un4_control_input1_31 ));
    InMux I__8359 (
            .O(N__39509),
            .I(N__39506));
    LocalMux I__8358 (
            .O(N__39506),
            .I(N__39503));
    Odrv12 I__8357 (
            .O(N__39503),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__8356 (
            .O(N__39500),
            .I(N__39497));
    LocalMux I__8355 (
            .O(N__39497),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__8354 (
            .O(N__39494),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__8353 (
            .O(N__39491),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__8352 (
            .O(N__39488),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__8351 (
            .O(N__39485),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__8350 (
            .O(N__39482),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__8349 (
            .O(N__39479),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__8348 (
            .O(N__39476),
            .I(N__39473));
    LocalMux I__8347 (
            .O(N__39473),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__8346 (
            .O(N__39470),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__8345 (
            .O(N__39467),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__8344 (
            .O(N__39464),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__8343 (
            .O(N__39461),
            .I(N__39458));
    LocalMux I__8342 (
            .O(N__39458),
            .I(N__39455));
    Odrv4 I__8341 (
            .O(N__39455),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__8340 (
            .O(N__39452),
            .I(bfn_16_18_0_));
    InMux I__8339 (
            .O(N__39449),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__8338 (
            .O(N__39446),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__8337 (
            .O(N__39443),
            .I(N__39439));
    CascadeMux I__8336 (
            .O(N__39442),
            .I(N__39436));
    LocalMux I__8335 (
            .O(N__39439),
            .I(N__39432));
    InMux I__8334 (
            .O(N__39436),
            .I(N__39427));
    InMux I__8333 (
            .O(N__39435),
            .I(N__39427));
    Odrv12 I__8332 (
            .O(N__39432),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__8331 (
            .O(N__39427),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__8330 (
            .O(N__39422),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__8329 (
            .O(N__39419),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__8328 (
            .O(N__39416),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__8327 (
            .O(N__39413),
            .I(N__39410));
    LocalMux I__8326 (
            .O(N__39410),
            .I(N__39407));
    Odrv4 I__8325 (
            .O(N__39407),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__8324 (
            .O(N__39404),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__8323 (
            .O(N__39401),
            .I(N__39398));
    LocalMux I__8322 (
            .O(N__39398),
            .I(N__39395));
    Span4Mux_h I__8321 (
            .O(N__39395),
            .I(N__39392));
    Odrv4 I__8320 (
            .O(N__39392),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__8319 (
            .O(N__39389),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__8318 (
            .O(N__39386),
            .I(N__39383));
    LocalMux I__8317 (
            .O(N__39383),
            .I(N__39380));
    Span4Mux_h I__8316 (
            .O(N__39380),
            .I(N__39377));
    Odrv4 I__8315 (
            .O(N__39377),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__8314 (
            .O(N__39374),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__8313 (
            .O(N__39371),
            .I(bfn_16_17_0_));
    InMux I__8312 (
            .O(N__39368),
            .I(N__39365));
    LocalMux I__8311 (
            .O(N__39365),
            .I(N__39362));
    Odrv4 I__8310 (
            .O(N__39362),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__8309 (
            .O(N__39359),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__8308 (
            .O(N__39356),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__8307 (
            .O(N__39353),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__8306 (
            .O(N__39350),
            .I(N__39347));
    LocalMux I__8305 (
            .O(N__39347),
            .I(N__39344));
    Span4Mux_v I__8304 (
            .O(N__39344),
            .I(N__39341));
    Odrv4 I__8303 (
            .O(N__39341),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__8302 (
            .O(N__39338),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__8301 (
            .O(N__39335),
            .I(N__39332));
    LocalMux I__8300 (
            .O(N__39332),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__8299 (
            .O(N__39329),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__8298 (
            .O(N__39326),
            .I(N__39323));
    LocalMux I__8297 (
            .O(N__39323),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__8296 (
            .O(N__39320),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__8295 (
            .O(N__39317),
            .I(N__39314));
    LocalMux I__8294 (
            .O(N__39314),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__8293 (
            .O(N__39311),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__8292 (
            .O(N__39308),
            .I(N__39305));
    LocalMux I__8291 (
            .O(N__39305),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__8290 (
            .O(N__39302),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__8289 (
            .O(N__39299),
            .I(N__39296));
    LocalMux I__8288 (
            .O(N__39296),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__8287 (
            .O(N__39293),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__8286 (
            .O(N__39290),
            .I(bfn_16_16_0_));
    InMux I__8285 (
            .O(N__39287),
            .I(N__39284));
    LocalMux I__8284 (
            .O(N__39284),
            .I(N__39281));
    Span4Mux_h I__8283 (
            .O(N__39281),
            .I(N__39278));
    Odrv4 I__8282 (
            .O(N__39278),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__8281 (
            .O(N__39275),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__8280 (
            .O(N__39272),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__8279 (
            .O(N__39269),
            .I(N__39266));
    LocalMux I__8278 (
            .O(N__39266),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__8277 (
            .O(N__39263),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__8276 (
            .O(N__39260),
            .I(N__39257));
    LocalMux I__8275 (
            .O(N__39257),
            .I(N__39254));
    Span4Mux_h I__8274 (
            .O(N__39254),
            .I(N__39251));
    Span4Mux_v I__8273 (
            .O(N__39251),
            .I(N__39248));
    Odrv4 I__8272 (
            .O(N__39248),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__8271 (
            .O(N__39245),
            .I(N__39242));
    LocalMux I__8270 (
            .O(N__39242),
            .I(N__39239));
    Span4Mux_h I__8269 (
            .O(N__39239),
            .I(N__39236));
    Odrv4 I__8268 (
            .O(N__39236),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ));
    InMux I__8267 (
            .O(N__39233),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__8266 (
            .O(N__39230),
            .I(N__39227));
    LocalMux I__8265 (
            .O(N__39227),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__8264 (
            .O(N__39224),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__8263 (
            .O(N__39221),
            .I(N__39218));
    LocalMux I__8262 (
            .O(N__39218),
            .I(N__39214));
    InMux I__8261 (
            .O(N__39217),
            .I(N__39211));
    Span4Mux_v I__8260 (
            .O(N__39214),
            .I(N__39208));
    LocalMux I__8259 (
            .O(N__39211),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv4 I__8258 (
            .O(N__39208),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__8257 (
            .O(N__39203),
            .I(N__39200));
    InMux I__8256 (
            .O(N__39200),
            .I(N__39195));
    InMux I__8255 (
            .O(N__39199),
            .I(N__39192));
    InMux I__8254 (
            .O(N__39198),
            .I(N__39189));
    LocalMux I__8253 (
            .O(N__39195),
            .I(N__39184));
    LocalMux I__8252 (
            .O(N__39192),
            .I(N__39184));
    LocalMux I__8251 (
            .O(N__39189),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv12 I__8250 (
            .O(N__39184),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__8249 (
            .O(N__39179),
            .I(N__39176));
    LocalMux I__8248 (
            .O(N__39176),
            .I(N__39170));
    InMux I__8247 (
            .O(N__39175),
            .I(N__39167));
    InMux I__8246 (
            .O(N__39174),
            .I(N__39162));
    InMux I__8245 (
            .O(N__39173),
            .I(N__39162));
    Span4Mux_h I__8244 (
            .O(N__39170),
            .I(N__39159));
    LocalMux I__8243 (
            .O(N__39167),
            .I(N__39156));
    LocalMux I__8242 (
            .O(N__39162),
            .I(N__39153));
    Span4Mux_v I__8241 (
            .O(N__39159),
            .I(N__39150));
    Span4Mux_v I__8240 (
            .O(N__39156),
            .I(N__39147));
    Span4Mux_h I__8239 (
            .O(N__39153),
            .I(N__39144));
    Odrv4 I__8238 (
            .O(N__39150),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__8237 (
            .O(N__39147),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__8236 (
            .O(N__39144),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__8235 (
            .O(N__39137),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__8234 (
            .O(N__39134),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__8233 (
            .O(N__39131),
            .I(N__39128));
    LocalMux I__8232 (
            .O(N__39128),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    CascadeMux I__8231 (
            .O(N__39125),
            .I(N__39121));
    InMux I__8230 (
            .O(N__39124),
            .I(N__39116));
    InMux I__8229 (
            .O(N__39121),
            .I(N__39116));
    LocalMux I__8228 (
            .O(N__39116),
            .I(N__39112));
    InMux I__8227 (
            .O(N__39115),
            .I(N__39109));
    Span4Mux_h I__8226 (
            .O(N__39112),
            .I(N__39106));
    LocalMux I__8225 (
            .O(N__39109),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__8224 (
            .O(N__39106),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__8223 (
            .O(N__39101),
            .I(N__39096));
    InMux I__8222 (
            .O(N__39100),
            .I(N__39093));
    InMux I__8221 (
            .O(N__39099),
            .I(N__39088));
    InMux I__8220 (
            .O(N__39096),
            .I(N__39088));
    LocalMux I__8219 (
            .O(N__39093),
            .I(N__39083));
    LocalMux I__8218 (
            .O(N__39088),
            .I(N__39083));
    Odrv4 I__8217 (
            .O(N__39083),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__8216 (
            .O(N__39080),
            .I(N__39077));
    InMux I__8215 (
            .O(N__39077),
            .I(N__39074));
    LocalMux I__8214 (
            .O(N__39074),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    InMux I__8213 (
            .O(N__39071),
            .I(N__39065));
    InMux I__8212 (
            .O(N__39070),
            .I(N__39065));
    LocalMux I__8211 (
            .O(N__39065),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    InMux I__8210 (
            .O(N__39062),
            .I(N__39059));
    LocalMux I__8209 (
            .O(N__39059),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    InMux I__8208 (
            .O(N__39056),
            .I(N__39053));
    LocalMux I__8207 (
            .O(N__39053),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    InMux I__8206 (
            .O(N__39050),
            .I(N__39043));
    InMux I__8205 (
            .O(N__39049),
            .I(N__39043));
    InMux I__8204 (
            .O(N__39048),
            .I(N__39040));
    LocalMux I__8203 (
            .O(N__39043),
            .I(N__39037));
    LocalMux I__8202 (
            .O(N__39040),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv12 I__8201 (
            .O(N__39037),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__8200 (
            .O(N__39032),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__8199 (
            .O(N__39029),
            .I(N__39026));
    InMux I__8198 (
            .O(N__39026),
            .I(N__39021));
    InMux I__8197 (
            .O(N__39025),
            .I(N__39018));
    InMux I__8196 (
            .O(N__39024),
            .I(N__39015));
    LocalMux I__8195 (
            .O(N__39021),
            .I(N__39010));
    LocalMux I__8194 (
            .O(N__39018),
            .I(N__39010));
    LocalMux I__8193 (
            .O(N__39015),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv12 I__8192 (
            .O(N__39010),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__8191 (
            .O(N__39005),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__8190 (
            .O(N__39002),
            .I(N__38998));
    InMux I__8189 (
            .O(N__39001),
            .I(N__38995));
    InMux I__8188 (
            .O(N__38998),
            .I(N__38992));
    LocalMux I__8187 (
            .O(N__38995),
            .I(N__38988));
    LocalMux I__8186 (
            .O(N__38992),
            .I(N__38985));
    InMux I__8185 (
            .O(N__38991),
            .I(N__38982));
    Span4Mux_v I__8184 (
            .O(N__38988),
            .I(N__38977));
    Span4Mux_v I__8183 (
            .O(N__38985),
            .I(N__38977));
    LocalMux I__8182 (
            .O(N__38982),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv4 I__8181 (
            .O(N__38977),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__8180 (
            .O(N__38972),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__8179 (
            .O(N__38969),
            .I(N__38963));
    InMux I__8178 (
            .O(N__38968),
            .I(N__38963));
    LocalMux I__8177 (
            .O(N__38963),
            .I(N__38959));
    InMux I__8176 (
            .O(N__38962),
            .I(N__38956));
    Span4Mux_v I__8175 (
            .O(N__38959),
            .I(N__38953));
    LocalMux I__8174 (
            .O(N__38956),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__8173 (
            .O(N__38953),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__8172 (
            .O(N__38948),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__8171 (
            .O(N__38945),
            .I(N__38941));
    CascadeMux I__8170 (
            .O(N__38944),
            .I(N__38938));
    InMux I__8169 (
            .O(N__38941),
            .I(N__38933));
    InMux I__8168 (
            .O(N__38938),
            .I(N__38933));
    LocalMux I__8167 (
            .O(N__38933),
            .I(N__38929));
    InMux I__8166 (
            .O(N__38932),
            .I(N__38926));
    Span4Mux_v I__8165 (
            .O(N__38929),
            .I(N__38923));
    LocalMux I__8164 (
            .O(N__38926),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv4 I__8163 (
            .O(N__38923),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__8162 (
            .O(N__38918),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__8161 (
            .O(N__38915),
            .I(N__38911));
    CascadeMux I__8160 (
            .O(N__38914),
            .I(N__38908));
    InMux I__8159 (
            .O(N__38911),
            .I(N__38905));
    InMux I__8158 (
            .O(N__38908),
            .I(N__38902));
    LocalMux I__8157 (
            .O(N__38905),
            .I(N__38896));
    LocalMux I__8156 (
            .O(N__38902),
            .I(N__38896));
    InMux I__8155 (
            .O(N__38901),
            .I(N__38893));
    Span4Mux_v I__8154 (
            .O(N__38896),
            .I(N__38890));
    LocalMux I__8153 (
            .O(N__38893),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__8152 (
            .O(N__38890),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__8151 (
            .O(N__38885),
            .I(bfn_16_12_0_));
    CascadeMux I__8150 (
            .O(N__38882),
            .I(N__38879));
    InMux I__8149 (
            .O(N__38879),
            .I(N__38874));
    InMux I__8148 (
            .O(N__38878),
            .I(N__38871));
    InMux I__8147 (
            .O(N__38877),
            .I(N__38868));
    LocalMux I__8146 (
            .O(N__38874),
            .I(N__38863));
    LocalMux I__8145 (
            .O(N__38871),
            .I(N__38863));
    LocalMux I__8144 (
            .O(N__38868),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv12 I__8143 (
            .O(N__38863),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__8142 (
            .O(N__38858),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__8141 (
            .O(N__38855),
            .I(N__38848));
    InMux I__8140 (
            .O(N__38854),
            .I(N__38848));
    InMux I__8139 (
            .O(N__38853),
            .I(N__38845));
    LocalMux I__8138 (
            .O(N__38848),
            .I(N__38842));
    LocalMux I__8137 (
            .O(N__38845),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv12 I__8136 (
            .O(N__38842),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    CascadeMux I__8135 (
            .O(N__38837),
            .I(N__38834));
    InMux I__8134 (
            .O(N__38834),
            .I(N__38830));
    InMux I__8133 (
            .O(N__38833),
            .I(N__38827));
    LocalMux I__8132 (
            .O(N__38830),
            .I(N__38824));
    LocalMux I__8131 (
            .O(N__38827),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv12 I__8130 (
            .O(N__38824),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__8129 (
            .O(N__38819),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__8128 (
            .O(N__38816),
            .I(N__38811));
    InMux I__8127 (
            .O(N__38815),
            .I(N__38808));
    InMux I__8126 (
            .O(N__38814),
            .I(N__38805));
    LocalMux I__8125 (
            .O(N__38811),
            .I(N__38802));
    LocalMux I__8124 (
            .O(N__38808),
            .I(N__38797));
    LocalMux I__8123 (
            .O(N__38805),
            .I(N__38797));
    Span4Mux_v I__8122 (
            .O(N__38802),
            .I(N__38791));
    Span4Mux_v I__8121 (
            .O(N__38797),
            .I(N__38791));
    InMux I__8120 (
            .O(N__38796),
            .I(N__38788));
    Odrv4 I__8119 (
            .O(N__38791),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__8118 (
            .O(N__38788),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__8117 (
            .O(N__38783),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__8116 (
            .O(N__38780),
            .I(N__38774));
    InMux I__8115 (
            .O(N__38779),
            .I(N__38774));
    LocalMux I__8114 (
            .O(N__38774),
            .I(N__38770));
    InMux I__8113 (
            .O(N__38773),
            .I(N__38767));
    Span4Mux_v I__8112 (
            .O(N__38770),
            .I(N__38764));
    LocalMux I__8111 (
            .O(N__38767),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__8110 (
            .O(N__38764),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__8109 (
            .O(N__38759),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__8108 (
            .O(N__38756),
            .I(N__38752));
    CascadeMux I__8107 (
            .O(N__38755),
            .I(N__38749));
    InMux I__8106 (
            .O(N__38752),
            .I(N__38743));
    InMux I__8105 (
            .O(N__38749),
            .I(N__38743));
    InMux I__8104 (
            .O(N__38748),
            .I(N__38740));
    LocalMux I__8103 (
            .O(N__38743),
            .I(N__38737));
    LocalMux I__8102 (
            .O(N__38740),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv12 I__8101 (
            .O(N__38737),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__8100 (
            .O(N__38732),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__8099 (
            .O(N__38729),
            .I(N__38725));
    CascadeMux I__8098 (
            .O(N__38728),
            .I(N__38722));
    InMux I__8097 (
            .O(N__38725),
            .I(N__38716));
    InMux I__8096 (
            .O(N__38722),
            .I(N__38716));
    InMux I__8095 (
            .O(N__38721),
            .I(N__38713));
    LocalMux I__8094 (
            .O(N__38716),
            .I(N__38710));
    LocalMux I__8093 (
            .O(N__38713),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv12 I__8092 (
            .O(N__38710),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__8091 (
            .O(N__38705),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__8090 (
            .O(N__38702),
            .I(N__38696));
    InMux I__8089 (
            .O(N__38701),
            .I(N__38696));
    LocalMux I__8088 (
            .O(N__38696),
            .I(N__38692));
    InMux I__8087 (
            .O(N__38695),
            .I(N__38689));
    Span4Mux_v I__8086 (
            .O(N__38692),
            .I(N__38686));
    LocalMux I__8085 (
            .O(N__38689),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__8084 (
            .O(N__38686),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__8083 (
            .O(N__38681),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__8082 (
            .O(N__38678),
            .I(N__38675));
    InMux I__8081 (
            .O(N__38675),
            .I(N__38670));
    InMux I__8080 (
            .O(N__38674),
            .I(N__38667));
    InMux I__8079 (
            .O(N__38673),
            .I(N__38664));
    LocalMux I__8078 (
            .O(N__38670),
            .I(N__38659));
    LocalMux I__8077 (
            .O(N__38667),
            .I(N__38659));
    LocalMux I__8076 (
            .O(N__38664),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv12 I__8075 (
            .O(N__38659),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__8074 (
            .O(N__38654),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__8073 (
            .O(N__38651),
            .I(N__38647));
    InMux I__8072 (
            .O(N__38650),
            .I(N__38644));
    InMux I__8071 (
            .O(N__38647),
            .I(N__38641));
    LocalMux I__8070 (
            .O(N__38644),
            .I(N__38635));
    LocalMux I__8069 (
            .O(N__38641),
            .I(N__38635));
    InMux I__8068 (
            .O(N__38640),
            .I(N__38632));
    Span4Mux_v I__8067 (
            .O(N__38635),
            .I(N__38629));
    LocalMux I__8066 (
            .O(N__38632),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__8065 (
            .O(N__38629),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__8064 (
            .O(N__38624),
            .I(bfn_16_11_0_));
    CascadeMux I__8063 (
            .O(N__38621),
            .I(N__38618));
    InMux I__8062 (
            .O(N__38618),
            .I(N__38613));
    InMux I__8061 (
            .O(N__38617),
            .I(N__38610));
    InMux I__8060 (
            .O(N__38616),
            .I(N__38607));
    LocalMux I__8059 (
            .O(N__38613),
            .I(N__38602));
    LocalMux I__8058 (
            .O(N__38610),
            .I(N__38602));
    LocalMux I__8057 (
            .O(N__38607),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv12 I__8056 (
            .O(N__38602),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__8055 (
            .O(N__38597),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__8054 (
            .O(N__38594),
            .I(N__38590));
    CascadeMux I__8053 (
            .O(N__38593),
            .I(N__38587));
    InMux I__8052 (
            .O(N__38590),
            .I(N__38581));
    InMux I__8051 (
            .O(N__38587),
            .I(N__38581));
    InMux I__8050 (
            .O(N__38586),
            .I(N__38578));
    LocalMux I__8049 (
            .O(N__38581),
            .I(N__38575));
    LocalMux I__8048 (
            .O(N__38578),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv12 I__8047 (
            .O(N__38575),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__8046 (
            .O(N__38570),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__8045 (
            .O(N__38567),
            .I(N__38563));
    CascadeMux I__8044 (
            .O(N__38566),
            .I(N__38560));
    LocalMux I__8043 (
            .O(N__38563),
            .I(N__38556));
    InMux I__8042 (
            .O(N__38560),
            .I(N__38553));
    InMux I__8041 (
            .O(N__38559),
            .I(N__38550));
    Sp12to4 I__8040 (
            .O(N__38556),
            .I(N__38545));
    LocalMux I__8039 (
            .O(N__38553),
            .I(N__38545));
    LocalMux I__8038 (
            .O(N__38550),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv12 I__8037 (
            .O(N__38545),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__8036 (
            .O(N__38540),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__8035 (
            .O(N__38537),
            .I(N__38531));
    InMux I__8034 (
            .O(N__38536),
            .I(N__38531));
    LocalMux I__8033 (
            .O(N__38531),
            .I(N__38527));
    InMux I__8032 (
            .O(N__38530),
            .I(N__38524));
    Span4Mux_v I__8031 (
            .O(N__38527),
            .I(N__38521));
    LocalMux I__8030 (
            .O(N__38524),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__8029 (
            .O(N__38521),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__8028 (
            .O(N__38516),
            .I(N__38513));
    LocalMux I__8027 (
            .O(N__38513),
            .I(N__38509));
    InMux I__8026 (
            .O(N__38512),
            .I(N__38506));
    Span4Mux_v I__8025 (
            .O(N__38509),
            .I(N__38501));
    LocalMux I__8024 (
            .O(N__38506),
            .I(N__38498));
    InMux I__8023 (
            .O(N__38505),
            .I(N__38495));
    InMux I__8022 (
            .O(N__38504),
            .I(N__38492));
    Odrv4 I__8021 (
            .O(N__38501),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    Odrv4 I__8020 (
            .O(N__38498),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    LocalMux I__8019 (
            .O(N__38495),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    LocalMux I__8018 (
            .O(N__38492),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__8017 (
            .O(N__38483),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__8016 (
            .O(N__38480),
            .I(N__38476));
    CascadeMux I__8015 (
            .O(N__38479),
            .I(N__38473));
    InMux I__8014 (
            .O(N__38476),
            .I(N__38467));
    InMux I__8013 (
            .O(N__38473),
            .I(N__38467));
    InMux I__8012 (
            .O(N__38472),
            .I(N__38464));
    LocalMux I__8011 (
            .O(N__38467),
            .I(N__38461));
    LocalMux I__8010 (
            .O(N__38464),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv12 I__8009 (
            .O(N__38461),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__8008 (
            .O(N__38456),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__8007 (
            .O(N__38453),
            .I(N__38449));
    CascadeMux I__8006 (
            .O(N__38452),
            .I(N__38446));
    InMux I__8005 (
            .O(N__38449),
            .I(N__38440));
    InMux I__8004 (
            .O(N__38446),
            .I(N__38440));
    InMux I__8003 (
            .O(N__38445),
            .I(N__38437));
    LocalMux I__8002 (
            .O(N__38440),
            .I(N__38434));
    LocalMux I__8001 (
            .O(N__38437),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv12 I__8000 (
            .O(N__38434),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__7999 (
            .O(N__38429),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__7998 (
            .O(N__38426),
            .I(N__38420));
    InMux I__7997 (
            .O(N__38425),
            .I(N__38420));
    LocalMux I__7996 (
            .O(N__38420),
            .I(N__38416));
    InMux I__7995 (
            .O(N__38419),
            .I(N__38413));
    Span4Mux_v I__7994 (
            .O(N__38416),
            .I(N__38410));
    LocalMux I__7993 (
            .O(N__38413),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__7992 (
            .O(N__38410),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__7991 (
            .O(N__38405),
            .I(N__38401));
    InMux I__7990 (
            .O(N__38404),
            .I(N__38396));
    LocalMux I__7989 (
            .O(N__38401),
            .I(N__38393));
    CascadeMux I__7988 (
            .O(N__38400),
            .I(N__38390));
    InMux I__7987 (
            .O(N__38399),
            .I(N__38387));
    LocalMux I__7986 (
            .O(N__38396),
            .I(N__38384));
    Span4Mux_v I__7985 (
            .O(N__38393),
            .I(N__38381));
    InMux I__7984 (
            .O(N__38390),
            .I(N__38378));
    LocalMux I__7983 (
            .O(N__38387),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__7982 (
            .O(N__38384),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__7981 (
            .O(N__38381),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    LocalMux I__7980 (
            .O(N__38378),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__7979 (
            .O(N__38369),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__7978 (
            .O(N__38366),
            .I(N__38360));
    InMux I__7977 (
            .O(N__38365),
            .I(N__38360));
    LocalMux I__7976 (
            .O(N__38360),
            .I(N__38356));
    InMux I__7975 (
            .O(N__38359),
            .I(N__38353));
    Span4Mux_v I__7974 (
            .O(N__38356),
            .I(N__38350));
    LocalMux I__7973 (
            .O(N__38353),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__7972 (
            .O(N__38350),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__7971 (
            .O(N__38345),
            .I(N__38342));
    LocalMux I__7970 (
            .O(N__38342),
            .I(N__38339));
    Span4Mux_h I__7969 (
            .O(N__38339),
            .I(N__38333));
    InMux I__7968 (
            .O(N__38338),
            .I(N__38328));
    InMux I__7967 (
            .O(N__38337),
            .I(N__38328));
    InMux I__7966 (
            .O(N__38336),
            .I(N__38325));
    Odrv4 I__7965 (
            .O(N__38333),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__7964 (
            .O(N__38328),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__7963 (
            .O(N__38325),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__7962 (
            .O(N__38318),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__7961 (
            .O(N__38315),
            .I(N__38311));
    CascadeMux I__7960 (
            .O(N__38314),
            .I(N__38308));
    InMux I__7959 (
            .O(N__38311),
            .I(N__38305));
    InMux I__7958 (
            .O(N__38308),
            .I(N__38302));
    LocalMux I__7957 (
            .O(N__38305),
            .I(N__38296));
    LocalMux I__7956 (
            .O(N__38302),
            .I(N__38296));
    InMux I__7955 (
            .O(N__38301),
            .I(N__38293));
    Span4Mux_v I__7954 (
            .O(N__38296),
            .I(N__38290));
    LocalMux I__7953 (
            .O(N__38293),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__7952 (
            .O(N__38290),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__7951 (
            .O(N__38285),
            .I(N__38281));
    InMux I__7950 (
            .O(N__38284),
            .I(N__38278));
    LocalMux I__7949 (
            .O(N__38281),
            .I(N__38275));
    LocalMux I__7948 (
            .O(N__38278),
            .I(N__38270));
    Span4Mux_h I__7947 (
            .O(N__38275),
            .I(N__38267));
    InMux I__7946 (
            .O(N__38274),
            .I(N__38262));
    InMux I__7945 (
            .O(N__38273),
            .I(N__38262));
    Odrv4 I__7944 (
            .O(N__38270),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    Odrv4 I__7943 (
            .O(N__38267),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__7942 (
            .O(N__38262),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__7941 (
            .O(N__38255),
            .I(bfn_16_10_0_));
    CascadeMux I__7940 (
            .O(N__38252),
            .I(N__38248));
    CascadeMux I__7939 (
            .O(N__38251),
            .I(N__38245));
    InMux I__7938 (
            .O(N__38248),
            .I(N__38242));
    InMux I__7937 (
            .O(N__38245),
            .I(N__38239));
    LocalMux I__7936 (
            .O(N__38242),
            .I(N__38233));
    LocalMux I__7935 (
            .O(N__38239),
            .I(N__38233));
    InMux I__7934 (
            .O(N__38238),
            .I(N__38230));
    Span4Mux_v I__7933 (
            .O(N__38233),
            .I(N__38227));
    LocalMux I__7932 (
            .O(N__38230),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__7931 (
            .O(N__38227),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__7930 (
            .O(N__38222),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__7929 (
            .O(N__38219),
            .I(N__38213));
    InMux I__7928 (
            .O(N__38218),
            .I(N__38213));
    LocalMux I__7927 (
            .O(N__38213),
            .I(N__38209));
    InMux I__7926 (
            .O(N__38212),
            .I(N__38206));
    Span4Mux_v I__7925 (
            .O(N__38209),
            .I(N__38203));
    LocalMux I__7924 (
            .O(N__38206),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__7923 (
            .O(N__38203),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__7922 (
            .O(N__38198),
            .I(bfn_16_8_0_));
    InMux I__7921 (
            .O(N__38195),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__7920 (
            .O(N__38192),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__7919 (
            .O(N__38189),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__7918 (
            .O(N__38186),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__7917 (
            .O(N__38183),
            .I(N__38149));
    InMux I__7916 (
            .O(N__38182),
            .I(N__38149));
    InMux I__7915 (
            .O(N__38181),
            .I(N__38140));
    InMux I__7914 (
            .O(N__38180),
            .I(N__38140));
    InMux I__7913 (
            .O(N__38179),
            .I(N__38140));
    InMux I__7912 (
            .O(N__38178),
            .I(N__38140));
    InMux I__7911 (
            .O(N__38177),
            .I(N__38131));
    InMux I__7910 (
            .O(N__38176),
            .I(N__38131));
    InMux I__7909 (
            .O(N__38175),
            .I(N__38131));
    InMux I__7908 (
            .O(N__38174),
            .I(N__38131));
    InMux I__7907 (
            .O(N__38173),
            .I(N__38122));
    InMux I__7906 (
            .O(N__38172),
            .I(N__38122));
    InMux I__7905 (
            .O(N__38171),
            .I(N__38122));
    InMux I__7904 (
            .O(N__38170),
            .I(N__38122));
    InMux I__7903 (
            .O(N__38169),
            .I(N__38113));
    InMux I__7902 (
            .O(N__38168),
            .I(N__38113));
    InMux I__7901 (
            .O(N__38167),
            .I(N__38113));
    InMux I__7900 (
            .O(N__38166),
            .I(N__38113));
    InMux I__7899 (
            .O(N__38165),
            .I(N__38104));
    InMux I__7898 (
            .O(N__38164),
            .I(N__38104));
    InMux I__7897 (
            .O(N__38163),
            .I(N__38104));
    InMux I__7896 (
            .O(N__38162),
            .I(N__38104));
    InMux I__7895 (
            .O(N__38161),
            .I(N__38095));
    InMux I__7894 (
            .O(N__38160),
            .I(N__38095));
    InMux I__7893 (
            .O(N__38159),
            .I(N__38095));
    InMux I__7892 (
            .O(N__38158),
            .I(N__38095));
    InMux I__7891 (
            .O(N__38157),
            .I(N__38086));
    InMux I__7890 (
            .O(N__38156),
            .I(N__38086));
    InMux I__7889 (
            .O(N__38155),
            .I(N__38086));
    InMux I__7888 (
            .O(N__38154),
            .I(N__38086));
    LocalMux I__7887 (
            .O(N__38149),
            .I(N__38081));
    LocalMux I__7886 (
            .O(N__38140),
            .I(N__38081));
    LocalMux I__7885 (
            .O(N__38131),
            .I(N__38068));
    LocalMux I__7884 (
            .O(N__38122),
            .I(N__38068));
    LocalMux I__7883 (
            .O(N__38113),
            .I(N__38068));
    LocalMux I__7882 (
            .O(N__38104),
            .I(N__38068));
    LocalMux I__7881 (
            .O(N__38095),
            .I(N__38068));
    LocalMux I__7880 (
            .O(N__38086),
            .I(N__38068));
    Span4Mux_v I__7879 (
            .O(N__38081),
            .I(N__38063));
    Span4Mux_v I__7878 (
            .O(N__38068),
            .I(N__38063));
    Odrv4 I__7877 (
            .O(N__38063),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__7876 (
            .O(N__38060),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    CEMux I__7875 (
            .O(N__38057),
            .I(N__38051));
    CEMux I__7874 (
            .O(N__38056),
            .I(N__38048));
    CEMux I__7873 (
            .O(N__38055),
            .I(N__38045));
    CEMux I__7872 (
            .O(N__38054),
            .I(N__38042));
    LocalMux I__7871 (
            .O(N__38051),
            .I(N__38039));
    LocalMux I__7870 (
            .O(N__38048),
            .I(N__38036));
    LocalMux I__7869 (
            .O(N__38045),
            .I(N__38033));
    LocalMux I__7868 (
            .O(N__38042),
            .I(N__38030));
    Span4Mux_h I__7867 (
            .O(N__38039),
            .I(N__38027));
    Span4Mux_h I__7866 (
            .O(N__38036),
            .I(N__38024));
    Span4Mux_h I__7865 (
            .O(N__38033),
            .I(N__38021));
    Span4Mux_v I__7864 (
            .O(N__38030),
            .I(N__38018));
    Odrv4 I__7863 (
            .O(N__38027),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    Odrv4 I__7862 (
            .O(N__38024),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    Odrv4 I__7861 (
            .O(N__38021),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    Odrv4 I__7860 (
            .O(N__38018),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    InMux I__7859 (
            .O(N__38009),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__7858 (
            .O(N__38006),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__7857 (
            .O(N__38003),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__7856 (
            .O(N__38000),
            .I(bfn_16_7_0_));
    InMux I__7855 (
            .O(N__37997),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__7854 (
            .O(N__37994),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__7853 (
            .O(N__37991),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__7852 (
            .O(N__37988),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__7851 (
            .O(N__37985),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__7850 (
            .O(N__37982),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__7849 (
            .O(N__37979),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__7848 (
            .O(N__37976),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__7847 (
            .O(N__37973),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__7846 (
            .O(N__37970),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__7845 (
            .O(N__37967),
            .I(bfn_16_6_0_));
    InMux I__7844 (
            .O(N__37964),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__7843 (
            .O(N__37961),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__7842 (
            .O(N__37958),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__7841 (
            .O(N__37955),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__7840 (
            .O(N__37952),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__7839 (
            .O(N__37949),
            .I(N__37944));
    InMux I__7838 (
            .O(N__37948),
            .I(N__37940));
    InMux I__7837 (
            .O(N__37947),
            .I(N__37937));
    LocalMux I__7836 (
            .O(N__37944),
            .I(N__37934));
    InMux I__7835 (
            .O(N__37943),
            .I(N__37931));
    LocalMux I__7834 (
            .O(N__37940),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7833 (
            .O(N__37937),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__7832 (
            .O(N__37934),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7831 (
            .O(N__37931),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__7830 (
            .O(N__37922),
            .I(bfn_16_5_0_));
    InMux I__7829 (
            .O(N__37919),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__7828 (
            .O(N__37916),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__7827 (
            .O(N__37913),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__7826 (
            .O(N__37910),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__7825 (
            .O(N__37907),
            .I(N__37904));
    InMux I__7824 (
            .O(N__37904),
            .I(N__37901));
    LocalMux I__7823 (
            .O(N__37901),
            .I(N__37898));
    Odrv4 I__7822 (
            .O(N__37898),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__7821 (
            .O(N__37895),
            .I(N__37892));
    LocalMux I__7820 (
            .O(N__37892),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    CascadeMux I__7819 (
            .O(N__37889),
            .I(N__37886));
    InMux I__7818 (
            .O(N__37886),
            .I(N__37883));
    LocalMux I__7817 (
            .O(N__37883),
            .I(N__37880));
    Odrv12 I__7816 (
            .O(N__37880),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    CascadeMux I__7815 (
            .O(N__37877),
            .I(N__37874));
    InMux I__7814 (
            .O(N__37874),
            .I(N__37871));
    LocalMux I__7813 (
            .O(N__37871),
            .I(N__37868));
    Span4Mux_v I__7812 (
            .O(N__37868),
            .I(N__37865));
    Span4Mux_h I__7811 (
            .O(N__37865),
            .I(N__37862));
    Odrv4 I__7810 (
            .O(N__37862),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    InMux I__7809 (
            .O(N__37859),
            .I(N__37856));
    LocalMux I__7808 (
            .O(N__37856),
            .I(N__37853));
    Odrv12 I__7807 (
            .O(N__37853),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__7806 (
            .O(N__37850),
            .I(N__37847));
    LocalMux I__7805 (
            .O(N__37847),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ));
    CascadeMux I__7804 (
            .O(N__37844),
            .I(N__37841));
    InMux I__7803 (
            .O(N__37841),
            .I(N__37838));
    LocalMux I__7802 (
            .O(N__37838),
            .I(N__37835));
    Odrv4 I__7801 (
            .O(N__37835),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__7800 (
            .O(N__37832),
            .I(N__37829));
    LocalMux I__7799 (
            .O(N__37829),
            .I(N__37826));
    Odrv12 I__7798 (
            .O(N__37826),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    CascadeMux I__7797 (
            .O(N__37823),
            .I(N__37820));
    InMux I__7796 (
            .O(N__37820),
            .I(N__37817));
    LocalMux I__7795 (
            .O(N__37817),
            .I(N__37814));
    Odrv4 I__7794 (
            .O(N__37814),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__7793 (
            .O(N__37811),
            .I(N__37808));
    LocalMux I__7792 (
            .O(N__37808),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    CascadeMux I__7791 (
            .O(N__37805),
            .I(N__37802));
    InMux I__7790 (
            .O(N__37802),
            .I(N__37799));
    LocalMux I__7789 (
            .O(N__37799),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    CascadeMux I__7788 (
            .O(N__37796),
            .I(N__37793));
    InMux I__7787 (
            .O(N__37793),
            .I(N__37790));
    LocalMux I__7786 (
            .O(N__37790),
            .I(N__37787));
    Span4Mux_h I__7785 (
            .O(N__37787),
            .I(N__37784));
    Odrv4 I__7784 (
            .O(N__37784),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__7783 (
            .O(N__37781),
            .I(N__37778));
    LocalMux I__7782 (
            .O(N__37778),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ));
    CascadeMux I__7781 (
            .O(N__37775),
            .I(N__37772));
    InMux I__7780 (
            .O(N__37772),
            .I(N__37769));
    LocalMux I__7779 (
            .O(N__37769),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ));
    InMux I__7778 (
            .O(N__37766),
            .I(N__37763));
    LocalMux I__7777 (
            .O(N__37763),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ));
    InMux I__7776 (
            .O(N__37760),
            .I(N__37757));
    LocalMux I__7775 (
            .O(N__37757),
            .I(N__37754));
    Odrv12 I__7774 (
            .O(N__37754),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ));
    InMux I__7773 (
            .O(N__37751),
            .I(N__37748));
    LocalMux I__7772 (
            .O(N__37748),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__7771 (
            .O(N__37745),
            .I(N__37742));
    LocalMux I__7770 (
            .O(N__37742),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ));
    CascadeMux I__7769 (
            .O(N__37739),
            .I(N__37736));
    InMux I__7768 (
            .O(N__37736),
            .I(N__37733));
    LocalMux I__7767 (
            .O(N__37733),
            .I(N__37730));
    Span4Mux_h I__7766 (
            .O(N__37730),
            .I(N__37727));
    Odrv4 I__7765 (
            .O(N__37727),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ));
    InMux I__7764 (
            .O(N__37724),
            .I(N__37721));
    LocalMux I__7763 (
            .O(N__37721),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__7762 (
            .O(N__37718),
            .I(N__37715));
    LocalMux I__7761 (
            .O(N__37715),
            .I(N__37712));
    Span4Mux_h I__7760 (
            .O(N__37712),
            .I(N__37709));
    Odrv4 I__7759 (
            .O(N__37709),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ));
    CascadeMux I__7758 (
            .O(N__37706),
            .I(N__37703));
    InMux I__7757 (
            .O(N__37703),
            .I(N__37700));
    LocalMux I__7756 (
            .O(N__37700),
            .I(N__37697));
    Span4Mux_v I__7755 (
            .O(N__37697),
            .I(N__37694));
    Odrv4 I__7754 (
            .O(N__37694),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt24 ));
    InMux I__7753 (
            .O(N__37691),
            .I(N__37688));
    LocalMux I__7752 (
            .O(N__37688),
            .I(N__37685));
    Span4Mux_v I__7751 (
            .O(N__37685),
            .I(N__37682));
    Odrv4 I__7750 (
            .O(N__37682),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    CascadeMux I__7749 (
            .O(N__37679),
            .I(N__37676));
    InMux I__7748 (
            .O(N__37676),
            .I(N__37673));
    LocalMux I__7747 (
            .O(N__37673),
            .I(N__37670));
    Span4Mux_v I__7746 (
            .O(N__37670),
            .I(N__37667));
    Odrv4 I__7745 (
            .O(N__37667),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    InMux I__7744 (
            .O(N__37664),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ));
    InMux I__7743 (
            .O(N__37661),
            .I(N__37658));
    LocalMux I__7742 (
            .O(N__37658),
            .I(N__37653));
    InMux I__7741 (
            .O(N__37657),
            .I(N__37648));
    InMux I__7740 (
            .O(N__37656),
            .I(N__37648));
    Span4Mux_v I__7739 (
            .O(N__37653),
            .I(N__37645));
    LocalMux I__7738 (
            .O(N__37648),
            .I(N__37642));
    Span4Mux_h I__7737 (
            .O(N__37645),
            .I(N__37637));
    Span4Mux_v I__7736 (
            .O(N__37642),
            .I(N__37637));
    Odrv4 I__7735 (
            .O(N__37637),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__7734 (
            .O(N__37634),
            .I(N__37631));
    LocalMux I__7733 (
            .O(N__37631),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ));
    CascadeMux I__7732 (
            .O(N__37628),
            .I(N__37625));
    InMux I__7731 (
            .O(N__37625),
            .I(N__37622));
    LocalMux I__7730 (
            .O(N__37622),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ));
    CascadeMux I__7729 (
            .O(N__37619),
            .I(N__37616));
    InMux I__7728 (
            .O(N__37616),
            .I(N__37613));
    LocalMux I__7727 (
            .O(N__37613),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ));
    InMux I__7726 (
            .O(N__37610),
            .I(N__37607));
    LocalMux I__7725 (
            .O(N__37607),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ));
    InMux I__7724 (
            .O(N__37604),
            .I(N__37601));
    LocalMux I__7723 (
            .O(N__37601),
            .I(N__37598));
    Odrv12 I__7722 (
            .O(N__37598),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    InMux I__7721 (
            .O(N__37595),
            .I(N__37591));
    InMux I__7720 (
            .O(N__37594),
            .I(N__37588));
    LocalMux I__7719 (
            .O(N__37591),
            .I(N__37585));
    LocalMux I__7718 (
            .O(N__37588),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__7717 (
            .O(N__37585),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__7716 (
            .O(N__37580),
            .I(N__37577));
    InMux I__7715 (
            .O(N__37577),
            .I(N__37574));
    LocalMux I__7714 (
            .O(N__37574),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__7713 (
            .O(N__37571),
            .I(N__37567));
    InMux I__7712 (
            .O(N__37570),
            .I(N__37564));
    LocalMux I__7711 (
            .O(N__37567),
            .I(N__37561));
    LocalMux I__7710 (
            .O(N__37564),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__7709 (
            .O(N__37561),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__7708 (
            .O(N__37556),
            .I(N__37553));
    LocalMux I__7707 (
            .O(N__37553),
            .I(N__37550));
    Span4Mux_v I__7706 (
            .O(N__37550),
            .I(N__37547));
    Odrv4 I__7705 (
            .O(N__37547),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__7704 (
            .O(N__37544),
            .I(N__37541));
    InMux I__7703 (
            .O(N__37541),
            .I(N__37538));
    LocalMux I__7702 (
            .O(N__37538),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__7701 (
            .O(N__37535),
            .I(N__37531));
    InMux I__7700 (
            .O(N__37534),
            .I(N__37528));
    LocalMux I__7699 (
            .O(N__37531),
            .I(N__37525));
    LocalMux I__7698 (
            .O(N__37528),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__7697 (
            .O(N__37525),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__7696 (
            .O(N__37520),
            .I(N__37517));
    InMux I__7695 (
            .O(N__37517),
            .I(N__37514));
    LocalMux I__7694 (
            .O(N__37514),
            .I(N__37511));
    Odrv4 I__7693 (
            .O(N__37511),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__7692 (
            .O(N__37508),
            .I(N__37505));
    LocalMux I__7691 (
            .O(N__37505),
            .I(N__37502));
    Span4Mux_v I__7690 (
            .O(N__37502),
            .I(N__37499));
    Odrv4 I__7689 (
            .O(N__37499),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    InMux I__7688 (
            .O(N__37496),
            .I(N__37492));
    InMux I__7687 (
            .O(N__37495),
            .I(N__37489));
    LocalMux I__7686 (
            .O(N__37492),
            .I(N__37486));
    LocalMux I__7685 (
            .O(N__37489),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__7684 (
            .O(N__37486),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__7683 (
            .O(N__37481),
            .I(N__37478));
    InMux I__7682 (
            .O(N__37478),
            .I(N__37475));
    LocalMux I__7681 (
            .O(N__37475),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__7680 (
            .O(N__37472),
            .I(N__37469));
    LocalMux I__7679 (
            .O(N__37469),
            .I(N__37466));
    Odrv12 I__7678 (
            .O(N__37466),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    CascadeMux I__7677 (
            .O(N__37463),
            .I(N__37460));
    InMux I__7676 (
            .O(N__37460),
            .I(N__37457));
    LocalMux I__7675 (
            .O(N__37457),
            .I(N__37454));
    Odrv12 I__7674 (
            .O(N__37454),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    InMux I__7673 (
            .O(N__37451),
            .I(N__37448));
    LocalMux I__7672 (
            .O(N__37448),
            .I(N__37445));
    Odrv12 I__7671 (
            .O(N__37445),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ));
    CascadeMux I__7670 (
            .O(N__37442),
            .I(N__37439));
    InMux I__7669 (
            .O(N__37439),
            .I(N__37436));
    LocalMux I__7668 (
            .O(N__37436),
            .I(N__37433));
    Span4Mux_v I__7667 (
            .O(N__37433),
            .I(N__37430));
    Odrv4 I__7666 (
            .O(N__37430),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt20 ));
    InMux I__7665 (
            .O(N__37427),
            .I(N__37424));
    LocalMux I__7664 (
            .O(N__37424),
            .I(N__37421));
    Span4Mux_v I__7663 (
            .O(N__37421),
            .I(N__37418));
    Odrv4 I__7662 (
            .O(N__37418),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt22 ));
    CascadeMux I__7661 (
            .O(N__37415),
            .I(N__37412));
    InMux I__7660 (
            .O(N__37412),
            .I(N__37409));
    LocalMux I__7659 (
            .O(N__37409),
            .I(N__37406));
    Span4Mux_v I__7658 (
            .O(N__37406),
            .I(N__37403));
    Odrv4 I__7657 (
            .O(N__37403),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ));
    InMux I__7656 (
            .O(N__37400),
            .I(N__37396));
    InMux I__7655 (
            .O(N__37399),
            .I(N__37393));
    LocalMux I__7654 (
            .O(N__37396),
            .I(N__37390));
    LocalMux I__7653 (
            .O(N__37393),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__7652 (
            .O(N__37390),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__7651 (
            .O(N__37385),
            .I(N__37382));
    InMux I__7650 (
            .O(N__37382),
            .I(N__37379));
    LocalMux I__7649 (
            .O(N__37379),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    InMux I__7648 (
            .O(N__37376),
            .I(N__37373));
    LocalMux I__7647 (
            .O(N__37373),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__7646 (
            .O(N__37370),
            .I(N__37366));
    InMux I__7645 (
            .O(N__37369),
            .I(N__37363));
    LocalMux I__7644 (
            .O(N__37366),
            .I(N__37360));
    LocalMux I__7643 (
            .O(N__37363),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__7642 (
            .O(N__37360),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__7641 (
            .O(N__37355),
            .I(N__37352));
    LocalMux I__7640 (
            .O(N__37352),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__7639 (
            .O(N__37349),
            .I(N__37346));
    InMux I__7638 (
            .O(N__37346),
            .I(N__37343));
    LocalMux I__7637 (
            .O(N__37343),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__7636 (
            .O(N__37340),
            .I(N__37337));
    InMux I__7635 (
            .O(N__37337),
            .I(N__37334));
    LocalMux I__7634 (
            .O(N__37334),
            .I(N__37331));
    Odrv4 I__7633 (
            .O(N__37331),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    InMux I__7632 (
            .O(N__37328),
            .I(N__37324));
    InMux I__7631 (
            .O(N__37327),
            .I(N__37321));
    LocalMux I__7630 (
            .O(N__37324),
            .I(N__37318));
    LocalMux I__7629 (
            .O(N__37321),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__7628 (
            .O(N__37318),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__7627 (
            .O(N__37313),
            .I(N__37310));
    LocalMux I__7626 (
            .O(N__37310),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__7625 (
            .O(N__37307),
            .I(N__37303));
    InMux I__7624 (
            .O(N__37306),
            .I(N__37300));
    LocalMux I__7623 (
            .O(N__37303),
            .I(N__37297));
    LocalMux I__7622 (
            .O(N__37300),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__7621 (
            .O(N__37297),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__7620 (
            .O(N__37292),
            .I(N__37289));
    LocalMux I__7619 (
            .O(N__37289),
            .I(N__37286));
    Odrv4 I__7618 (
            .O(N__37286),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__7617 (
            .O(N__37283),
            .I(N__37280));
    InMux I__7616 (
            .O(N__37280),
            .I(N__37277));
    LocalMux I__7615 (
            .O(N__37277),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__7614 (
            .O(N__37274),
            .I(N__37271));
    LocalMux I__7613 (
            .O(N__37271),
            .I(N__37268));
    Span4Mux_h I__7612 (
            .O(N__37268),
            .I(N__37265));
    Odrv4 I__7611 (
            .O(N__37265),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    InMux I__7610 (
            .O(N__37262),
            .I(N__37259));
    LocalMux I__7609 (
            .O(N__37259),
            .I(N__37255));
    InMux I__7608 (
            .O(N__37258),
            .I(N__37252));
    Span4Mux_v I__7607 (
            .O(N__37255),
            .I(N__37249));
    LocalMux I__7606 (
            .O(N__37252),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__7605 (
            .O(N__37249),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__7604 (
            .O(N__37244),
            .I(N__37241));
    InMux I__7603 (
            .O(N__37241),
            .I(N__37238));
    LocalMux I__7602 (
            .O(N__37238),
            .I(N__37235));
    Odrv4 I__7601 (
            .O(N__37235),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__7600 (
            .O(N__37232),
            .I(N__37229));
    LocalMux I__7599 (
            .O(N__37229),
            .I(N__37226));
    Span4Mux_v I__7598 (
            .O(N__37226),
            .I(N__37223));
    Odrv4 I__7597 (
            .O(N__37223),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    InMux I__7596 (
            .O(N__37220),
            .I(N__37216));
    InMux I__7595 (
            .O(N__37219),
            .I(N__37213));
    LocalMux I__7594 (
            .O(N__37216),
            .I(N__37210));
    LocalMux I__7593 (
            .O(N__37213),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__7592 (
            .O(N__37210),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__7591 (
            .O(N__37205),
            .I(N__37202));
    InMux I__7590 (
            .O(N__37202),
            .I(N__37199));
    LocalMux I__7589 (
            .O(N__37199),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__7588 (
            .O(N__37196),
            .I(N__37193));
    LocalMux I__7587 (
            .O(N__37193),
            .I(N__37190));
    Span4Mux_v I__7586 (
            .O(N__37190),
            .I(N__37187));
    Odrv4 I__7585 (
            .O(N__37187),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    InMux I__7584 (
            .O(N__37184),
            .I(N__37181));
    LocalMux I__7583 (
            .O(N__37181),
            .I(N__37177));
    InMux I__7582 (
            .O(N__37180),
            .I(N__37174));
    Span4Mux_v I__7581 (
            .O(N__37177),
            .I(N__37171));
    LocalMux I__7580 (
            .O(N__37174),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__7579 (
            .O(N__37171),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__7578 (
            .O(N__37166),
            .I(N__37163));
    InMux I__7577 (
            .O(N__37163),
            .I(N__37160));
    LocalMux I__7576 (
            .O(N__37160),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    InMux I__7575 (
            .O(N__37157),
            .I(N__37153));
    InMux I__7574 (
            .O(N__37156),
            .I(N__37149));
    LocalMux I__7573 (
            .O(N__37153),
            .I(N__37146));
    InMux I__7572 (
            .O(N__37152),
            .I(N__37143));
    LocalMux I__7571 (
            .O(N__37149),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    Odrv4 I__7570 (
            .O(N__37146),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    LocalMux I__7569 (
            .O(N__37143),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    CascadeMux I__7568 (
            .O(N__37136),
            .I(N__37133));
    InMux I__7567 (
            .O(N__37133),
            .I(N__37130));
    LocalMux I__7566 (
            .O(N__37130),
            .I(N__37127));
    Odrv12 I__7565 (
            .O(N__37127),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__7564 (
            .O(N__37124),
            .I(N__37121));
    InMux I__7563 (
            .O(N__37121),
            .I(N__37118));
    LocalMux I__7562 (
            .O(N__37118),
            .I(N__37113));
    InMux I__7561 (
            .O(N__37117),
            .I(N__37110));
    InMux I__7560 (
            .O(N__37116),
            .I(N__37107));
    Span4Mux_h I__7559 (
            .O(N__37113),
            .I(N__37104));
    LocalMux I__7558 (
            .O(N__37110),
            .I(N__37101));
    LocalMux I__7557 (
            .O(N__37107),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__7556 (
            .O(N__37104),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__7555 (
            .O(N__37101),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__7554 (
            .O(N__37094),
            .I(N__37091));
    LocalMux I__7553 (
            .O(N__37091),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__7552 (
            .O(N__37088),
            .I(N__37084));
    InMux I__7551 (
            .O(N__37087),
            .I(N__37081));
    LocalMux I__7550 (
            .O(N__37084),
            .I(N__37078));
    LocalMux I__7549 (
            .O(N__37081),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__7548 (
            .O(N__37078),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__7547 (
            .O(N__37073),
            .I(N__37070));
    InMux I__7546 (
            .O(N__37070),
            .I(N__37067));
    LocalMux I__7545 (
            .O(N__37067),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    InMux I__7544 (
            .O(N__37064),
            .I(N__37061));
    LocalMux I__7543 (
            .O(N__37061),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    InMux I__7542 (
            .O(N__37058),
            .I(N__37055));
    LocalMux I__7541 (
            .O(N__37055),
            .I(N__37051));
    InMux I__7540 (
            .O(N__37054),
            .I(N__37048));
    Span4Mux_v I__7539 (
            .O(N__37051),
            .I(N__37045));
    LocalMux I__7538 (
            .O(N__37048),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__7537 (
            .O(N__37045),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__7536 (
            .O(N__37040),
            .I(N__37037));
    InMux I__7535 (
            .O(N__37037),
            .I(N__37034));
    LocalMux I__7534 (
            .O(N__37034),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__7533 (
            .O(N__37031),
            .I(N__37028));
    LocalMux I__7532 (
            .O(N__37028),
            .I(N__37024));
    InMux I__7531 (
            .O(N__37027),
            .I(N__37021));
    Span4Mux_v I__7530 (
            .O(N__37024),
            .I(N__37018));
    LocalMux I__7529 (
            .O(N__37021),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__7528 (
            .O(N__37018),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__7527 (
            .O(N__37013),
            .I(N__37010));
    LocalMux I__7526 (
            .O(N__37010),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__7525 (
            .O(N__37007),
            .I(N__37004));
    InMux I__7524 (
            .O(N__37004),
            .I(N__37001));
    LocalMux I__7523 (
            .O(N__37001),
            .I(N__36998));
    Odrv4 I__7522 (
            .O(N__36998),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__7521 (
            .O(N__36995),
            .I(N__36992));
    InMux I__7520 (
            .O(N__36992),
            .I(N__36988));
    InMux I__7519 (
            .O(N__36991),
            .I(N__36984));
    LocalMux I__7518 (
            .O(N__36988),
            .I(N__36981));
    InMux I__7517 (
            .O(N__36987),
            .I(N__36978));
    LocalMux I__7516 (
            .O(N__36984),
            .I(N__36975));
    Span4Mux_h I__7515 (
            .O(N__36981),
            .I(N__36972));
    LocalMux I__7514 (
            .O(N__36978),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    Odrv4 I__7513 (
            .O(N__36975),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    Odrv4 I__7512 (
            .O(N__36972),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    CascadeMux I__7511 (
            .O(N__36965),
            .I(N__36961));
    InMux I__7510 (
            .O(N__36964),
            .I(N__36955));
    InMux I__7509 (
            .O(N__36961),
            .I(N__36955));
    InMux I__7508 (
            .O(N__36960),
            .I(N__36952));
    LocalMux I__7507 (
            .O(N__36955),
            .I(N__36949));
    LocalMux I__7506 (
            .O(N__36952),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__7505 (
            .O(N__36949),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    CascadeMux I__7504 (
            .O(N__36944),
            .I(N__36941));
    InMux I__7503 (
            .O(N__36941),
            .I(N__36937));
    InMux I__7502 (
            .O(N__36940),
            .I(N__36934));
    LocalMux I__7501 (
            .O(N__36937),
            .I(N__36928));
    LocalMux I__7500 (
            .O(N__36934),
            .I(N__36928));
    InMux I__7499 (
            .O(N__36933),
            .I(N__36925));
    Span4Mux_v I__7498 (
            .O(N__36928),
            .I(N__36922));
    LocalMux I__7497 (
            .O(N__36925),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__7496 (
            .O(N__36922),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__7495 (
            .O(N__36917),
            .I(N__36913));
    InMux I__7494 (
            .O(N__36916),
            .I(N__36910));
    LocalMux I__7493 (
            .O(N__36913),
            .I(N__36905));
    LocalMux I__7492 (
            .O(N__36910),
            .I(N__36905));
    Odrv4 I__7491 (
            .O(N__36905),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ));
    InMux I__7490 (
            .O(N__36902),
            .I(N__36896));
    InMux I__7489 (
            .O(N__36901),
            .I(N__36896));
    LocalMux I__7488 (
            .O(N__36896),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ));
    InMux I__7487 (
            .O(N__36893),
            .I(N__36889));
    InMux I__7486 (
            .O(N__36892),
            .I(N__36886));
    LocalMux I__7485 (
            .O(N__36889),
            .I(N__36880));
    LocalMux I__7484 (
            .O(N__36886),
            .I(N__36880));
    InMux I__7483 (
            .O(N__36885),
            .I(N__36877));
    Span4Mux_v I__7482 (
            .O(N__36880),
            .I(N__36874));
    LocalMux I__7481 (
            .O(N__36877),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    Odrv4 I__7480 (
            .O(N__36874),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    CascadeMux I__7479 (
            .O(N__36869),
            .I(N__36865));
    InMux I__7478 (
            .O(N__36868),
            .I(N__36860));
    InMux I__7477 (
            .O(N__36865),
            .I(N__36860));
    LocalMux I__7476 (
            .O(N__36860),
            .I(N__36857));
    Span4Mux_v I__7475 (
            .O(N__36857),
            .I(N__36854));
    Odrv4 I__7474 (
            .O(N__36854),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__7473 (
            .O(N__36851),
            .I(N__36846));
    InMux I__7472 (
            .O(N__36850),
            .I(N__36843));
    InMux I__7471 (
            .O(N__36849),
            .I(N__36838));
    InMux I__7470 (
            .O(N__36846),
            .I(N__36838));
    LocalMux I__7469 (
            .O(N__36843),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__7468 (
            .O(N__36838),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__7467 (
            .O(N__36833),
            .I(N__36828));
    InMux I__7466 (
            .O(N__36832),
            .I(N__36823));
    InMux I__7465 (
            .O(N__36831),
            .I(N__36823));
    LocalMux I__7464 (
            .O(N__36828),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__7463 (
            .O(N__36823),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__7462 (
            .O(N__36818),
            .I(N__36815));
    LocalMux I__7461 (
            .O(N__36815),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ));
    CascadeMux I__7460 (
            .O(N__36812),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ));
    InMux I__7459 (
            .O(N__36809),
            .I(N__36806));
    LocalMux I__7458 (
            .O(N__36806),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ));
    InMux I__7457 (
            .O(N__36803),
            .I(N__36800));
    LocalMux I__7456 (
            .O(N__36800),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ));
    CascadeMux I__7455 (
            .O(N__36797),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ));
    InMux I__7454 (
            .O(N__36794),
            .I(N__36791));
    LocalMux I__7453 (
            .O(N__36791),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ));
    InMux I__7452 (
            .O(N__36788),
            .I(N__36785));
    LocalMux I__7451 (
            .O(N__36785),
            .I(N__36782));
    Span4Mux_v I__7450 (
            .O(N__36782),
            .I(N__36778));
    InMux I__7449 (
            .O(N__36781),
            .I(N__36775));
    Odrv4 I__7448 (
            .O(N__36778),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    LocalMux I__7447 (
            .O(N__36775),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    CascadeMux I__7446 (
            .O(N__36770),
            .I(elapsed_time_ns_1_RNITUBN9_0_10_cascade_));
    CascadeMux I__7445 (
            .O(N__36767),
            .I(N__36764));
    InMux I__7444 (
            .O(N__36764),
            .I(N__36761));
    LocalMux I__7443 (
            .O(N__36761),
            .I(N__36758));
    Span4Mux_v I__7442 (
            .O(N__36758),
            .I(N__36755));
    Odrv4 I__7441 (
            .O(N__36755),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__7440 (
            .O(N__36752),
            .I(N__36744));
    InMux I__7439 (
            .O(N__36751),
            .I(N__36744));
    InMux I__7438 (
            .O(N__36750),
            .I(N__36741));
    InMux I__7437 (
            .O(N__36749),
            .I(N__36738));
    LocalMux I__7436 (
            .O(N__36744),
            .I(N__36733));
    LocalMux I__7435 (
            .O(N__36741),
            .I(N__36733));
    LocalMux I__7434 (
            .O(N__36738),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv4 I__7433 (
            .O(N__36733),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__7432 (
            .O(N__36728),
            .I(N__36720));
    InMux I__7431 (
            .O(N__36727),
            .I(N__36720));
    InMux I__7430 (
            .O(N__36726),
            .I(N__36717));
    InMux I__7429 (
            .O(N__36725),
            .I(N__36714));
    LocalMux I__7428 (
            .O(N__36720),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7427 (
            .O(N__36717),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7426 (
            .O(N__36714),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    CascadeMux I__7425 (
            .O(N__36707),
            .I(N__36704));
    InMux I__7424 (
            .O(N__36704),
            .I(N__36701));
    LocalMux I__7423 (
            .O(N__36701),
            .I(N__36698));
    Span4Mux_v I__7422 (
            .O(N__36698),
            .I(N__36695));
    Odrv4 I__7421 (
            .O(N__36695),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__7420 (
            .O(N__36692),
            .I(N__36689));
    LocalMux I__7419 (
            .O(N__36689),
            .I(N__36686));
    Span4Mux_v I__7418 (
            .O(N__36686),
            .I(N__36681));
    InMux I__7417 (
            .O(N__36685),
            .I(N__36678));
    InMux I__7416 (
            .O(N__36684),
            .I(N__36675));
    Span4Mux_v I__7415 (
            .O(N__36681),
            .I(N__36670));
    LocalMux I__7414 (
            .O(N__36678),
            .I(N__36670));
    LocalMux I__7413 (
            .O(N__36675),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv4 I__7412 (
            .O(N__36670),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__7411 (
            .O(N__36665),
            .I(N__36662));
    LocalMux I__7410 (
            .O(N__36662),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__7409 (
            .O(N__36659),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__7408 (
            .O(N__36656),
            .I(N__36653));
    LocalMux I__7407 (
            .O(N__36653),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__7406 (
            .O(N__36650),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__7405 (
            .O(N__36647),
            .I(N__36644));
    LocalMux I__7404 (
            .O(N__36644),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__7403 (
            .O(N__36641),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__7402 (
            .O(N__36638),
            .I(N__36635));
    LocalMux I__7401 (
            .O(N__36635),
            .I(N__36632));
    Odrv4 I__7400 (
            .O(N__36632),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__7399 (
            .O(N__36629),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__7398 (
            .O(N__36626),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__7397 (
            .O(N__36623),
            .I(N__36620));
    LocalMux I__7396 (
            .O(N__36620),
            .I(N__36617));
    Span4Mux_h I__7395 (
            .O(N__36617),
            .I(N__36614));
    Odrv4 I__7394 (
            .O(N__36614),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__7393 (
            .O(N__36611),
            .I(N__36608));
    LocalMux I__7392 (
            .O(N__36608),
            .I(N__36605));
    Span4Mux_v I__7391 (
            .O(N__36605),
            .I(N__36602));
    Odrv4 I__7390 (
            .O(N__36602),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ));
    InMux I__7389 (
            .O(N__36599),
            .I(N__36596));
    LocalMux I__7388 (
            .O(N__36596),
            .I(N__36593));
    Span4Mux_v I__7387 (
            .O(N__36593),
            .I(N__36590));
    Odrv4 I__7386 (
            .O(N__36590),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ));
    InMux I__7385 (
            .O(N__36587),
            .I(N__36584));
    LocalMux I__7384 (
            .O(N__36584),
            .I(\current_shift_inst.un38_control_input_0_s1_18 ));
    InMux I__7383 (
            .O(N__36581),
            .I(\current_shift_inst.un38_control_input_cry_17_s1 ));
    InMux I__7382 (
            .O(N__36578),
            .I(N__36575));
    LocalMux I__7381 (
            .O(N__36575),
            .I(\current_shift_inst.un38_control_input_0_s1_19 ));
    InMux I__7380 (
            .O(N__36572),
            .I(\current_shift_inst.un38_control_input_cry_18_s1 ));
    InMux I__7379 (
            .O(N__36569),
            .I(N__36566));
    LocalMux I__7378 (
            .O(N__36566),
            .I(N__36563));
    Span4Mux_h I__7377 (
            .O(N__36563),
            .I(N__36560));
    Odrv4 I__7376 (
            .O(N__36560),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__7375 (
            .O(N__36557),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__7374 (
            .O(N__36554),
            .I(N__36551));
    LocalMux I__7373 (
            .O(N__36551),
            .I(N__36548));
    Span4Mux_h I__7372 (
            .O(N__36548),
            .I(N__36545));
    Odrv4 I__7371 (
            .O(N__36545),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__7370 (
            .O(N__36542),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    CascadeMux I__7369 (
            .O(N__36539),
            .I(N__36536));
    InMux I__7368 (
            .O(N__36536),
            .I(N__36533));
    LocalMux I__7367 (
            .O(N__36533),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__7366 (
            .O(N__36530),
            .I(N__36527));
    LocalMux I__7365 (
            .O(N__36527),
            .I(N__36524));
    Odrv12 I__7364 (
            .O(N__36524),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__7363 (
            .O(N__36521),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__7362 (
            .O(N__36518),
            .I(N__36515));
    LocalMux I__7361 (
            .O(N__36515),
            .I(N__36512));
    Odrv4 I__7360 (
            .O(N__36512),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__7359 (
            .O(N__36509),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__7358 (
            .O(N__36506),
            .I(N__36503));
    LocalMux I__7357 (
            .O(N__36503),
            .I(N__36500));
    Span4Mux_h I__7356 (
            .O(N__36500),
            .I(N__36497));
    Odrv4 I__7355 (
            .O(N__36497),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__7354 (
            .O(N__36494),
            .I(bfn_14_18_0_));
    InMux I__7353 (
            .O(N__36491),
            .I(N__36488));
    LocalMux I__7352 (
            .O(N__36488),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__7351 (
            .O(N__36485),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    InMux I__7350 (
            .O(N__36482),
            .I(N__36479));
    LocalMux I__7349 (
            .O(N__36479),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__7348 (
            .O(N__36476),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__7347 (
            .O(N__36473),
            .I(N__36470));
    LocalMux I__7346 (
            .O(N__36470),
            .I(\current_shift_inst.un38_control_input_0_s1_10 ));
    InMux I__7345 (
            .O(N__36467),
            .I(\current_shift_inst.un38_control_input_cry_9_s1 ));
    InMux I__7344 (
            .O(N__36464),
            .I(N__36461));
    LocalMux I__7343 (
            .O(N__36461),
            .I(N__36458));
    Span4Mux_v I__7342 (
            .O(N__36458),
            .I(N__36455));
    Odrv4 I__7341 (
            .O(N__36455),
            .I(\current_shift_inst.un38_control_input_0_s1_11 ));
    InMux I__7340 (
            .O(N__36452),
            .I(\current_shift_inst.un38_control_input_cry_10_s1 ));
    InMux I__7339 (
            .O(N__36449),
            .I(N__36446));
    LocalMux I__7338 (
            .O(N__36446),
            .I(N__36443));
    Span4Mux_h I__7337 (
            .O(N__36443),
            .I(N__36440));
    Odrv4 I__7336 (
            .O(N__36440),
            .I(\current_shift_inst.un38_control_input_0_s1_12 ));
    InMux I__7335 (
            .O(N__36437),
            .I(\current_shift_inst.un38_control_input_cry_11_s1 ));
    InMux I__7334 (
            .O(N__36434),
            .I(N__36431));
    LocalMux I__7333 (
            .O(N__36431),
            .I(N__36428));
    Odrv12 I__7332 (
            .O(N__36428),
            .I(\current_shift_inst.un38_control_input_0_s1_13 ));
    InMux I__7331 (
            .O(N__36425),
            .I(\current_shift_inst.un38_control_input_cry_12_s1 ));
    InMux I__7330 (
            .O(N__36422),
            .I(N__36419));
    LocalMux I__7329 (
            .O(N__36419),
            .I(\current_shift_inst.un38_control_input_0_s1_14 ));
    InMux I__7328 (
            .O(N__36416),
            .I(\current_shift_inst.un38_control_input_cry_13_s1 ));
    InMux I__7327 (
            .O(N__36413),
            .I(N__36410));
    LocalMux I__7326 (
            .O(N__36410),
            .I(\current_shift_inst.un38_control_input_0_s1_15 ));
    InMux I__7325 (
            .O(N__36407),
            .I(\current_shift_inst.un38_control_input_cry_14_s1 ));
    InMux I__7324 (
            .O(N__36404),
            .I(N__36401));
    LocalMux I__7323 (
            .O(N__36401),
            .I(\current_shift_inst.un38_control_input_0_s1_16 ));
    InMux I__7322 (
            .O(N__36398),
            .I(bfn_14_17_0_));
    InMux I__7321 (
            .O(N__36395),
            .I(N__36392));
    LocalMux I__7320 (
            .O(N__36392),
            .I(\current_shift_inst.un38_control_input_0_s1_17 ));
    InMux I__7319 (
            .O(N__36389),
            .I(\current_shift_inst.un38_control_input_cry_16_s1 ));
    InMux I__7318 (
            .O(N__36386),
            .I(N__36383));
    LocalMux I__7317 (
            .O(N__36383),
            .I(N__36380));
    Odrv12 I__7316 (
            .O(N__36380),
            .I(\current_shift_inst.un38_control_input_0_s1_3 ));
    InMux I__7315 (
            .O(N__36377),
            .I(\current_shift_inst.un38_control_input_cry_2_s1 ));
    InMux I__7314 (
            .O(N__36374),
            .I(N__36371));
    LocalMux I__7313 (
            .O(N__36371),
            .I(N__36368));
    Odrv4 I__7312 (
            .O(N__36368),
            .I(\current_shift_inst.un38_control_input_0_s1_4 ));
    InMux I__7311 (
            .O(N__36365),
            .I(\current_shift_inst.un38_control_input_cry_3_s1 ));
    InMux I__7310 (
            .O(N__36362),
            .I(N__36359));
    LocalMux I__7309 (
            .O(N__36359),
            .I(N__36356));
    Odrv4 I__7308 (
            .O(N__36356),
            .I(\current_shift_inst.un38_control_input_0_s1_5 ));
    InMux I__7307 (
            .O(N__36353),
            .I(\current_shift_inst.un38_control_input_cry_4_s1 ));
    CascadeMux I__7306 (
            .O(N__36350),
            .I(N__36347));
    InMux I__7305 (
            .O(N__36347),
            .I(N__36344));
    LocalMux I__7304 (
            .O(N__36344),
            .I(N__36341));
    Span4Mux_h I__7303 (
            .O(N__36341),
            .I(N__36338));
    Odrv4 I__7302 (
            .O(N__36338),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ));
    InMux I__7301 (
            .O(N__36335),
            .I(N__36332));
    LocalMux I__7300 (
            .O(N__36332),
            .I(N__36329));
    Odrv12 I__7299 (
            .O(N__36329),
            .I(\current_shift_inst.un38_control_input_0_s1_6 ));
    InMux I__7298 (
            .O(N__36326),
            .I(\current_shift_inst.un38_control_input_cry_5_s1 ));
    InMux I__7297 (
            .O(N__36323),
            .I(N__36320));
    LocalMux I__7296 (
            .O(N__36320),
            .I(N__36317));
    Odrv4 I__7295 (
            .O(N__36317),
            .I(\current_shift_inst.un38_control_input_0_s1_7 ));
    InMux I__7294 (
            .O(N__36314),
            .I(\current_shift_inst.un38_control_input_cry_6_s1 ));
    InMux I__7293 (
            .O(N__36311),
            .I(N__36308));
    LocalMux I__7292 (
            .O(N__36308),
            .I(N__36305));
    Span4Mux_v I__7291 (
            .O(N__36305),
            .I(N__36302));
    Odrv4 I__7290 (
            .O(N__36302),
            .I(\current_shift_inst.un38_control_input_0_s1_8 ));
    InMux I__7289 (
            .O(N__36299),
            .I(bfn_14_16_0_));
    InMux I__7288 (
            .O(N__36296),
            .I(N__36293));
    LocalMux I__7287 (
            .O(N__36293),
            .I(N__36290));
    Span4Mux_v I__7286 (
            .O(N__36290),
            .I(N__36287));
    Span4Mux_h I__7285 (
            .O(N__36287),
            .I(N__36284));
    Odrv4 I__7284 (
            .O(N__36284),
            .I(\current_shift_inst.un38_control_input_0_s1_9 ));
    InMux I__7283 (
            .O(N__36281),
            .I(\current_shift_inst.un38_control_input_cry_8_s1 ));
    InMux I__7282 (
            .O(N__36278),
            .I(N__36273));
    InMux I__7281 (
            .O(N__36277),
            .I(N__36268));
    InMux I__7280 (
            .O(N__36276),
            .I(N__36268));
    LocalMux I__7279 (
            .O(N__36273),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__7278 (
            .O(N__36268),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__7277 (
            .O(N__36263),
            .I(bfn_14_14_0_));
    InMux I__7276 (
            .O(N__36260),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__7275 (
            .O(N__36257),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__7274 (
            .O(N__36254),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__7273 (
            .O(N__36251),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__7272 (
            .O(N__36248),
            .I(N__36243));
    InMux I__7271 (
            .O(N__36247),
            .I(N__36238));
    InMux I__7270 (
            .O(N__36246),
            .I(N__36238));
    LocalMux I__7269 (
            .O(N__36243),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    LocalMux I__7268 (
            .O(N__36238),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__7267 (
            .O(N__36233),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    IoInMux I__7266 (
            .O(N__36230),
            .I(N__36213));
    InMux I__7265 (
            .O(N__36229),
            .I(N__36206));
    InMux I__7264 (
            .O(N__36228),
            .I(N__36206));
    InMux I__7263 (
            .O(N__36227),
            .I(N__36206));
    InMux I__7262 (
            .O(N__36226),
            .I(N__36197));
    InMux I__7261 (
            .O(N__36225),
            .I(N__36197));
    InMux I__7260 (
            .O(N__36224),
            .I(N__36197));
    InMux I__7259 (
            .O(N__36223),
            .I(N__36197));
    InMux I__7258 (
            .O(N__36222),
            .I(N__36186));
    InMux I__7257 (
            .O(N__36221),
            .I(N__36186));
    InMux I__7256 (
            .O(N__36220),
            .I(N__36186));
    InMux I__7255 (
            .O(N__36219),
            .I(N__36177));
    InMux I__7254 (
            .O(N__36218),
            .I(N__36177));
    InMux I__7253 (
            .O(N__36217),
            .I(N__36177));
    InMux I__7252 (
            .O(N__36216),
            .I(N__36177));
    LocalMux I__7251 (
            .O(N__36213),
            .I(N__36170));
    LocalMux I__7250 (
            .O(N__36206),
            .I(N__36158));
    LocalMux I__7249 (
            .O(N__36197),
            .I(N__36155));
    InMux I__7248 (
            .O(N__36196),
            .I(N__36146));
    InMux I__7247 (
            .O(N__36195),
            .I(N__36146));
    InMux I__7246 (
            .O(N__36194),
            .I(N__36146));
    InMux I__7245 (
            .O(N__36193),
            .I(N__36146));
    LocalMux I__7244 (
            .O(N__36186),
            .I(N__36141));
    LocalMux I__7243 (
            .O(N__36177),
            .I(N__36141));
    InMux I__7242 (
            .O(N__36176),
            .I(N__36132));
    InMux I__7241 (
            .O(N__36175),
            .I(N__36132));
    InMux I__7240 (
            .O(N__36174),
            .I(N__36132));
    InMux I__7239 (
            .O(N__36173),
            .I(N__36132));
    IoSpan4Mux I__7238 (
            .O(N__36170),
            .I(N__36129));
    InMux I__7237 (
            .O(N__36169),
            .I(N__36126));
    InMux I__7236 (
            .O(N__36168),
            .I(N__36117));
    InMux I__7235 (
            .O(N__36167),
            .I(N__36117));
    InMux I__7234 (
            .O(N__36166),
            .I(N__36117));
    InMux I__7233 (
            .O(N__36165),
            .I(N__36117));
    InMux I__7232 (
            .O(N__36164),
            .I(N__36108));
    InMux I__7231 (
            .O(N__36163),
            .I(N__36108));
    InMux I__7230 (
            .O(N__36162),
            .I(N__36108));
    InMux I__7229 (
            .O(N__36161),
            .I(N__36108));
    Span4Mux_v I__7228 (
            .O(N__36158),
            .I(N__36097));
    Span4Mux_v I__7227 (
            .O(N__36155),
            .I(N__36097));
    LocalMux I__7226 (
            .O(N__36146),
            .I(N__36097));
    Span4Mux_v I__7225 (
            .O(N__36141),
            .I(N__36097));
    LocalMux I__7224 (
            .O(N__36132),
            .I(N__36097));
    Span4Mux_s1_v I__7223 (
            .O(N__36129),
            .I(N__36094));
    LocalMux I__7222 (
            .O(N__36126),
            .I(N__36087));
    LocalMux I__7221 (
            .O(N__36117),
            .I(N__36087));
    LocalMux I__7220 (
            .O(N__36108),
            .I(N__36087));
    Span4Mux_h I__7219 (
            .O(N__36097),
            .I(N__36084));
    Sp12to4 I__7218 (
            .O(N__36094),
            .I(N__36081));
    Span12Mux_h I__7217 (
            .O(N__36087),
            .I(N__36078));
    Span4Mux_h I__7216 (
            .O(N__36084),
            .I(N__36075));
    Span12Mux_s9_v I__7215 (
            .O(N__36081),
            .I(N__36072));
    Odrv12 I__7214 (
            .O(N__36078),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__7213 (
            .O(N__36075),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv12 I__7212 (
            .O(N__36072),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__7211 (
            .O(N__36065),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    CascadeMux I__7210 (
            .O(N__36062),
            .I(N__36058));
    InMux I__7209 (
            .O(N__36061),
            .I(N__36054));
    InMux I__7208 (
            .O(N__36058),
            .I(N__36049));
    InMux I__7207 (
            .O(N__36057),
            .I(N__36049));
    LocalMux I__7206 (
            .O(N__36054),
            .I(N__36044));
    LocalMux I__7205 (
            .O(N__36049),
            .I(N__36044));
    Odrv4 I__7204 (
            .O(N__36044),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__7203 (
            .O(N__36041),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__7202 (
            .O(N__36038),
            .I(bfn_14_13_0_));
    InMux I__7201 (
            .O(N__36035),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__7200 (
            .O(N__36032),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__7199 (
            .O(N__36029),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__7198 (
            .O(N__36026),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__7197 (
            .O(N__36023),
            .I(N__36018));
    InMux I__7196 (
            .O(N__36022),
            .I(N__36015));
    InMux I__7195 (
            .O(N__36021),
            .I(N__36010));
    InMux I__7194 (
            .O(N__36018),
            .I(N__36010));
    LocalMux I__7193 (
            .O(N__36015),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    LocalMux I__7192 (
            .O(N__36010),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__7191 (
            .O(N__36005),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    CascadeMux I__7190 (
            .O(N__36002),
            .I(N__35997));
    InMux I__7189 (
            .O(N__36001),
            .I(N__35994));
    InMux I__7188 (
            .O(N__36000),
            .I(N__35989));
    InMux I__7187 (
            .O(N__35997),
            .I(N__35989));
    LocalMux I__7186 (
            .O(N__35994),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    LocalMux I__7185 (
            .O(N__35989),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__7184 (
            .O(N__35984),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    CascadeMux I__7183 (
            .O(N__35981),
            .I(N__35977));
    InMux I__7182 (
            .O(N__35980),
            .I(N__35973));
    InMux I__7181 (
            .O(N__35977),
            .I(N__35968));
    InMux I__7180 (
            .O(N__35976),
            .I(N__35968));
    LocalMux I__7179 (
            .O(N__35973),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    LocalMux I__7178 (
            .O(N__35968),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__7177 (
            .O(N__35963),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__7176 (
            .O(N__35960),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__7175 (
            .O(N__35957),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__7174 (
            .O(N__35954),
            .I(bfn_14_12_0_));
    InMux I__7173 (
            .O(N__35951),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__7172 (
            .O(N__35948),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__7171 (
            .O(N__35945),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__7170 (
            .O(N__35942),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__7169 (
            .O(N__35939),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__7168 (
            .O(N__35936),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__7167 (
            .O(N__35933),
            .I(N__35929));
    InMux I__7166 (
            .O(N__35932),
            .I(N__35925));
    LocalMux I__7165 (
            .O(N__35929),
            .I(N__35922));
    InMux I__7164 (
            .O(N__35928),
            .I(N__35919));
    LocalMux I__7163 (
            .O(N__35925),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    Odrv4 I__7162 (
            .O(N__35922),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    LocalMux I__7161 (
            .O(N__35919),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    InMux I__7160 (
            .O(N__35912),
            .I(N__35909));
    LocalMux I__7159 (
            .O(N__35909),
            .I(N__35906));
    Span4Mux_h I__7158 (
            .O(N__35906),
            .I(N__35903));
    Odrv4 I__7157 (
            .O(N__35903),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    InMux I__7156 (
            .O(N__35900),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__7155 (
            .O(N__35897),
            .I(N__35894));
    InMux I__7154 (
            .O(N__35894),
            .I(N__35891));
    LocalMux I__7153 (
            .O(N__35891),
            .I(N__35888));
    Span4Mux_h I__7152 (
            .O(N__35888),
            .I(N__35885));
    Odrv4 I__7151 (
            .O(N__35885),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ));
    InMux I__7150 (
            .O(N__35882),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__7149 (
            .O(N__35879),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__7148 (
            .O(N__35876),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__7147 (
            .O(N__35873),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    IoInMux I__7146 (
            .O(N__35870),
            .I(N__35867));
    LocalMux I__7145 (
            .O(N__35867),
            .I(s2_phy_c));
    InMux I__7144 (
            .O(N__35864),
            .I(N__35861));
    LocalMux I__7143 (
            .O(N__35861),
            .I(N__35857));
    InMux I__7142 (
            .O(N__35860),
            .I(N__35854));
    Span4Mux_v I__7141 (
            .O(N__35857),
            .I(N__35847));
    LocalMux I__7140 (
            .O(N__35854),
            .I(N__35847));
    InMux I__7139 (
            .O(N__35853),
            .I(N__35844));
    InMux I__7138 (
            .O(N__35852),
            .I(N__35841));
    Span4Mux_v I__7137 (
            .O(N__35847),
            .I(N__35838));
    LocalMux I__7136 (
            .O(N__35844),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__7135 (
            .O(N__35841),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__7134 (
            .O(N__35838),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__7133 (
            .O(N__35831),
            .I(N__35828));
    LocalMux I__7132 (
            .O(N__35828),
            .I(N__35823));
    InMux I__7131 (
            .O(N__35827),
            .I(N__35818));
    InMux I__7130 (
            .O(N__35826),
            .I(N__35818));
    Span4Mux_h I__7129 (
            .O(N__35823),
            .I(N__35812));
    LocalMux I__7128 (
            .O(N__35818),
            .I(N__35812));
    InMux I__7127 (
            .O(N__35817),
            .I(N__35809));
    Span4Mux_v I__7126 (
            .O(N__35812),
            .I(N__35806));
    LocalMux I__7125 (
            .O(N__35809),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__7124 (
            .O(N__35806),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__7123 (
            .O(N__35801),
            .I(N__35798));
    LocalMux I__7122 (
            .O(N__35798),
            .I(N__35793));
    InMux I__7121 (
            .O(N__35797),
            .I(N__35790));
    InMux I__7120 (
            .O(N__35796),
            .I(N__35787));
    Span4Mux_v I__7119 (
            .O(N__35793),
            .I(N__35782));
    LocalMux I__7118 (
            .O(N__35790),
            .I(N__35782));
    LocalMux I__7117 (
            .O(N__35787),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__7116 (
            .O(N__35782),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__7115 (
            .O(N__35777),
            .I(N__35774));
    LocalMux I__7114 (
            .O(N__35774),
            .I(N__35770));
    InMux I__7113 (
            .O(N__35773),
            .I(N__35766));
    Span4Mux_v I__7112 (
            .O(N__35770),
            .I(N__35763));
    InMux I__7111 (
            .O(N__35769),
            .I(N__35760));
    LocalMux I__7110 (
            .O(N__35766),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    Odrv4 I__7109 (
            .O(N__35763),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    LocalMux I__7108 (
            .O(N__35760),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    InMux I__7107 (
            .O(N__35753),
            .I(N__35750));
    LocalMux I__7106 (
            .O(N__35750),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__7105 (
            .O(N__35747),
            .I(N__35744));
    LocalMux I__7104 (
            .O(N__35744),
            .I(N__35741));
    Span4Mux_v I__7103 (
            .O(N__35741),
            .I(N__35738));
    Odrv4 I__7102 (
            .O(N__35738),
            .I(\current_shift_inst.control_input_axb_21 ));
    InMux I__7101 (
            .O(N__35735),
            .I(N__35732));
    LocalMux I__7100 (
            .O(N__35732),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__7099 (
            .O(N__35729),
            .I(N__35726));
    LocalMux I__7098 (
            .O(N__35726),
            .I(N__35723));
    Span4Mux_h I__7097 (
            .O(N__35723),
            .I(N__35720));
    Odrv4 I__7096 (
            .O(N__35720),
            .I(\current_shift_inst.control_input_axb_22 ));
    CascadeMux I__7095 (
            .O(N__35717),
            .I(N__35714));
    InMux I__7094 (
            .O(N__35714),
            .I(N__35711));
    LocalMux I__7093 (
            .O(N__35711),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__7092 (
            .O(N__35708),
            .I(N__35705));
    LocalMux I__7091 (
            .O(N__35705),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__7090 (
            .O(N__35702),
            .I(N__35699));
    LocalMux I__7089 (
            .O(N__35699),
            .I(N__35696));
    Span4Mux_h I__7088 (
            .O(N__35696),
            .I(N__35693));
    Odrv4 I__7087 (
            .O(N__35693),
            .I(\current_shift_inst.control_input_axb_23 ));
    CascadeMux I__7086 (
            .O(N__35690),
            .I(N__35687));
    InMux I__7085 (
            .O(N__35687),
            .I(N__35684));
    LocalMux I__7084 (
            .O(N__35684),
            .I(N__35681));
    Span4Mux_h I__7083 (
            .O(N__35681),
            .I(N__35677));
    InMux I__7082 (
            .O(N__35680),
            .I(N__35673));
    Sp12to4 I__7081 (
            .O(N__35677),
            .I(N__35670));
    InMux I__7080 (
            .O(N__35676),
            .I(N__35667));
    LocalMux I__7079 (
            .O(N__35673),
            .I(N__35660));
    Span12Mux_v I__7078 (
            .O(N__35670),
            .I(N__35660));
    LocalMux I__7077 (
            .O(N__35667),
            .I(N__35660));
    Span12Mux_v I__7076 (
            .O(N__35660),
            .I(N__35657));
    Odrv12 I__7075 (
            .O(N__35657),
            .I(il_max_comp1_D2));
    IoInMux I__7074 (
            .O(N__35654),
            .I(N__35651));
    LocalMux I__7073 (
            .O(N__35651),
            .I(N__35648));
    Span4Mux_s3_v I__7072 (
            .O(N__35648),
            .I(N__35645));
    Sp12to4 I__7071 (
            .O(N__35645),
            .I(N__35642));
    Span12Mux_h I__7070 (
            .O(N__35642),
            .I(N__35638));
    InMux I__7069 (
            .O(N__35641),
            .I(N__35635));
    Odrv12 I__7068 (
            .O(N__35638),
            .I(T01_c));
    LocalMux I__7067 (
            .O(N__35635),
            .I(T01_c));
    CascadeMux I__7066 (
            .O(N__35630),
            .I(N__35625));
    InMux I__7065 (
            .O(N__35629),
            .I(N__35618));
    InMux I__7064 (
            .O(N__35628),
            .I(N__35618));
    InMux I__7063 (
            .O(N__35625),
            .I(N__35615));
    InMux I__7062 (
            .O(N__35624),
            .I(N__35610));
    InMux I__7061 (
            .O(N__35623),
            .I(N__35610));
    LocalMux I__7060 (
            .O(N__35618),
            .I(N__35603));
    LocalMux I__7059 (
            .O(N__35615),
            .I(N__35603));
    LocalMux I__7058 (
            .O(N__35610),
            .I(N__35603));
    Span4Mux_v I__7057 (
            .O(N__35603),
            .I(N__35598));
    InMux I__7056 (
            .O(N__35602),
            .I(N__35593));
    InMux I__7055 (
            .O(N__35601),
            .I(N__35593));
    Odrv4 I__7054 (
            .O(N__35598),
            .I(state_3));
    LocalMux I__7053 (
            .O(N__35593),
            .I(state_3));
    IoInMux I__7052 (
            .O(N__35588),
            .I(N__35585));
    LocalMux I__7051 (
            .O(N__35585),
            .I(N__35582));
    Span4Mux_s2_v I__7050 (
            .O(N__35582),
            .I(N__35579));
    Span4Mux_h I__7049 (
            .O(N__35579),
            .I(N__35576));
    Span4Mux_v I__7048 (
            .O(N__35576),
            .I(N__35571));
    InMux I__7047 (
            .O(N__35575),
            .I(N__35568));
    InMux I__7046 (
            .O(N__35574),
            .I(N__35565));
    Odrv4 I__7045 (
            .O(N__35571),
            .I(s1_phy_c));
    LocalMux I__7044 (
            .O(N__35568),
            .I(s1_phy_c));
    LocalMux I__7043 (
            .O(N__35565),
            .I(s1_phy_c));
    IoInMux I__7042 (
            .O(N__35558),
            .I(N__35555));
    LocalMux I__7041 (
            .O(N__35555),
            .I(N__35552));
    Span12Mux_s0_v I__7040 (
            .O(N__35552),
            .I(N__35549));
    Odrv12 I__7039 (
            .O(N__35549),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    InMux I__7038 (
            .O(N__35546),
            .I(N__35543));
    LocalMux I__7037 (
            .O(N__35543),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ));
    InMux I__7036 (
            .O(N__35540),
            .I(N__35537));
    LocalMux I__7035 (
            .O(N__35537),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__7034 (
            .O(N__35534),
            .I(N__35531));
    LocalMux I__7033 (
            .O(N__35531),
            .I(N__35528));
    Odrv4 I__7032 (
            .O(N__35528),
            .I(\current_shift_inst.control_input_axb_24 ));
    InMux I__7031 (
            .O(N__35525),
            .I(N__35522));
    LocalMux I__7030 (
            .O(N__35522),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    CascadeMux I__7029 (
            .O(N__35519),
            .I(N__35516));
    InMux I__7028 (
            .O(N__35516),
            .I(N__35513));
    LocalMux I__7027 (
            .O(N__35513),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ));
    CascadeMux I__7026 (
            .O(N__35510),
            .I(N__35507));
    InMux I__7025 (
            .O(N__35507),
            .I(N__35504));
    LocalMux I__7024 (
            .O(N__35504),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ));
    InMux I__7023 (
            .O(N__35501),
            .I(N__35498));
    LocalMux I__7022 (
            .O(N__35498),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    CascadeMux I__7021 (
            .O(N__35495),
            .I(N__35492));
    InMux I__7020 (
            .O(N__35492),
            .I(N__35489));
    LocalMux I__7019 (
            .O(N__35489),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__7018 (
            .O(N__35486),
            .I(N__35483));
    LocalMux I__7017 (
            .O(N__35483),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__7016 (
            .O(N__35480),
            .I(N__35477));
    LocalMux I__7015 (
            .O(N__35477),
            .I(N__35474));
    Span4Mux_v I__7014 (
            .O(N__35474),
            .I(N__35471));
    Odrv4 I__7013 (
            .O(N__35471),
            .I(\current_shift_inst.control_input_axb_26 ));
    InMux I__7012 (
            .O(N__35468),
            .I(N__35465));
    LocalMux I__7011 (
            .O(N__35465),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__7010 (
            .O(N__35462),
            .I(N__35459));
    LocalMux I__7009 (
            .O(N__35459),
            .I(N__35456));
    Span4Mux_v I__7008 (
            .O(N__35456),
            .I(N__35453));
    Odrv4 I__7007 (
            .O(N__35453),
            .I(\current_shift_inst.control_input_axb_20 ));
    CascadeMux I__7006 (
            .O(N__35450),
            .I(N__35447));
    InMux I__7005 (
            .O(N__35447),
            .I(N__35444));
    LocalMux I__7004 (
            .O(N__35444),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ));
    CascadeMux I__7003 (
            .O(N__35441),
            .I(N__35438));
    InMux I__7002 (
            .O(N__35438),
            .I(N__35435));
    LocalMux I__7001 (
            .O(N__35435),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    CascadeMux I__7000 (
            .O(N__35432),
            .I(N__35429));
    InMux I__6999 (
            .O(N__35429),
            .I(N__35426));
    LocalMux I__6998 (
            .O(N__35426),
            .I(N__35423));
    Odrv12 I__6997 (
            .O(N__35423),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ));
    CascadeMux I__6996 (
            .O(N__35420),
            .I(N__35417));
    InMux I__6995 (
            .O(N__35417),
            .I(N__35414));
    LocalMux I__6994 (
            .O(N__35414),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ));
    InMux I__6993 (
            .O(N__35411),
            .I(N__35408));
    LocalMux I__6992 (
            .O(N__35408),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ));
    InMux I__6991 (
            .O(N__35405),
            .I(N__35402));
    LocalMux I__6990 (
            .O(N__35402),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ));
    InMux I__6989 (
            .O(N__35399),
            .I(N__35396));
    LocalMux I__6988 (
            .O(N__35396),
            .I(\current_shift_inst.un38_control_input_0_s0_19 ));
    InMux I__6987 (
            .O(N__35393),
            .I(N__35390));
    LocalMux I__6986 (
            .O(N__35390),
            .I(N__35387));
    Odrv4 I__6985 (
            .O(N__35387),
            .I(\current_shift_inst.control_input_axb_16 ));
    InMux I__6984 (
            .O(N__35384),
            .I(N__35381));
    LocalMux I__6983 (
            .O(N__35381),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__6982 (
            .O(N__35378),
            .I(N__35375));
    LocalMux I__6981 (
            .O(N__35375),
            .I(N__35372));
    Odrv4 I__6980 (
            .O(N__35372),
            .I(\current_shift_inst.control_input_axb_25 ));
    InMux I__6979 (
            .O(N__35369),
            .I(N__35366));
    LocalMux I__6978 (
            .O(N__35366),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ));
    InMux I__6977 (
            .O(N__35363),
            .I(N__35360));
    LocalMux I__6976 (
            .O(N__35360),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ));
    CascadeMux I__6975 (
            .O(N__35357),
            .I(N__35354));
    InMux I__6974 (
            .O(N__35354),
            .I(N__35351));
    LocalMux I__6973 (
            .O(N__35351),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ));
    CascadeMux I__6972 (
            .O(N__35348),
            .I(N__35345));
    InMux I__6971 (
            .O(N__35345),
            .I(N__35342));
    LocalMux I__6970 (
            .O(N__35342),
            .I(\current_shift_inst.un38_control_input_0_s0_14 ));
    CascadeMux I__6969 (
            .O(N__35339),
            .I(N__35336));
    InMux I__6968 (
            .O(N__35336),
            .I(N__35333));
    LocalMux I__6967 (
            .O(N__35333),
            .I(N__35330));
    Odrv4 I__6966 (
            .O(N__35330),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__6965 (
            .O(N__35327),
            .I(N__35324));
    LocalMux I__6964 (
            .O(N__35324),
            .I(\current_shift_inst.un38_control_input_0_s0_15 ));
    InMux I__6963 (
            .O(N__35321),
            .I(N__35318));
    LocalMux I__6962 (
            .O(N__35318),
            .I(N__35315));
    Odrv4 I__6961 (
            .O(N__35315),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__6960 (
            .O(N__35312),
            .I(N__35309));
    LocalMux I__6959 (
            .O(N__35309),
            .I(N__35306));
    Odrv4 I__6958 (
            .O(N__35306),
            .I(\current_shift_inst.un38_control_input_0_s0_16 ));
    InMux I__6957 (
            .O(N__35303),
            .I(N__35300));
    LocalMux I__6956 (
            .O(N__35300),
            .I(N__35297));
    Odrv4 I__6955 (
            .O(N__35297),
            .I(\current_shift_inst.control_input_axb_13 ));
    InMux I__6954 (
            .O(N__35294),
            .I(N__35291));
    LocalMux I__6953 (
            .O(N__35291),
            .I(N__35288));
    Odrv4 I__6952 (
            .O(N__35288),
            .I(\current_shift_inst.un38_control_input_0_s0_17 ));
    InMux I__6951 (
            .O(N__35285),
            .I(N__35282));
    LocalMux I__6950 (
            .O(N__35282),
            .I(N__35279));
    Odrv4 I__6949 (
            .O(N__35279),
            .I(\current_shift_inst.control_input_axb_14 ));
    InMux I__6948 (
            .O(N__35276),
            .I(N__35273));
    LocalMux I__6947 (
            .O(N__35273),
            .I(N__35270));
    Odrv4 I__6946 (
            .O(N__35270),
            .I(\current_shift_inst.un38_control_input_0_s0_18 ));
    InMux I__6945 (
            .O(N__35267),
            .I(N__35264));
    LocalMux I__6944 (
            .O(N__35264),
            .I(N__35261));
    Odrv4 I__6943 (
            .O(N__35261),
            .I(\current_shift_inst.control_input_axb_15 ));
    InMux I__6942 (
            .O(N__35258),
            .I(N__35255));
    LocalMux I__6941 (
            .O(N__35255),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ));
    InMux I__6940 (
            .O(N__35252),
            .I(N__35246));
    InMux I__6939 (
            .O(N__35251),
            .I(N__35246));
    LocalMux I__6938 (
            .O(N__35246),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ));
    CascadeMux I__6937 (
            .O(N__35243),
            .I(N__35240));
    InMux I__6936 (
            .O(N__35240),
            .I(N__35234));
    InMux I__6935 (
            .O(N__35239),
            .I(N__35234));
    LocalMux I__6934 (
            .O(N__35234),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ));
    CascadeMux I__6933 (
            .O(N__35231),
            .I(N__35228));
    InMux I__6932 (
            .O(N__35228),
            .I(N__35222));
    InMux I__6931 (
            .O(N__35227),
            .I(N__35222));
    LocalMux I__6930 (
            .O(N__35222),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    InMux I__6929 (
            .O(N__35219),
            .I(N__35213));
    InMux I__6928 (
            .O(N__35218),
            .I(N__35213));
    LocalMux I__6927 (
            .O(N__35213),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    InMux I__6926 (
            .O(N__35210),
            .I(N__35207));
    LocalMux I__6925 (
            .O(N__35207),
            .I(N__35204));
    Odrv4 I__6924 (
            .O(N__35204),
            .I(\current_shift_inst.un38_control_input_0_s0_10 ));
    InMux I__6923 (
            .O(N__35201),
            .I(N__35198));
    LocalMux I__6922 (
            .O(N__35198),
            .I(N__35195));
    Odrv4 I__6921 (
            .O(N__35195),
            .I(\current_shift_inst.control_input_axb_7 ));
    CascadeMux I__6920 (
            .O(N__35192),
            .I(N__35189));
    InMux I__6919 (
            .O(N__35189),
            .I(N__35186));
    LocalMux I__6918 (
            .O(N__35186),
            .I(N__35183));
    Odrv4 I__6917 (
            .O(N__35183),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ));
    InMux I__6916 (
            .O(N__35180),
            .I(N__35174));
    InMux I__6915 (
            .O(N__35179),
            .I(N__35174));
    LocalMux I__6914 (
            .O(N__35174),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    CascadeMux I__6913 (
            .O(N__35171),
            .I(N__35165));
    InMux I__6912 (
            .O(N__35170),
            .I(N__35161));
    InMux I__6911 (
            .O(N__35169),
            .I(N__35158));
    InMux I__6910 (
            .O(N__35168),
            .I(N__35155));
    InMux I__6909 (
            .O(N__35165),
            .I(N__35152));
    InMux I__6908 (
            .O(N__35164),
            .I(N__35149));
    LocalMux I__6907 (
            .O(N__35161),
            .I(N__35146));
    LocalMux I__6906 (
            .O(N__35158),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__6905 (
            .O(N__35155),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__6904 (
            .O(N__35152),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__6903 (
            .O(N__35149),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv12 I__6902 (
            .O(N__35146),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__6901 (
            .O(N__35135),
            .I(N__35131));
    InMux I__6900 (
            .O(N__35134),
            .I(N__35128));
    LocalMux I__6899 (
            .O(N__35131),
            .I(N__35124));
    LocalMux I__6898 (
            .O(N__35128),
            .I(N__35121));
    InMux I__6897 (
            .O(N__35127),
            .I(N__35118));
    Span4Mux_h I__6896 (
            .O(N__35124),
            .I(N__35111));
    Span4Mux_v I__6895 (
            .O(N__35121),
            .I(N__35111));
    LocalMux I__6894 (
            .O(N__35118),
            .I(N__35111));
    Odrv4 I__6893 (
            .O(N__35111),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__6892 (
            .O(N__35108),
            .I(N__35104));
    InMux I__6891 (
            .O(N__35107),
            .I(N__35101));
    LocalMux I__6890 (
            .O(N__35104),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    LocalMux I__6889 (
            .O(N__35101),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    InMux I__6888 (
            .O(N__35096),
            .I(N__35093));
    LocalMux I__6887 (
            .O(N__35093),
            .I(N__35088));
    InMux I__6886 (
            .O(N__35092),
            .I(N__35083));
    InMux I__6885 (
            .O(N__35091),
            .I(N__35083));
    Odrv4 I__6884 (
            .O(N__35088),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__6883 (
            .O(N__35083),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__6882 (
            .O(N__35078),
            .I(N__35075));
    InMux I__6881 (
            .O(N__35075),
            .I(N__35071));
    InMux I__6880 (
            .O(N__35074),
            .I(N__35068));
    LocalMux I__6879 (
            .O(N__35071),
            .I(N__35061));
    LocalMux I__6878 (
            .O(N__35068),
            .I(N__35061));
    InMux I__6877 (
            .O(N__35067),
            .I(N__35056));
    InMux I__6876 (
            .O(N__35066),
            .I(N__35056));
    Odrv12 I__6875 (
            .O(N__35061),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    LocalMux I__6874 (
            .O(N__35056),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__6873 (
            .O(N__35051),
            .I(N__35048));
    LocalMux I__6872 (
            .O(N__35048),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    InMux I__6871 (
            .O(N__35045),
            .I(N__35042));
    LocalMux I__6870 (
            .O(N__35042),
            .I(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ));
    InMux I__6869 (
            .O(N__35039),
            .I(N__35031));
    InMux I__6868 (
            .O(N__35038),
            .I(N__35031));
    InMux I__6867 (
            .O(N__35037),
            .I(N__35026));
    InMux I__6866 (
            .O(N__35036),
            .I(N__35026));
    LocalMux I__6865 (
            .O(N__35031),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__6864 (
            .O(N__35026),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__6863 (
            .O(N__35021),
            .I(N__35017));
    CascadeMux I__6862 (
            .O(N__35020),
            .I(N__35014));
    InMux I__6861 (
            .O(N__35017),
            .I(N__35008));
    InMux I__6860 (
            .O(N__35014),
            .I(N__35005));
    InMux I__6859 (
            .O(N__35013),
            .I(N__35000));
    InMux I__6858 (
            .O(N__35012),
            .I(N__35000));
    InMux I__6857 (
            .O(N__35011),
            .I(N__34997));
    LocalMux I__6856 (
            .O(N__35008),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__6855 (
            .O(N__35005),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__6854 (
            .O(N__35000),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__6853 (
            .O(N__34997),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    InMux I__6852 (
            .O(N__34988),
            .I(N__34983));
    InMux I__6851 (
            .O(N__34987),
            .I(N__34980));
    InMux I__6850 (
            .O(N__34986),
            .I(N__34977));
    LocalMux I__6849 (
            .O(N__34983),
            .I(N__34974));
    LocalMux I__6848 (
            .O(N__34980),
            .I(N__34969));
    LocalMux I__6847 (
            .O(N__34977),
            .I(N__34969));
    Sp12to4 I__6846 (
            .O(N__34974),
            .I(N__34964));
    Sp12to4 I__6845 (
            .O(N__34969),
            .I(N__34964));
    Span12Mux_v I__6844 (
            .O(N__34964),
            .I(N__34961));
    Odrv12 I__6843 (
            .O(N__34961),
            .I(il_min_comp1_D2));
    CascadeMux I__6842 (
            .O(N__34958),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24_cascade_));
    InMux I__6841 (
            .O(N__34955),
            .I(N__34949));
    InMux I__6840 (
            .O(N__34954),
            .I(N__34949));
    LocalMux I__6839 (
            .O(N__34949),
            .I(N__34945));
    InMux I__6838 (
            .O(N__34948),
            .I(N__34942));
    Span4Mux_h I__6837 (
            .O(N__34945),
            .I(N__34939));
    LocalMux I__6836 (
            .O(N__34942),
            .I(N__34935));
    Span4Mux_h I__6835 (
            .O(N__34939),
            .I(N__34932));
    InMux I__6834 (
            .O(N__34938),
            .I(N__34929));
    Odrv4 I__6833 (
            .O(N__34935),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv4 I__6832 (
            .O(N__34932),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    LocalMux I__6831 (
            .O(N__34929),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__6830 (
            .O(N__34922),
            .I(N__34916));
    InMux I__6829 (
            .O(N__34921),
            .I(N__34916));
    LocalMux I__6828 (
            .O(N__34916),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ));
    InMux I__6827 (
            .O(N__34913),
            .I(N__34910));
    LocalMux I__6826 (
            .O(N__34910),
            .I(N__34906));
    InMux I__6825 (
            .O(N__34909),
            .I(N__34902));
    Span4Mux_h I__6824 (
            .O(N__34906),
            .I(N__34899));
    InMux I__6823 (
            .O(N__34905),
            .I(N__34896));
    LocalMux I__6822 (
            .O(N__34902),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv4 I__6821 (
            .O(N__34899),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    LocalMux I__6820 (
            .O(N__34896),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    InMux I__6819 (
            .O(N__34889),
            .I(N__34886));
    LocalMux I__6818 (
            .O(N__34886),
            .I(N__34882));
    InMux I__6817 (
            .O(N__34885),
            .I(N__34878));
    Span4Mux_v I__6816 (
            .O(N__34882),
            .I(N__34875));
    InMux I__6815 (
            .O(N__34881),
            .I(N__34872));
    LocalMux I__6814 (
            .O(N__34878),
            .I(N__34868));
    Sp12to4 I__6813 (
            .O(N__34875),
            .I(N__34863));
    LocalMux I__6812 (
            .O(N__34872),
            .I(N__34863));
    InMux I__6811 (
            .O(N__34871),
            .I(N__34860));
    Odrv4 I__6810 (
            .O(N__34868),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv12 I__6809 (
            .O(N__34863),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    LocalMux I__6808 (
            .O(N__34860),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__6807 (
            .O(N__34853),
            .I(N__34850));
    LocalMux I__6806 (
            .O(N__34850),
            .I(N__34847));
    Odrv12 I__6805 (
            .O(N__34847),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__6804 (
            .O(N__34844),
            .I(N__34825));
    InMux I__6803 (
            .O(N__34843),
            .I(N__34818));
    InMux I__6802 (
            .O(N__34842),
            .I(N__34818));
    InMux I__6801 (
            .O(N__34841),
            .I(N__34818));
    InMux I__6800 (
            .O(N__34840),
            .I(N__34810));
    InMux I__6799 (
            .O(N__34839),
            .I(N__34810));
    InMux I__6798 (
            .O(N__34838),
            .I(N__34795));
    InMux I__6797 (
            .O(N__34837),
            .I(N__34795));
    InMux I__6796 (
            .O(N__34836),
            .I(N__34795));
    InMux I__6795 (
            .O(N__34835),
            .I(N__34795));
    InMux I__6794 (
            .O(N__34834),
            .I(N__34795));
    InMux I__6793 (
            .O(N__34833),
            .I(N__34795));
    InMux I__6792 (
            .O(N__34832),
            .I(N__34795));
    InMux I__6791 (
            .O(N__34831),
            .I(N__34786));
    InMux I__6790 (
            .O(N__34830),
            .I(N__34786));
    InMux I__6789 (
            .O(N__34829),
            .I(N__34786));
    InMux I__6788 (
            .O(N__34828),
            .I(N__34786));
    LocalMux I__6787 (
            .O(N__34825),
            .I(N__34781));
    LocalMux I__6786 (
            .O(N__34818),
            .I(N__34781));
    InMux I__6785 (
            .O(N__34817),
            .I(N__34762));
    InMux I__6784 (
            .O(N__34816),
            .I(N__34759));
    InMux I__6783 (
            .O(N__34815),
            .I(N__34743));
    LocalMux I__6782 (
            .O(N__34810),
            .I(N__34723));
    LocalMux I__6781 (
            .O(N__34795),
            .I(N__34723));
    LocalMux I__6780 (
            .O(N__34786),
            .I(N__34723));
    Span4Mux_v I__6779 (
            .O(N__34781),
            .I(N__34723));
    InMux I__6778 (
            .O(N__34780),
            .I(N__34712));
    InMux I__6777 (
            .O(N__34779),
            .I(N__34712));
    InMux I__6776 (
            .O(N__34778),
            .I(N__34712));
    InMux I__6775 (
            .O(N__34777),
            .I(N__34712));
    InMux I__6774 (
            .O(N__34776),
            .I(N__34712));
    InMux I__6773 (
            .O(N__34775),
            .I(N__34704));
    InMux I__6772 (
            .O(N__34774),
            .I(N__34704));
    InMux I__6771 (
            .O(N__34773),
            .I(N__34691));
    InMux I__6770 (
            .O(N__34772),
            .I(N__34691));
    InMux I__6769 (
            .O(N__34771),
            .I(N__34691));
    InMux I__6768 (
            .O(N__34770),
            .I(N__34691));
    InMux I__6767 (
            .O(N__34769),
            .I(N__34691));
    InMux I__6766 (
            .O(N__34768),
            .I(N__34691));
    InMux I__6765 (
            .O(N__34767),
            .I(N__34686));
    InMux I__6764 (
            .O(N__34766),
            .I(N__34686));
    CascadeMux I__6763 (
            .O(N__34765),
            .I(N__34680));
    LocalMux I__6762 (
            .O(N__34762),
            .I(N__34674));
    LocalMux I__6761 (
            .O(N__34759),
            .I(N__34674));
    InMux I__6760 (
            .O(N__34758),
            .I(N__34663));
    InMux I__6759 (
            .O(N__34757),
            .I(N__34660));
    InMux I__6758 (
            .O(N__34756),
            .I(N__34647));
    InMux I__6757 (
            .O(N__34755),
            .I(N__34647));
    InMux I__6756 (
            .O(N__34754),
            .I(N__34647));
    InMux I__6755 (
            .O(N__34753),
            .I(N__34647));
    InMux I__6754 (
            .O(N__34752),
            .I(N__34647));
    InMux I__6753 (
            .O(N__34751),
            .I(N__34647));
    InMux I__6752 (
            .O(N__34750),
            .I(N__34636));
    InMux I__6751 (
            .O(N__34749),
            .I(N__34636));
    InMux I__6750 (
            .O(N__34748),
            .I(N__34636));
    InMux I__6749 (
            .O(N__34747),
            .I(N__34636));
    InMux I__6748 (
            .O(N__34746),
            .I(N__34636));
    LocalMux I__6747 (
            .O(N__34743),
            .I(N__34633));
    InMux I__6746 (
            .O(N__34742),
            .I(N__34630));
    InMux I__6745 (
            .O(N__34741),
            .I(N__34623));
    InMux I__6744 (
            .O(N__34740),
            .I(N__34623));
    InMux I__6743 (
            .O(N__34739),
            .I(N__34623));
    InMux I__6742 (
            .O(N__34738),
            .I(N__34620));
    InMux I__6741 (
            .O(N__34737),
            .I(N__34615));
    InMux I__6740 (
            .O(N__34736),
            .I(N__34615));
    InMux I__6739 (
            .O(N__34735),
            .I(N__34590));
    InMux I__6738 (
            .O(N__34734),
            .I(N__34590));
    InMux I__6737 (
            .O(N__34733),
            .I(N__34590));
    InMux I__6736 (
            .O(N__34732),
            .I(N__34590));
    Span4Mux_v I__6735 (
            .O(N__34723),
            .I(N__34585));
    LocalMux I__6734 (
            .O(N__34712),
            .I(N__34585));
    CascadeMux I__6733 (
            .O(N__34711),
            .I(N__34582));
    InMux I__6732 (
            .O(N__34710),
            .I(N__34578));
    InMux I__6731 (
            .O(N__34709),
            .I(N__34575));
    LocalMux I__6730 (
            .O(N__34704),
            .I(N__34568));
    LocalMux I__6729 (
            .O(N__34691),
            .I(N__34568));
    LocalMux I__6728 (
            .O(N__34686),
            .I(N__34568));
    InMux I__6727 (
            .O(N__34685),
            .I(N__34557));
    InMux I__6726 (
            .O(N__34684),
            .I(N__34557));
    InMux I__6725 (
            .O(N__34683),
            .I(N__34557));
    InMux I__6724 (
            .O(N__34680),
            .I(N__34557));
    InMux I__6723 (
            .O(N__34679),
            .I(N__34557));
    Span4Mux_v I__6722 (
            .O(N__34674),
            .I(N__34554));
    InMux I__6721 (
            .O(N__34673),
            .I(N__34551));
    InMux I__6720 (
            .O(N__34672),
            .I(N__34536));
    InMux I__6719 (
            .O(N__34671),
            .I(N__34536));
    InMux I__6718 (
            .O(N__34670),
            .I(N__34536));
    InMux I__6717 (
            .O(N__34669),
            .I(N__34536));
    InMux I__6716 (
            .O(N__34668),
            .I(N__34536));
    InMux I__6715 (
            .O(N__34667),
            .I(N__34536));
    InMux I__6714 (
            .O(N__34666),
            .I(N__34536));
    LocalMux I__6713 (
            .O(N__34663),
            .I(N__34533));
    LocalMux I__6712 (
            .O(N__34660),
            .I(N__34530));
    LocalMux I__6711 (
            .O(N__34647),
            .I(N__34525));
    LocalMux I__6710 (
            .O(N__34636),
            .I(N__34525));
    Span4Mux_v I__6709 (
            .O(N__34633),
            .I(N__34520));
    LocalMux I__6708 (
            .O(N__34630),
            .I(N__34520));
    LocalMux I__6707 (
            .O(N__34623),
            .I(N__34517));
    LocalMux I__6706 (
            .O(N__34620),
            .I(N__34512));
    LocalMux I__6705 (
            .O(N__34615),
            .I(N__34512));
    InMux I__6704 (
            .O(N__34614),
            .I(N__34507));
    InMux I__6703 (
            .O(N__34613),
            .I(N__34507));
    InMux I__6702 (
            .O(N__34612),
            .I(N__34504));
    InMux I__6701 (
            .O(N__34611),
            .I(N__34491));
    InMux I__6700 (
            .O(N__34610),
            .I(N__34491));
    InMux I__6699 (
            .O(N__34609),
            .I(N__34491));
    InMux I__6698 (
            .O(N__34608),
            .I(N__34491));
    InMux I__6697 (
            .O(N__34607),
            .I(N__34491));
    InMux I__6696 (
            .O(N__34606),
            .I(N__34491));
    InMux I__6695 (
            .O(N__34605),
            .I(N__34486));
    InMux I__6694 (
            .O(N__34604),
            .I(N__34486));
    InMux I__6693 (
            .O(N__34603),
            .I(N__34475));
    InMux I__6692 (
            .O(N__34602),
            .I(N__34475));
    InMux I__6691 (
            .O(N__34601),
            .I(N__34475));
    InMux I__6690 (
            .O(N__34600),
            .I(N__34475));
    InMux I__6689 (
            .O(N__34599),
            .I(N__34475));
    LocalMux I__6688 (
            .O(N__34590),
            .I(N__34472));
    Span4Mux_h I__6687 (
            .O(N__34585),
            .I(N__34469));
    InMux I__6686 (
            .O(N__34582),
            .I(N__34464));
    InMux I__6685 (
            .O(N__34581),
            .I(N__34464));
    LocalMux I__6684 (
            .O(N__34578),
            .I(N__34459));
    LocalMux I__6683 (
            .O(N__34575),
            .I(N__34459));
    Span4Mux_v I__6682 (
            .O(N__34568),
            .I(N__34452));
    LocalMux I__6681 (
            .O(N__34557),
            .I(N__34452));
    Span4Mux_h I__6680 (
            .O(N__34554),
            .I(N__34452));
    LocalMux I__6679 (
            .O(N__34551),
            .I(N__34435));
    LocalMux I__6678 (
            .O(N__34536),
            .I(N__34435));
    Span4Mux_v I__6677 (
            .O(N__34533),
            .I(N__34435));
    Span4Mux_v I__6676 (
            .O(N__34530),
            .I(N__34435));
    Span4Mux_v I__6675 (
            .O(N__34525),
            .I(N__34435));
    Span4Mux_v I__6674 (
            .O(N__34520),
            .I(N__34435));
    Span4Mux_h I__6673 (
            .O(N__34517),
            .I(N__34435));
    Span4Mux_v I__6672 (
            .O(N__34512),
            .I(N__34435));
    LocalMux I__6671 (
            .O(N__34507),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__6670 (
            .O(N__34504),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__6669 (
            .O(N__34491),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__6668 (
            .O(N__34486),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__6667 (
            .O(N__34475),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__6666 (
            .O(N__34472),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__6665 (
            .O(N__34469),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__6664 (
            .O(N__34464),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__6663 (
            .O(N__34459),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__6662 (
            .O(N__34452),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__6661 (
            .O(N__34435),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    InMux I__6660 (
            .O(N__34412),
            .I(N__34409));
    LocalMux I__6659 (
            .O(N__34409),
            .I(N__34405));
    InMux I__6658 (
            .O(N__34408),
            .I(N__34401));
    Span4Mux_h I__6657 (
            .O(N__34405),
            .I(N__34398));
    InMux I__6656 (
            .O(N__34404),
            .I(N__34395));
    LocalMux I__6655 (
            .O(N__34401),
            .I(N__34390));
    Span4Mux_v I__6654 (
            .O(N__34398),
            .I(N__34390));
    LocalMux I__6653 (
            .O(N__34395),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    Odrv4 I__6652 (
            .O(N__34390),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    InMux I__6651 (
            .O(N__34385),
            .I(N__34381));
    InMux I__6650 (
            .O(N__34384),
            .I(N__34378));
    LocalMux I__6649 (
            .O(N__34381),
            .I(N__34375));
    LocalMux I__6648 (
            .O(N__34378),
            .I(N__34371));
    Span4Mux_v I__6647 (
            .O(N__34375),
            .I(N__34368));
    InMux I__6646 (
            .O(N__34374),
            .I(N__34365));
    Span12Mux_h I__6645 (
            .O(N__34371),
            .I(N__34361));
    Sp12to4 I__6644 (
            .O(N__34368),
            .I(N__34356));
    LocalMux I__6643 (
            .O(N__34365),
            .I(N__34356));
    InMux I__6642 (
            .O(N__34364),
            .I(N__34353));
    Odrv12 I__6641 (
            .O(N__34361),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv12 I__6640 (
            .O(N__34356),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    LocalMux I__6639 (
            .O(N__34353),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__6638 (
            .O(N__34346),
            .I(N__34343));
    LocalMux I__6637 (
            .O(N__34343),
            .I(N__34340));
    Odrv4 I__6636 (
            .O(N__34340),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CEMux I__6635 (
            .O(N__34337),
            .I(N__34334));
    LocalMux I__6634 (
            .O(N__34334),
            .I(N__34313));
    InMux I__6633 (
            .O(N__34333),
            .I(N__34302));
    InMux I__6632 (
            .O(N__34332),
            .I(N__34302));
    InMux I__6631 (
            .O(N__34331),
            .I(N__34302));
    InMux I__6630 (
            .O(N__34330),
            .I(N__34293));
    InMux I__6629 (
            .O(N__34329),
            .I(N__34293));
    InMux I__6628 (
            .O(N__34328),
            .I(N__34293));
    InMux I__6627 (
            .O(N__34327),
            .I(N__34293));
    InMux I__6626 (
            .O(N__34326),
            .I(N__34284));
    InMux I__6625 (
            .O(N__34325),
            .I(N__34284));
    InMux I__6624 (
            .O(N__34324),
            .I(N__34284));
    InMux I__6623 (
            .O(N__34323),
            .I(N__34284));
    CEMux I__6622 (
            .O(N__34322),
            .I(N__34281));
    CEMux I__6621 (
            .O(N__34321),
            .I(N__34277));
    InMux I__6620 (
            .O(N__34320),
            .I(N__34267));
    InMux I__6619 (
            .O(N__34319),
            .I(N__34267));
    InMux I__6618 (
            .O(N__34318),
            .I(N__34267));
    InMux I__6617 (
            .O(N__34317),
            .I(N__34267));
    CEMux I__6616 (
            .O(N__34316),
            .I(N__34264));
    Span4Mux_v I__6615 (
            .O(N__34313),
            .I(N__34258));
    CEMux I__6614 (
            .O(N__34312),
            .I(N__34255));
    InMux I__6613 (
            .O(N__34311),
            .I(N__34247));
    InMux I__6612 (
            .O(N__34310),
            .I(N__34247));
    InMux I__6611 (
            .O(N__34309),
            .I(N__34247));
    LocalMux I__6610 (
            .O(N__34302),
            .I(N__34238));
    LocalMux I__6609 (
            .O(N__34293),
            .I(N__34238));
    LocalMux I__6608 (
            .O(N__34284),
            .I(N__34238));
    LocalMux I__6607 (
            .O(N__34281),
            .I(N__34238));
    CEMux I__6606 (
            .O(N__34280),
            .I(N__34223));
    LocalMux I__6605 (
            .O(N__34277),
            .I(N__34220));
    CEMux I__6604 (
            .O(N__34276),
            .I(N__34217));
    LocalMux I__6603 (
            .O(N__34267),
            .I(N__34212));
    LocalMux I__6602 (
            .O(N__34264),
            .I(N__34212));
    CEMux I__6601 (
            .O(N__34263),
            .I(N__34209));
    CEMux I__6600 (
            .O(N__34262),
            .I(N__34206));
    CEMux I__6599 (
            .O(N__34261),
            .I(N__34203));
    Span4Mux_h I__6598 (
            .O(N__34258),
            .I(N__34197));
    LocalMux I__6597 (
            .O(N__34255),
            .I(N__34197));
    CEMux I__6596 (
            .O(N__34254),
            .I(N__34194));
    LocalMux I__6595 (
            .O(N__34247),
            .I(N__34189));
    Span4Mux_v I__6594 (
            .O(N__34238),
            .I(N__34189));
    InMux I__6593 (
            .O(N__34237),
            .I(N__34180));
    InMux I__6592 (
            .O(N__34236),
            .I(N__34180));
    InMux I__6591 (
            .O(N__34235),
            .I(N__34180));
    InMux I__6590 (
            .O(N__34234),
            .I(N__34180));
    InMux I__6589 (
            .O(N__34233),
            .I(N__34171));
    InMux I__6588 (
            .O(N__34232),
            .I(N__34171));
    InMux I__6587 (
            .O(N__34231),
            .I(N__34171));
    InMux I__6586 (
            .O(N__34230),
            .I(N__34171));
    InMux I__6585 (
            .O(N__34229),
            .I(N__34162));
    InMux I__6584 (
            .O(N__34228),
            .I(N__34162));
    InMux I__6583 (
            .O(N__34227),
            .I(N__34162));
    InMux I__6582 (
            .O(N__34226),
            .I(N__34162));
    LocalMux I__6581 (
            .O(N__34223),
            .I(N__34159));
    Span4Mux_v I__6580 (
            .O(N__34220),
            .I(N__34154));
    LocalMux I__6579 (
            .O(N__34217),
            .I(N__34154));
    Span4Mux_h I__6578 (
            .O(N__34212),
            .I(N__34151));
    LocalMux I__6577 (
            .O(N__34209),
            .I(N__34148));
    LocalMux I__6576 (
            .O(N__34206),
            .I(N__34145));
    LocalMux I__6575 (
            .O(N__34203),
            .I(N__34142));
    CEMux I__6574 (
            .O(N__34202),
            .I(N__34138));
    Span4Mux_h I__6573 (
            .O(N__34197),
            .I(N__34135));
    LocalMux I__6572 (
            .O(N__34194),
            .I(N__34132));
    Span4Mux_h I__6571 (
            .O(N__34189),
            .I(N__34121));
    LocalMux I__6570 (
            .O(N__34180),
            .I(N__34121));
    LocalMux I__6569 (
            .O(N__34171),
            .I(N__34121));
    LocalMux I__6568 (
            .O(N__34162),
            .I(N__34121));
    Span4Mux_h I__6567 (
            .O(N__34159),
            .I(N__34121));
    Span4Mux_v I__6566 (
            .O(N__34154),
            .I(N__34118));
    Span4Mux_v I__6565 (
            .O(N__34151),
            .I(N__34115));
    Span4Mux_h I__6564 (
            .O(N__34148),
            .I(N__34110));
    Span4Mux_v I__6563 (
            .O(N__34145),
            .I(N__34110));
    Span4Mux_v I__6562 (
            .O(N__34142),
            .I(N__34107));
    InMux I__6561 (
            .O(N__34141),
            .I(N__34104));
    LocalMux I__6560 (
            .O(N__34138),
            .I(N__34099));
    Sp12to4 I__6559 (
            .O(N__34135),
            .I(N__34099));
    Span4Mux_h I__6558 (
            .O(N__34132),
            .I(N__34094));
    Span4Mux_v I__6557 (
            .O(N__34121),
            .I(N__34094));
    Span4Mux_h I__6556 (
            .O(N__34118),
            .I(N__34089));
    Span4Mux_h I__6555 (
            .O(N__34115),
            .I(N__34089));
    Odrv4 I__6554 (
            .O(N__34110),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__6553 (
            .O(N__34107),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__6552 (
            .O(N__34104),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv12 I__6551 (
            .O(N__34099),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__6550 (
            .O(N__34094),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__6549 (
            .O(N__34089),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    InMux I__6548 (
            .O(N__34076),
            .I(N__34070));
    InMux I__6547 (
            .O(N__34075),
            .I(N__34070));
    LocalMux I__6546 (
            .O(N__34070),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ));
    IoInMux I__6545 (
            .O(N__34067),
            .I(N__34064));
    LocalMux I__6544 (
            .O(N__34064),
            .I(N__34061));
    Span4Mux_s0_v I__6543 (
            .O(N__34061),
            .I(N__34058));
    Odrv4 I__6542 (
            .O(N__34058),
            .I(\pll_inst.red_c_i ));
    ClkMux I__6541 (
            .O(N__34055),
            .I(N__34049));
    ClkMux I__6540 (
            .O(N__34054),
            .I(N__34049));
    GlobalMux I__6539 (
            .O(N__34049),
            .I(N__34046));
    gio2CtrlBuf I__6538 (
            .O(N__34046),
            .I(delay_hc_input_c_g));
    InMux I__6537 (
            .O(N__34043),
            .I(N__34040));
    LocalMux I__6536 (
            .O(N__34040),
            .I(N__34035));
    InMux I__6535 (
            .O(N__34039),
            .I(N__34032));
    InMux I__6534 (
            .O(N__34038),
            .I(N__34029));
    Span4Mux_v I__6533 (
            .O(N__34035),
            .I(N__34026));
    LocalMux I__6532 (
            .O(N__34032),
            .I(N__34023));
    LocalMux I__6531 (
            .O(N__34029),
            .I(N__34020));
    Span4Mux_v I__6530 (
            .O(N__34026),
            .I(N__34014));
    Span4Mux_v I__6529 (
            .O(N__34023),
            .I(N__34014));
    Span12Mux_v I__6528 (
            .O(N__34020),
            .I(N__34011));
    InMux I__6527 (
            .O(N__34019),
            .I(N__34008));
    Odrv4 I__6526 (
            .O(N__34014),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    Odrv12 I__6525 (
            .O(N__34011),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__6524 (
            .O(N__34008),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__6523 (
            .O(N__34001),
            .I(N__33998));
    LocalMux I__6522 (
            .O(N__33998),
            .I(N__33993));
    InMux I__6521 (
            .O(N__33997),
            .I(N__33990));
    InMux I__6520 (
            .O(N__33996),
            .I(N__33987));
    Span4Mux_h I__6519 (
            .O(N__33993),
            .I(N__33984));
    LocalMux I__6518 (
            .O(N__33990),
            .I(N__33981));
    LocalMux I__6517 (
            .O(N__33987),
            .I(N__33974));
    Span4Mux_v I__6516 (
            .O(N__33984),
            .I(N__33974));
    Span4Mux_v I__6515 (
            .O(N__33981),
            .I(N__33974));
    Odrv4 I__6514 (
            .O(N__33974),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    CascadeMux I__6513 (
            .O(N__33971),
            .I(N__33968));
    InMux I__6512 (
            .O(N__33968),
            .I(N__33965));
    LocalMux I__6511 (
            .O(N__33965),
            .I(N__33962));
    Span4Mux_h I__6510 (
            .O(N__33962),
            .I(N__33959));
    Odrv4 I__6509 (
            .O(N__33959),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt24 ));
    InMux I__6508 (
            .O(N__33956),
            .I(N__33951));
    InMux I__6507 (
            .O(N__33955),
            .I(N__33946));
    InMux I__6506 (
            .O(N__33954),
            .I(N__33946));
    LocalMux I__6505 (
            .O(N__33951),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    LocalMux I__6504 (
            .O(N__33946),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    CascadeMux I__6503 (
            .O(N__33941),
            .I(N__33938));
    InMux I__6502 (
            .O(N__33938),
            .I(N__33931));
    InMux I__6501 (
            .O(N__33937),
            .I(N__33931));
    InMux I__6500 (
            .O(N__33936),
            .I(N__33928));
    LocalMux I__6499 (
            .O(N__33931),
            .I(N__33925));
    LocalMux I__6498 (
            .O(N__33928),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__6497 (
            .O(N__33925),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__6496 (
            .O(N__33920),
            .I(N__33917));
    LocalMux I__6495 (
            .O(N__33917),
            .I(N__33914));
    Span4Mux_h I__6494 (
            .O(N__33914),
            .I(N__33911));
    Odrv4 I__6493 (
            .O(N__33911),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ));
    InMux I__6492 (
            .O(N__33908),
            .I(N__33905));
    LocalMux I__6491 (
            .O(N__33905),
            .I(N__33902));
    Span4Mux_v I__6490 (
            .O(N__33902),
            .I(N__33897));
    InMux I__6489 (
            .O(N__33901),
            .I(N__33894));
    InMux I__6488 (
            .O(N__33900),
            .I(N__33891));
    Span4Mux_h I__6487 (
            .O(N__33897),
            .I(N__33888));
    LocalMux I__6486 (
            .O(N__33894),
            .I(N__33885));
    LocalMux I__6485 (
            .O(N__33891),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    Odrv4 I__6484 (
            .O(N__33888),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    Odrv4 I__6483 (
            .O(N__33885),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    InMux I__6482 (
            .O(N__33878),
            .I(N__33875));
    LocalMux I__6481 (
            .O(N__33875),
            .I(N__33871));
    InMux I__6480 (
            .O(N__33874),
            .I(N__33867));
    Span4Mux_h I__6479 (
            .O(N__33871),
            .I(N__33864));
    InMux I__6478 (
            .O(N__33870),
            .I(N__33861));
    LocalMux I__6477 (
            .O(N__33867),
            .I(N__33857));
    Span4Mux_h I__6476 (
            .O(N__33864),
            .I(N__33852));
    LocalMux I__6475 (
            .O(N__33861),
            .I(N__33852));
    InMux I__6474 (
            .O(N__33860),
            .I(N__33849));
    Odrv4 I__6473 (
            .O(N__33857),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__6472 (
            .O(N__33852),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    LocalMux I__6471 (
            .O(N__33849),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    CascadeMux I__6470 (
            .O(N__33842),
            .I(N__33839));
    InMux I__6469 (
            .O(N__33839),
            .I(N__33833));
    InMux I__6468 (
            .O(N__33838),
            .I(N__33833));
    LocalMux I__6467 (
            .O(N__33833),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ));
    InMux I__6466 (
            .O(N__33830),
            .I(N__33827));
    LocalMux I__6465 (
            .O(N__33827),
            .I(N__33824));
    Span4Mux_h I__6464 (
            .O(N__33824),
            .I(N__33820));
    InMux I__6463 (
            .O(N__33823),
            .I(N__33817));
    Odrv4 I__6462 (
            .O(N__33820),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    LocalMux I__6461 (
            .O(N__33817),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__6460 (
            .O(N__33812),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__6459 (
            .O(N__33809),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__6458 (
            .O(N__33806),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__6457 (
            .O(N__33803),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__6456 (
            .O(N__33800),
            .I(N__33797));
    LocalMux I__6455 (
            .O(N__33797),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__6454 (
            .O(N__33794),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__6453 (
            .O(N__33791),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__6452 (
            .O(N__33788),
            .I(N__33785));
    LocalMux I__6451 (
            .O(N__33785),
            .I(\current_shift_inst.control_input_axb_28 ));
    InMux I__6450 (
            .O(N__33782),
            .I(N__33779));
    LocalMux I__6449 (
            .O(N__33779),
            .I(N__33776));
    Odrv4 I__6448 (
            .O(N__33776),
            .I(\current_shift_inst.control_input_axb_29 ));
    InMux I__6447 (
            .O(N__33773),
            .I(\current_shift_inst.un38_control_input_cry_16_s0 ));
    InMux I__6446 (
            .O(N__33770),
            .I(\current_shift_inst.un38_control_input_cry_17_s0 ));
    InMux I__6445 (
            .O(N__33767),
            .I(\current_shift_inst.un38_control_input_cry_18_s0 ));
    InMux I__6444 (
            .O(N__33764),
            .I(N__33761));
    LocalMux I__6443 (
            .O(N__33761),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__6442 (
            .O(N__33758),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__6441 (
            .O(N__33755),
            .I(N__33752));
    LocalMux I__6440 (
            .O(N__33752),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__6439 (
            .O(N__33749),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__6438 (
            .O(N__33746),
            .I(N__33743));
    LocalMux I__6437 (
            .O(N__33743),
            .I(N__33740));
    Span4Mux_h I__6436 (
            .O(N__33740),
            .I(N__33737));
    Odrv4 I__6435 (
            .O(N__33737),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__6434 (
            .O(N__33734),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__6433 (
            .O(N__33731),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__6432 (
            .O(N__33728),
            .I(bfn_12_19_0_));
    InMux I__6431 (
            .O(N__33725),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__6430 (
            .O(N__33722),
            .I(N__33719));
    LocalMux I__6429 (
            .O(N__33719),
            .I(N__33716));
    Odrv4 I__6428 (
            .O(N__33716),
            .I(\current_shift_inst.un38_control_input_0_s0_9 ));
    InMux I__6427 (
            .O(N__33713),
            .I(\current_shift_inst.un38_control_input_cry_8_s0 ));
    InMux I__6426 (
            .O(N__33710),
            .I(\current_shift_inst.un38_control_input_cry_9_s0 ));
    InMux I__6425 (
            .O(N__33707),
            .I(N__33704));
    LocalMux I__6424 (
            .O(N__33704),
            .I(N__33701));
    Span4Mux_v I__6423 (
            .O(N__33701),
            .I(N__33698));
    Odrv4 I__6422 (
            .O(N__33698),
            .I(\current_shift_inst.un38_control_input_0_s0_11 ));
    InMux I__6421 (
            .O(N__33695),
            .I(\current_shift_inst.un38_control_input_cry_10_s0 ));
    InMux I__6420 (
            .O(N__33692),
            .I(N__33689));
    LocalMux I__6419 (
            .O(N__33689),
            .I(N__33686));
    Span4Mux_h I__6418 (
            .O(N__33686),
            .I(N__33683));
    Odrv4 I__6417 (
            .O(N__33683),
            .I(\current_shift_inst.un38_control_input_0_s0_12 ));
    InMux I__6416 (
            .O(N__33680),
            .I(\current_shift_inst.un38_control_input_cry_11_s0 ));
    InMux I__6415 (
            .O(N__33677),
            .I(N__33674));
    LocalMux I__6414 (
            .O(N__33674),
            .I(N__33671));
    Span4Mux_h I__6413 (
            .O(N__33671),
            .I(N__33668));
    Odrv4 I__6412 (
            .O(N__33668),
            .I(\current_shift_inst.un38_control_input_0_s0_13 ));
    InMux I__6411 (
            .O(N__33665),
            .I(\current_shift_inst.un38_control_input_cry_12_s0 ));
    InMux I__6410 (
            .O(N__33662),
            .I(\current_shift_inst.un38_control_input_cry_13_s0 ));
    InMux I__6409 (
            .O(N__33659),
            .I(\current_shift_inst.un38_control_input_cry_14_s0 ));
    InMux I__6408 (
            .O(N__33656),
            .I(bfn_12_18_0_));
    InMux I__6407 (
            .O(N__33653),
            .I(N__33650));
    LocalMux I__6406 (
            .O(N__33650),
            .I(N__33647));
    Span4Mux_h I__6405 (
            .O(N__33647),
            .I(N__33644));
    Odrv4 I__6404 (
            .O(N__33644),
            .I(\current_shift_inst.un38_control_input_0_s0_3 ));
    InMux I__6403 (
            .O(N__33641),
            .I(\current_shift_inst.un38_control_input_cry_2_s0 ));
    CascadeMux I__6402 (
            .O(N__33638),
            .I(N__33635));
    InMux I__6401 (
            .O(N__33635),
            .I(N__33632));
    LocalMux I__6400 (
            .O(N__33632),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ));
    InMux I__6399 (
            .O(N__33629),
            .I(N__33626));
    LocalMux I__6398 (
            .O(N__33626),
            .I(\current_shift_inst.un38_control_input_0_s0_4 ));
    InMux I__6397 (
            .O(N__33623),
            .I(\current_shift_inst.un38_control_input_cry_3_s0 ));
    InMux I__6396 (
            .O(N__33620),
            .I(N__33617));
    LocalMux I__6395 (
            .O(N__33617),
            .I(\current_shift_inst.un38_control_input_0_s0_5 ));
    InMux I__6394 (
            .O(N__33614),
            .I(\current_shift_inst.un38_control_input_cry_4_s0 ));
    InMux I__6393 (
            .O(N__33611),
            .I(N__33608));
    LocalMux I__6392 (
            .O(N__33608),
            .I(\current_shift_inst.un38_control_input_0_s0_6 ));
    InMux I__6391 (
            .O(N__33605),
            .I(\current_shift_inst.un38_control_input_cry_5_s0 ));
    InMux I__6390 (
            .O(N__33602),
            .I(N__33599));
    LocalMux I__6389 (
            .O(N__33599),
            .I(\current_shift_inst.un38_control_input_0_s0_7 ));
    InMux I__6388 (
            .O(N__33596),
            .I(\current_shift_inst.un38_control_input_cry_6_s0 ));
    InMux I__6387 (
            .O(N__33593),
            .I(N__33590));
    LocalMux I__6386 (
            .O(N__33590),
            .I(N__33587));
    Odrv4 I__6385 (
            .O(N__33587),
            .I(\current_shift_inst.un38_control_input_0_s0_8 ));
    InMux I__6384 (
            .O(N__33584),
            .I(bfn_12_17_0_));
    InMux I__6383 (
            .O(N__33581),
            .I(N__33578));
    LocalMux I__6382 (
            .O(N__33578),
            .I(N__33575));
    Span4Mux_h I__6381 (
            .O(N__33575),
            .I(N__33572));
    Span4Mux_h I__6380 (
            .O(N__33572),
            .I(N__33568));
    InMux I__6379 (
            .O(N__33571),
            .I(N__33565));
    Odrv4 I__6378 (
            .O(N__33568),
            .I(state_ns_i_a3_1));
    LocalMux I__6377 (
            .O(N__33565),
            .I(state_ns_i_a3_1));
    InMux I__6376 (
            .O(N__33560),
            .I(N__33557));
    LocalMux I__6375 (
            .O(N__33557),
            .I(N__33554));
    Span4Mux_h I__6374 (
            .O(N__33554),
            .I(N__33550));
    InMux I__6373 (
            .O(N__33553),
            .I(N__33547));
    Span4Mux_v I__6372 (
            .O(N__33550),
            .I(N__33540));
    LocalMux I__6371 (
            .O(N__33547),
            .I(N__33540));
    InMux I__6370 (
            .O(N__33546),
            .I(N__33535));
    InMux I__6369 (
            .O(N__33545),
            .I(N__33535));
    Sp12to4 I__6368 (
            .O(N__33540),
            .I(N__33532));
    LocalMux I__6367 (
            .O(N__33535),
            .I(N__33529));
    Span12Mux_v I__6366 (
            .O(N__33532),
            .I(N__33526));
    Span4Mux_v I__6365 (
            .O(N__33529),
            .I(N__33523));
    Span12Mux_v I__6364 (
            .O(N__33526),
            .I(N__33520));
    Sp12to4 I__6363 (
            .O(N__33523),
            .I(N__33517));
    Span12Mux_h I__6362 (
            .O(N__33520),
            .I(N__33514));
    Span12Mux_h I__6361 (
            .O(N__33517),
            .I(N__33511));
    Odrv12 I__6360 (
            .O(N__33514),
            .I(start_stop_c));
    Odrv12 I__6359 (
            .O(N__33511),
            .I(start_stop_c));
    InMux I__6358 (
            .O(N__33506),
            .I(N__33503));
    LocalMux I__6357 (
            .O(N__33503),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__6356 (
            .O(N__33500),
            .I(N__33497));
    LocalMux I__6355 (
            .O(N__33497),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__6354 (
            .O(N__33494),
            .I(N__33491));
    LocalMux I__6353 (
            .O(N__33491),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__6352 (
            .O(N__33488),
            .I(N__33485));
    LocalMux I__6351 (
            .O(N__33485),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__6350 (
            .O(N__33482),
            .I(N__33479));
    LocalMux I__6349 (
            .O(N__33479),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__6348 (
            .O(N__33476),
            .I(N__33473));
    LocalMux I__6347 (
            .O(N__33473),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__6346 (
            .O(N__33470),
            .I(N__33461));
    InMux I__6345 (
            .O(N__33469),
            .I(N__33461));
    InMux I__6344 (
            .O(N__33468),
            .I(N__33461));
    LocalMux I__6343 (
            .O(N__33461),
            .I(\phase_controller_inst1.tr_time_passed ));
    CascadeMux I__6342 (
            .O(N__33458),
            .I(N__33454));
    InMux I__6341 (
            .O(N__33457),
            .I(N__33450));
    InMux I__6340 (
            .O(N__33454),
            .I(N__33447));
    InMux I__6339 (
            .O(N__33453),
            .I(N__33444));
    LocalMux I__6338 (
            .O(N__33450),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__6337 (
            .O(N__33447),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__6336 (
            .O(N__33444),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    CascadeMux I__6335 (
            .O(N__33437),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_ ));
    InMux I__6334 (
            .O(N__33434),
            .I(N__33431));
    LocalMux I__6333 (
            .O(N__33431),
            .I(N__33428));
    Span4Mux_h I__6332 (
            .O(N__33428),
            .I(N__33424));
    InMux I__6331 (
            .O(N__33427),
            .I(N__33421));
    Odrv4 I__6330 (
            .O(N__33424),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    LocalMux I__6329 (
            .O(N__33421),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    CascadeMux I__6328 (
            .O(N__33416),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17_cascade_));
    CascadeMux I__6327 (
            .O(N__33413),
            .I(N__33408));
    InMux I__6326 (
            .O(N__33412),
            .I(N__33405));
    InMux I__6325 (
            .O(N__33411),
            .I(N__33400));
    InMux I__6324 (
            .O(N__33408),
            .I(N__33400));
    LocalMux I__6323 (
            .O(N__33405),
            .I(N__33396));
    LocalMux I__6322 (
            .O(N__33400),
            .I(N__33393));
    CascadeMux I__6321 (
            .O(N__33399),
            .I(N__33390));
    Span12Mux_v I__6320 (
            .O(N__33396),
            .I(N__33387));
    Span4Mux_h I__6319 (
            .O(N__33393),
            .I(N__33384));
    InMux I__6318 (
            .O(N__33390),
            .I(N__33381));
    Odrv12 I__6317 (
            .O(N__33387),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    Odrv4 I__6316 (
            .O(N__33384),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    LocalMux I__6315 (
            .O(N__33381),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    CascadeMux I__6314 (
            .O(N__33374),
            .I(N__33371));
    InMux I__6313 (
            .O(N__33371),
            .I(N__33368));
    LocalMux I__6312 (
            .O(N__33368),
            .I(N__33365));
    Span4Mux_h I__6311 (
            .O(N__33365),
            .I(N__33362));
    Odrv4 I__6310 (
            .O(N__33362),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    CascadeMux I__6309 (
            .O(N__33359),
            .I(N__33356));
    InMux I__6308 (
            .O(N__33356),
            .I(N__33349));
    InMux I__6307 (
            .O(N__33355),
            .I(N__33349));
    InMux I__6306 (
            .O(N__33354),
            .I(N__33346));
    LocalMux I__6305 (
            .O(N__33349),
            .I(N__33343));
    LocalMux I__6304 (
            .O(N__33346),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__6303 (
            .O(N__33343),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__6302 (
            .O(N__33338),
            .I(N__33335));
    InMux I__6301 (
            .O(N__33335),
            .I(N__33329));
    InMux I__6300 (
            .O(N__33334),
            .I(N__33329));
    LocalMux I__6299 (
            .O(N__33329),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__6298 (
            .O(N__33326),
            .I(N__33319));
    InMux I__6297 (
            .O(N__33325),
            .I(N__33319));
    InMux I__6296 (
            .O(N__33324),
            .I(N__33316));
    LocalMux I__6295 (
            .O(N__33319),
            .I(N__33313));
    LocalMux I__6294 (
            .O(N__33316),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv12 I__6293 (
            .O(N__33313),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__6292 (
            .O(N__33308),
            .I(N__33305));
    LocalMux I__6291 (
            .O(N__33305),
            .I(N__33302));
    Odrv4 I__6290 (
            .O(N__33302),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    InMux I__6289 (
            .O(N__33299),
            .I(N__33296));
    LocalMux I__6288 (
            .O(N__33296),
            .I(N__33293));
    Span4Mux_h I__6287 (
            .O(N__33293),
            .I(N__33289));
    InMux I__6286 (
            .O(N__33292),
            .I(N__33286));
    Odrv4 I__6285 (
            .O(N__33289),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    LocalMux I__6284 (
            .O(N__33286),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    InMux I__6283 (
            .O(N__33281),
            .I(N__33278));
    LocalMux I__6282 (
            .O(N__33278),
            .I(N__33273));
    InMux I__6281 (
            .O(N__33277),
            .I(N__33268));
    InMux I__6280 (
            .O(N__33276),
            .I(N__33268));
    Span4Mux_v I__6279 (
            .O(N__33273),
            .I(N__33264));
    LocalMux I__6278 (
            .O(N__33268),
            .I(N__33261));
    CascadeMux I__6277 (
            .O(N__33267),
            .I(N__33258));
    Span4Mux_v I__6276 (
            .O(N__33264),
            .I(N__33255));
    Span4Mux_v I__6275 (
            .O(N__33261),
            .I(N__33252));
    InMux I__6274 (
            .O(N__33258),
            .I(N__33249));
    Odrv4 I__6273 (
            .O(N__33255),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    Odrv4 I__6272 (
            .O(N__33252),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__6271 (
            .O(N__33249),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    CascadeMux I__6270 (
            .O(N__33242),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_));
    InMux I__6269 (
            .O(N__33239),
            .I(N__33233));
    InMux I__6268 (
            .O(N__33238),
            .I(N__33233));
    LocalMux I__6267 (
            .O(N__33233),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__6266 (
            .O(N__33230),
            .I(N__33227));
    LocalMux I__6265 (
            .O(N__33227),
            .I(N__33223));
    InMux I__6264 (
            .O(N__33226),
            .I(N__33220));
    Span4Mux_v I__6263 (
            .O(N__33223),
            .I(N__33217));
    LocalMux I__6262 (
            .O(N__33220),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    Odrv4 I__6261 (
            .O(N__33217),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__6260 (
            .O(N__33212),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__6259 (
            .O(N__33209),
            .I(N__33206));
    LocalMux I__6258 (
            .O(N__33206),
            .I(N__33203));
    Span4Mux_v I__6257 (
            .O(N__33203),
            .I(N__33200));
    Odrv4 I__6256 (
            .O(N__33200),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ));
    CascadeMux I__6255 (
            .O(N__33197),
            .I(N__33192));
    InMux I__6254 (
            .O(N__33196),
            .I(N__33189));
    InMux I__6253 (
            .O(N__33195),
            .I(N__33184));
    InMux I__6252 (
            .O(N__33192),
            .I(N__33184));
    LocalMux I__6251 (
            .O(N__33189),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__6250 (
            .O(N__33184),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__6249 (
            .O(N__33179),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    CascadeMux I__6248 (
            .O(N__33176),
            .I(N__33171));
    InMux I__6247 (
            .O(N__33175),
            .I(N__33168));
    InMux I__6246 (
            .O(N__33174),
            .I(N__33163));
    InMux I__6245 (
            .O(N__33171),
            .I(N__33163));
    LocalMux I__6244 (
            .O(N__33168),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__6243 (
            .O(N__33163),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__6242 (
            .O(N__33158),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__6241 (
            .O(N__33155),
            .I(N__33148));
    InMux I__6240 (
            .O(N__33154),
            .I(N__33148));
    InMux I__6239 (
            .O(N__33153),
            .I(N__33145));
    LocalMux I__6238 (
            .O(N__33148),
            .I(N__33142));
    LocalMux I__6237 (
            .O(N__33145),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__6236 (
            .O(N__33142),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__6235 (
            .O(N__33137),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__6234 (
            .O(N__33134),
            .I(N__33127));
    InMux I__6233 (
            .O(N__33133),
            .I(N__33127));
    InMux I__6232 (
            .O(N__33132),
            .I(N__33124));
    LocalMux I__6231 (
            .O(N__33127),
            .I(N__33121));
    LocalMux I__6230 (
            .O(N__33124),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__6229 (
            .O(N__33121),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__6228 (
            .O(N__33116),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    CascadeMux I__6227 (
            .O(N__33113),
            .I(N__33108));
    InMux I__6226 (
            .O(N__33112),
            .I(N__33105));
    InMux I__6225 (
            .O(N__33111),
            .I(N__33102));
    InMux I__6224 (
            .O(N__33108),
            .I(N__33099));
    LocalMux I__6223 (
            .O(N__33105),
            .I(N__33096));
    LocalMux I__6222 (
            .O(N__33102),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    LocalMux I__6221 (
            .O(N__33099),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__6220 (
            .O(N__33096),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__6219 (
            .O(N__33089),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__6218 (
            .O(N__33086),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    CascadeMux I__6217 (
            .O(N__33083),
            .I(N__33080));
    InMux I__6216 (
            .O(N__33080),
            .I(N__33075));
    InMux I__6215 (
            .O(N__33079),
            .I(N__33072));
    InMux I__6214 (
            .O(N__33078),
            .I(N__33069));
    LocalMux I__6213 (
            .O(N__33075),
            .I(N__33066));
    LocalMux I__6212 (
            .O(N__33072),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__6211 (
            .O(N__33069),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__6210 (
            .O(N__33066),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__6209 (
            .O(N__33059),
            .I(N__33056));
    LocalMux I__6208 (
            .O(N__33056),
            .I(N__33052));
    InMux I__6207 (
            .O(N__33055),
            .I(N__33049));
    Span4Mux_h I__6206 (
            .O(N__33052),
            .I(N__33046));
    LocalMux I__6205 (
            .O(N__33049),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    Odrv4 I__6204 (
            .O(N__33046),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    InMux I__6203 (
            .O(N__33041),
            .I(N__33038));
    LocalMux I__6202 (
            .O(N__33038),
            .I(N__33033));
    InMux I__6201 (
            .O(N__33037),
            .I(N__33028));
    InMux I__6200 (
            .O(N__33036),
            .I(N__33028));
    Span4Mux_h I__6199 (
            .O(N__33033),
            .I(N__33023));
    LocalMux I__6198 (
            .O(N__33028),
            .I(N__33023));
    Span4Mux_v I__6197 (
            .O(N__33023),
            .I(N__33019));
    InMux I__6196 (
            .O(N__33022),
            .I(N__33016));
    Odrv4 I__6195 (
            .O(N__33019),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__6194 (
            .O(N__33016),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    CascadeMux I__6193 (
            .O(N__33011),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_));
    CascadeMux I__6192 (
            .O(N__33008),
            .I(N__33005));
    InMux I__6191 (
            .O(N__33005),
            .I(N__33002));
    LocalMux I__6190 (
            .O(N__33002),
            .I(N__32999));
    Odrv4 I__6189 (
            .O(N__32999),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__6188 (
            .O(N__32996),
            .I(bfn_12_9_0_));
    CascadeMux I__6187 (
            .O(N__32993),
            .I(N__32989));
    CascadeMux I__6186 (
            .O(N__32992),
            .I(N__32986));
    InMux I__6185 (
            .O(N__32989),
            .I(N__32980));
    InMux I__6184 (
            .O(N__32986),
            .I(N__32980));
    InMux I__6183 (
            .O(N__32985),
            .I(N__32977));
    LocalMux I__6182 (
            .O(N__32980),
            .I(N__32974));
    LocalMux I__6181 (
            .O(N__32977),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv12 I__6180 (
            .O(N__32974),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__6179 (
            .O(N__32969),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__6178 (
            .O(N__32966),
            .I(N__32959));
    InMux I__6177 (
            .O(N__32965),
            .I(N__32959));
    InMux I__6176 (
            .O(N__32964),
            .I(N__32956));
    LocalMux I__6175 (
            .O(N__32959),
            .I(N__32953));
    LocalMux I__6174 (
            .O(N__32956),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__6173 (
            .O(N__32953),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__6172 (
            .O(N__32948),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    CascadeMux I__6171 (
            .O(N__32945),
            .I(N__32941));
    InMux I__6170 (
            .O(N__32944),
            .I(N__32935));
    InMux I__6169 (
            .O(N__32941),
            .I(N__32935));
    InMux I__6168 (
            .O(N__32940),
            .I(N__32932));
    LocalMux I__6167 (
            .O(N__32935),
            .I(N__32929));
    LocalMux I__6166 (
            .O(N__32932),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv12 I__6165 (
            .O(N__32929),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__6164 (
            .O(N__32924),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__6163 (
            .O(N__32921),
            .I(N__32914));
    InMux I__6162 (
            .O(N__32920),
            .I(N__32914));
    InMux I__6161 (
            .O(N__32919),
            .I(N__32911));
    LocalMux I__6160 (
            .O(N__32914),
            .I(N__32908));
    LocalMux I__6159 (
            .O(N__32911),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__6158 (
            .O(N__32908),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__6157 (
            .O(N__32903),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__6156 (
            .O(N__32900),
            .I(N__32893));
    InMux I__6155 (
            .O(N__32899),
            .I(N__32893));
    InMux I__6154 (
            .O(N__32898),
            .I(N__32890));
    LocalMux I__6153 (
            .O(N__32893),
            .I(N__32887));
    LocalMux I__6152 (
            .O(N__32890),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__6151 (
            .O(N__32887),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__6150 (
            .O(N__32882),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__6149 (
            .O(N__32879),
            .I(N__32872));
    InMux I__6148 (
            .O(N__32878),
            .I(N__32872));
    InMux I__6147 (
            .O(N__32877),
            .I(N__32869));
    LocalMux I__6146 (
            .O(N__32872),
            .I(N__32866));
    LocalMux I__6145 (
            .O(N__32869),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__6144 (
            .O(N__32866),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__6143 (
            .O(N__32861),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__6142 (
            .O(N__32858),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__6141 (
            .O(N__32855),
            .I(bfn_12_10_0_));
    InMux I__6140 (
            .O(N__32852),
            .I(N__32848));
    InMux I__6139 (
            .O(N__32851),
            .I(N__32845));
    LocalMux I__6138 (
            .O(N__32848),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__6137 (
            .O(N__32845),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__6136 (
            .O(N__32840),
            .I(bfn_12_8_0_));
    InMux I__6135 (
            .O(N__32837),
            .I(N__32833));
    InMux I__6134 (
            .O(N__32836),
            .I(N__32830));
    LocalMux I__6133 (
            .O(N__32833),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__6132 (
            .O(N__32830),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__6131 (
            .O(N__32825),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__6130 (
            .O(N__32822),
            .I(N__32818));
    InMux I__6129 (
            .O(N__32821),
            .I(N__32815));
    LocalMux I__6128 (
            .O(N__32818),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__6127 (
            .O(N__32815),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__6126 (
            .O(N__32810),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__6125 (
            .O(N__32807),
            .I(N__32803));
    InMux I__6124 (
            .O(N__32806),
            .I(N__32800));
    LocalMux I__6123 (
            .O(N__32803),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__6122 (
            .O(N__32800),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__6121 (
            .O(N__32795),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__6120 (
            .O(N__32792),
            .I(N__32788));
    InMux I__6119 (
            .O(N__32791),
            .I(N__32785));
    LocalMux I__6118 (
            .O(N__32788),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__6117 (
            .O(N__32785),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__6116 (
            .O(N__32780),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__6115 (
            .O(N__32777),
            .I(N__32773));
    InMux I__6114 (
            .O(N__32776),
            .I(N__32770));
    LocalMux I__6113 (
            .O(N__32773),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__6112 (
            .O(N__32770),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__6111 (
            .O(N__32765),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__6110 (
            .O(N__32762),
            .I(N__32758));
    InMux I__6109 (
            .O(N__32761),
            .I(N__32755));
    LocalMux I__6108 (
            .O(N__32758),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__6107 (
            .O(N__32755),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__6106 (
            .O(N__32750),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__6105 (
            .O(N__32747),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__6104 (
            .O(N__32744),
            .I(N__32741));
    LocalMux I__6103 (
            .O(N__32741),
            .I(N__32738));
    Span4Mux_h I__6102 (
            .O(N__32738),
            .I(N__32734));
    InMux I__6101 (
            .O(N__32737),
            .I(N__32730));
    Span4Mux_v I__6100 (
            .O(N__32734),
            .I(N__32727));
    InMux I__6099 (
            .O(N__32733),
            .I(N__32724));
    LocalMux I__6098 (
            .O(N__32730),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__6097 (
            .O(N__32727),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    LocalMux I__6096 (
            .O(N__32724),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__6095 (
            .O(N__32717),
            .I(N__32714));
    LocalMux I__6094 (
            .O(N__32714),
            .I(N__32709));
    InMux I__6093 (
            .O(N__32713),
            .I(N__32706));
    InMux I__6092 (
            .O(N__32712),
            .I(N__32703));
    Span4Mux_v I__6091 (
            .O(N__32709),
            .I(N__32700));
    LocalMux I__6090 (
            .O(N__32706),
            .I(N__32697));
    LocalMux I__6089 (
            .O(N__32703),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__6088 (
            .O(N__32700),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__6087 (
            .O(N__32697),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__6086 (
            .O(N__32690),
            .I(N__32687));
    InMux I__6085 (
            .O(N__32687),
            .I(N__32684));
    LocalMux I__6084 (
            .O(N__32684),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    InMux I__6083 (
            .O(N__32681),
            .I(N__32677));
    InMux I__6082 (
            .O(N__32680),
            .I(N__32674));
    LocalMux I__6081 (
            .O(N__32677),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__6080 (
            .O(N__32674),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__6079 (
            .O(N__32669),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__6078 (
            .O(N__32666),
            .I(N__32663));
    InMux I__6077 (
            .O(N__32663),
            .I(N__32659));
    InMux I__6076 (
            .O(N__32662),
            .I(N__32656));
    LocalMux I__6075 (
            .O(N__32659),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__6074 (
            .O(N__32656),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__6073 (
            .O(N__32651),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__6072 (
            .O(N__32648),
            .I(N__32644));
    InMux I__6071 (
            .O(N__32647),
            .I(N__32641));
    LocalMux I__6070 (
            .O(N__32644),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__6069 (
            .O(N__32641),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__6068 (
            .O(N__32636),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__6067 (
            .O(N__32633),
            .I(N__32629));
    InMux I__6066 (
            .O(N__32632),
            .I(N__32626));
    LocalMux I__6065 (
            .O(N__32629),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__6064 (
            .O(N__32626),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__6063 (
            .O(N__32621),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__6062 (
            .O(N__32618),
            .I(N__32614));
    InMux I__6061 (
            .O(N__32617),
            .I(N__32611));
    LocalMux I__6060 (
            .O(N__32614),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__6059 (
            .O(N__32611),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__6058 (
            .O(N__32606),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__6057 (
            .O(N__32603),
            .I(N__32599));
    InMux I__6056 (
            .O(N__32602),
            .I(N__32596));
    LocalMux I__6055 (
            .O(N__32599),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__6054 (
            .O(N__32596),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__6053 (
            .O(N__32591),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__6052 (
            .O(N__32588),
            .I(N__32584));
    InMux I__6051 (
            .O(N__32587),
            .I(N__32581));
    LocalMux I__6050 (
            .O(N__32584),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__6049 (
            .O(N__32581),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__6048 (
            .O(N__32576),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__6047 (
            .O(N__32573),
            .I(N__32570));
    LocalMux I__6046 (
            .O(N__32570),
            .I(N__32567));
    Odrv4 I__6045 (
            .O(N__32567),
            .I(\current_shift_inst.control_input_axb_18 ));
    InMux I__6044 (
            .O(N__32564),
            .I(N__32561));
    LocalMux I__6043 (
            .O(N__32561),
            .I(N__32558));
    Odrv4 I__6042 (
            .O(N__32558),
            .I(\current_shift_inst.control_input_axb_17 ));
    InMux I__6041 (
            .O(N__32555),
            .I(N__32552));
    LocalMux I__6040 (
            .O(N__32552),
            .I(N__32548));
    InMux I__6039 (
            .O(N__32551),
            .I(N__32545));
    Span4Mux_h I__6038 (
            .O(N__32548),
            .I(N__32542));
    LocalMux I__6037 (
            .O(N__32545),
            .I(N__32539));
    Sp12to4 I__6036 (
            .O(N__32542),
            .I(N__32536));
    Span12Mux_v I__6035 (
            .O(N__32539),
            .I(N__32533));
    Span12Mux_s6_v I__6034 (
            .O(N__32536),
            .I(N__32530));
    Span12Mux_h I__6033 (
            .O(N__32533),
            .I(N__32527));
    Odrv12 I__6032 (
            .O(N__32530),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    Odrv12 I__6031 (
            .O(N__32527),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    InMux I__6030 (
            .O(N__32522),
            .I(N__32518));
    InMux I__6029 (
            .O(N__32521),
            .I(N__32515));
    LocalMux I__6028 (
            .O(N__32518),
            .I(N__32510));
    LocalMux I__6027 (
            .O(N__32515),
            .I(N__32510));
    Span4Mux_h I__6026 (
            .O(N__32510),
            .I(N__32507));
    Span4Mux_v I__6025 (
            .O(N__32507),
            .I(N__32498));
    InMux I__6024 (
            .O(N__32506),
            .I(N__32491));
    InMux I__6023 (
            .O(N__32505),
            .I(N__32491));
    InMux I__6022 (
            .O(N__32504),
            .I(N__32491));
    InMux I__6021 (
            .O(N__32503),
            .I(N__32484));
    InMux I__6020 (
            .O(N__32502),
            .I(N__32484));
    InMux I__6019 (
            .O(N__32501),
            .I(N__32484));
    Sp12to4 I__6018 (
            .O(N__32498),
            .I(N__32477));
    LocalMux I__6017 (
            .O(N__32491),
            .I(N__32477));
    LocalMux I__6016 (
            .O(N__32484),
            .I(N__32477));
    Span12Mux_h I__6015 (
            .O(N__32477),
            .I(N__32474));
    Odrv12 I__6014 (
            .O(N__32474),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    InMux I__6013 (
            .O(N__32471),
            .I(N__32440));
    InMux I__6012 (
            .O(N__32470),
            .I(N__32440));
    InMux I__6011 (
            .O(N__32469),
            .I(N__32440));
    InMux I__6010 (
            .O(N__32468),
            .I(N__32440));
    InMux I__6009 (
            .O(N__32467),
            .I(N__32440));
    InMux I__6008 (
            .O(N__32466),
            .I(N__32440));
    InMux I__6007 (
            .O(N__32465),
            .I(N__32440));
    InMux I__6006 (
            .O(N__32464),
            .I(N__32440));
    InMux I__6005 (
            .O(N__32463),
            .I(N__32425));
    InMux I__6004 (
            .O(N__32462),
            .I(N__32425));
    InMux I__6003 (
            .O(N__32461),
            .I(N__32425));
    InMux I__6002 (
            .O(N__32460),
            .I(N__32425));
    InMux I__6001 (
            .O(N__32459),
            .I(N__32425));
    InMux I__6000 (
            .O(N__32458),
            .I(N__32425));
    InMux I__5999 (
            .O(N__32457),
            .I(N__32425));
    LocalMux I__5998 (
            .O(N__32440),
            .I(N__32418));
    LocalMux I__5997 (
            .O(N__32425),
            .I(N__32418));
    InMux I__5996 (
            .O(N__32424),
            .I(N__32415));
    InMux I__5995 (
            .O(N__32423),
            .I(N__32412));
    Span4Mux_s3_h I__5994 (
            .O(N__32418),
            .I(N__32403));
    LocalMux I__5993 (
            .O(N__32415),
            .I(N__32400));
    LocalMux I__5992 (
            .O(N__32412),
            .I(N__32397));
    CascadeMux I__5991 (
            .O(N__32411),
            .I(N__32386));
    InMux I__5990 (
            .O(N__32410),
            .I(N__32381));
    InMux I__5989 (
            .O(N__32409),
            .I(N__32381));
    InMux I__5988 (
            .O(N__32408),
            .I(N__32374));
    InMux I__5987 (
            .O(N__32407),
            .I(N__32374));
    InMux I__5986 (
            .O(N__32406),
            .I(N__32374));
    Span4Mux_h I__5985 (
            .O(N__32403),
            .I(N__32371));
    Span4Mux_v I__5984 (
            .O(N__32400),
            .I(N__32368));
    Span4Mux_v I__5983 (
            .O(N__32397),
            .I(N__32364));
    InMux I__5982 (
            .O(N__32396),
            .I(N__32347));
    InMux I__5981 (
            .O(N__32395),
            .I(N__32347));
    InMux I__5980 (
            .O(N__32394),
            .I(N__32347));
    InMux I__5979 (
            .O(N__32393),
            .I(N__32347));
    InMux I__5978 (
            .O(N__32392),
            .I(N__32347));
    InMux I__5977 (
            .O(N__32391),
            .I(N__32347));
    InMux I__5976 (
            .O(N__32390),
            .I(N__32347));
    InMux I__5975 (
            .O(N__32389),
            .I(N__32347));
    InMux I__5974 (
            .O(N__32386),
            .I(N__32344));
    LocalMux I__5973 (
            .O(N__32381),
            .I(N__32339));
    LocalMux I__5972 (
            .O(N__32374),
            .I(N__32339));
    Span4Mux_h I__5971 (
            .O(N__32371),
            .I(N__32336));
    Span4Mux_h I__5970 (
            .O(N__32368),
            .I(N__32333));
    InMux I__5969 (
            .O(N__32367),
            .I(N__32330));
    Sp12to4 I__5968 (
            .O(N__32364),
            .I(N__32321));
    LocalMux I__5967 (
            .O(N__32347),
            .I(N__32321));
    LocalMux I__5966 (
            .O(N__32344),
            .I(N__32321));
    Span12Mux_s7_v I__5965 (
            .O(N__32339),
            .I(N__32321));
    Span4Mux_h I__5964 (
            .O(N__32336),
            .I(N__32318));
    Odrv4 I__5963 (
            .O(N__32333),
            .I(N_19_1));
    LocalMux I__5962 (
            .O(N__32330),
            .I(N_19_1));
    Odrv12 I__5961 (
            .O(N__32321),
            .I(N_19_1));
    Odrv4 I__5960 (
            .O(N__32318),
            .I(N_19_1));
    InMux I__5959 (
            .O(N__32309),
            .I(N__32306));
    LocalMux I__5958 (
            .O(N__32306),
            .I(N__32303));
    Span4Mux_v I__5957 (
            .O(N__32303),
            .I(N__32300));
    Sp12to4 I__5956 (
            .O(N__32300),
            .I(N__32297));
    Span12Mux_h I__5955 (
            .O(N__32297),
            .I(N__32294));
    Odrv12 I__5954 (
            .O(N__32294),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__5953 (
            .O(N__32291),
            .I(N__32288));
    LocalMux I__5952 (
            .O(N__32288),
            .I(N__32285));
    Span4Mux_v I__5951 (
            .O(N__32285),
            .I(N__32282));
    Odrv4 I__5950 (
            .O(N__32282),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    InMux I__5949 (
            .O(N__32279),
            .I(N__32276));
    LocalMux I__5948 (
            .O(N__32276),
            .I(N__32273));
    Span4Mux_v I__5947 (
            .O(N__32273),
            .I(N__32270));
    Span4Mux_h I__5946 (
            .O(N__32270),
            .I(N__32267));
    Odrv4 I__5945 (
            .O(N__32267),
            .I(il_max_comp1_c));
    InMux I__5944 (
            .O(N__32264),
            .I(N__32261));
    LocalMux I__5943 (
            .O(N__32261),
            .I(il_max_comp1_D1));
    InMux I__5942 (
            .O(N__32258),
            .I(N__32254));
    InMux I__5941 (
            .O(N__32257),
            .I(N__32250));
    LocalMux I__5940 (
            .O(N__32254),
            .I(N__32247));
    InMux I__5939 (
            .O(N__32253),
            .I(N__32244));
    LocalMux I__5938 (
            .O(N__32250),
            .I(N__32240));
    Span4Mux_h I__5937 (
            .O(N__32247),
            .I(N__32235));
    LocalMux I__5936 (
            .O(N__32244),
            .I(N__32235));
    InMux I__5935 (
            .O(N__32243),
            .I(N__32232));
    Span4Mux_v I__5934 (
            .O(N__32240),
            .I(N__32229));
    Span4Mux_v I__5933 (
            .O(N__32235),
            .I(N__32226));
    LocalMux I__5932 (
            .O(N__32232),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__5931 (
            .O(N__32229),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__5930 (
            .O(N__32226),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    InMux I__5929 (
            .O(N__32219),
            .I(N__32216));
    LocalMux I__5928 (
            .O(N__32216),
            .I(N__32212));
    InMux I__5927 (
            .O(N__32215),
            .I(N__32209));
    Span4Mux_v I__5926 (
            .O(N__32212),
            .I(N__32205));
    LocalMux I__5925 (
            .O(N__32209),
            .I(N__32202));
    InMux I__5924 (
            .O(N__32208),
            .I(N__32199));
    Span4Mux_h I__5923 (
            .O(N__32205),
            .I(N__32196));
    Span4Mux_v I__5922 (
            .O(N__32202),
            .I(N__32193));
    LocalMux I__5921 (
            .O(N__32199),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__5920 (
            .O(N__32196),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__5919 (
            .O(N__32193),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    InMux I__5918 (
            .O(N__32186),
            .I(N__32183));
    LocalMux I__5917 (
            .O(N__32183),
            .I(N__32180));
    Span4Mux_v I__5916 (
            .O(N__32180),
            .I(N__32175));
    InMux I__5915 (
            .O(N__32179),
            .I(N__32172));
    InMux I__5914 (
            .O(N__32178),
            .I(N__32169));
    Span4Mux_v I__5913 (
            .O(N__32175),
            .I(N__32165));
    LocalMux I__5912 (
            .O(N__32172),
            .I(N__32160));
    LocalMux I__5911 (
            .O(N__32169),
            .I(N__32160));
    InMux I__5910 (
            .O(N__32168),
            .I(N__32157));
    Odrv4 I__5909 (
            .O(N__32165),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    Odrv12 I__5908 (
            .O(N__32160),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__5907 (
            .O(N__32157),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__5906 (
            .O(N__32150),
            .I(N__32147));
    LocalMux I__5905 (
            .O(N__32147),
            .I(N__32144));
    Odrv4 I__5904 (
            .O(N__32144),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ));
    InMux I__5903 (
            .O(N__32141),
            .I(bfn_11_18_0_));
    CascadeMux I__5902 (
            .O(N__32138),
            .I(N__32135));
    InMux I__5901 (
            .O(N__32135),
            .I(N__32132));
    LocalMux I__5900 (
            .O(N__32132),
            .I(N__32129));
    Odrv4 I__5899 (
            .O(N__32129),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ));
    InMux I__5898 (
            .O(N__32126),
            .I(\current_shift_inst.control_input_cry_24 ));
    InMux I__5897 (
            .O(N__32123),
            .I(N__32120));
    LocalMux I__5896 (
            .O(N__32120),
            .I(N__32117));
    Odrv4 I__5895 (
            .O(N__32117),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ));
    InMux I__5894 (
            .O(N__32114),
            .I(\current_shift_inst.control_input_cry_25 ));
    InMux I__5893 (
            .O(N__32111),
            .I(N__32108));
    LocalMux I__5892 (
            .O(N__32108),
            .I(N__32105));
    Odrv4 I__5891 (
            .O(N__32105),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ));
    InMux I__5890 (
            .O(N__32102),
            .I(\current_shift_inst.control_input_cry_26 ));
    CascadeMux I__5889 (
            .O(N__32099),
            .I(N__32096));
    InMux I__5888 (
            .O(N__32096),
            .I(N__32093));
    LocalMux I__5887 (
            .O(N__32093),
            .I(N__32090));
    Odrv4 I__5886 (
            .O(N__32090),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ));
    InMux I__5885 (
            .O(N__32087),
            .I(\current_shift_inst.control_input_cry_27 ));
    InMux I__5884 (
            .O(N__32084),
            .I(N__32081));
    LocalMux I__5883 (
            .O(N__32081),
            .I(N__32078));
    Odrv4 I__5882 (
            .O(N__32078),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ));
    InMux I__5881 (
            .O(N__32075),
            .I(\current_shift_inst.control_input_cry_28 ));
    InMux I__5880 (
            .O(N__32072),
            .I(\current_shift_inst.control_input_cry_29 ));
    InMux I__5879 (
            .O(N__32069),
            .I(N__32066));
    LocalMux I__5878 (
            .O(N__32066),
            .I(N__32062));
    InMux I__5877 (
            .O(N__32065),
            .I(N__32059));
    Odrv4 I__5876 (
            .O(N__32062),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__5875 (
            .O(N__32059),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__5874 (
            .O(N__32054),
            .I(N__32051));
    LocalMux I__5873 (
            .O(N__32051),
            .I(\current_shift_inst.control_input_axb_27 ));
    CascadeMux I__5872 (
            .O(N__32048),
            .I(N__32045));
    InMux I__5871 (
            .O(N__32045),
            .I(N__32042));
    LocalMux I__5870 (
            .O(N__32042),
            .I(N__32039));
    Odrv12 I__5869 (
            .O(N__32039),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ));
    InMux I__5868 (
            .O(N__32036),
            .I(bfn_11_17_0_));
    CascadeMux I__5867 (
            .O(N__32033),
            .I(N__32030));
    InMux I__5866 (
            .O(N__32030),
            .I(N__32027));
    LocalMux I__5865 (
            .O(N__32027),
            .I(N__32024));
    Odrv4 I__5864 (
            .O(N__32024),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ));
    InMux I__5863 (
            .O(N__32021),
            .I(\current_shift_inst.control_input_cry_16 ));
    InMux I__5862 (
            .O(N__32018),
            .I(N__32015));
    LocalMux I__5861 (
            .O(N__32015),
            .I(N__32012));
    Span4Mux_h I__5860 (
            .O(N__32012),
            .I(N__32009));
    Odrv4 I__5859 (
            .O(N__32009),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ));
    InMux I__5858 (
            .O(N__32006),
            .I(\current_shift_inst.control_input_cry_17 ));
    InMux I__5857 (
            .O(N__32003),
            .I(N__32000));
    LocalMux I__5856 (
            .O(N__32000),
            .I(\current_shift_inst.control_input_axb_19 ));
    InMux I__5855 (
            .O(N__31997),
            .I(N__31994));
    LocalMux I__5854 (
            .O(N__31994),
            .I(N__31991));
    Odrv4 I__5853 (
            .O(N__31991),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ));
    InMux I__5852 (
            .O(N__31988),
            .I(\current_shift_inst.control_input_cry_18 ));
    InMux I__5851 (
            .O(N__31985),
            .I(N__31982));
    LocalMux I__5850 (
            .O(N__31982),
            .I(N__31979));
    Odrv4 I__5849 (
            .O(N__31979),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ));
    InMux I__5848 (
            .O(N__31976),
            .I(\current_shift_inst.control_input_cry_19 ));
    InMux I__5847 (
            .O(N__31973),
            .I(N__31970));
    LocalMux I__5846 (
            .O(N__31970),
            .I(N__31967));
    Odrv4 I__5845 (
            .O(N__31967),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ));
    InMux I__5844 (
            .O(N__31964),
            .I(\current_shift_inst.control_input_cry_20 ));
    InMux I__5843 (
            .O(N__31961),
            .I(N__31958));
    LocalMux I__5842 (
            .O(N__31958),
            .I(N__31955));
    Odrv4 I__5841 (
            .O(N__31955),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ));
    InMux I__5840 (
            .O(N__31952),
            .I(\current_shift_inst.control_input_cry_21 ));
    CascadeMux I__5839 (
            .O(N__31949),
            .I(N__31946));
    InMux I__5838 (
            .O(N__31946),
            .I(N__31943));
    LocalMux I__5837 (
            .O(N__31943),
            .I(N__31940));
    Odrv4 I__5836 (
            .O(N__31940),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ));
    InMux I__5835 (
            .O(N__31937),
            .I(\current_shift_inst.control_input_cry_22 ));
    InMux I__5834 (
            .O(N__31934),
            .I(N__31931));
    LocalMux I__5833 (
            .O(N__31931),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__5832 (
            .O(N__31928),
            .I(N__31925));
    LocalMux I__5831 (
            .O(N__31925),
            .I(N__31922));
    Odrv4 I__5830 (
            .O(N__31922),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__5829 (
            .O(N__31919),
            .I(bfn_11_16_0_));
    InMux I__5828 (
            .O(N__31916),
            .I(N__31913));
    LocalMux I__5827 (
            .O(N__31913),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__5826 (
            .O(N__31910),
            .I(N__31907));
    LocalMux I__5825 (
            .O(N__31907),
            .I(N__31904));
    Odrv4 I__5824 (
            .O(N__31904),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__5823 (
            .O(N__31901),
            .I(\current_shift_inst.control_input_cry_8 ));
    CascadeMux I__5822 (
            .O(N__31898),
            .I(N__31895));
    InMux I__5821 (
            .O(N__31895),
            .I(N__31892));
    LocalMux I__5820 (
            .O(N__31892),
            .I(\current_shift_inst.control_input_axb_10 ));
    InMux I__5819 (
            .O(N__31889),
            .I(N__31886));
    LocalMux I__5818 (
            .O(N__31886),
            .I(N__31883));
    Span4Mux_h I__5817 (
            .O(N__31883),
            .I(N__31880));
    Odrv4 I__5816 (
            .O(N__31880),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__5815 (
            .O(N__31877),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__5814 (
            .O(N__31874),
            .I(N__31871));
    LocalMux I__5813 (
            .O(N__31871),
            .I(N__31868));
    Odrv4 I__5812 (
            .O(N__31868),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__5811 (
            .O(N__31865),
            .I(\current_shift_inst.control_input_cry_10 ));
    CascadeMux I__5810 (
            .O(N__31862),
            .I(N__31859));
    InMux I__5809 (
            .O(N__31859),
            .I(N__31856));
    LocalMux I__5808 (
            .O(N__31856),
            .I(N__31853));
    Odrv4 I__5807 (
            .O(N__31853),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__5806 (
            .O(N__31850),
            .I(\current_shift_inst.control_input_cry_11 ));
    CascadeMux I__5805 (
            .O(N__31847),
            .I(N__31844));
    InMux I__5804 (
            .O(N__31844),
            .I(N__31841));
    LocalMux I__5803 (
            .O(N__31841),
            .I(N__31838));
    Odrv4 I__5802 (
            .O(N__31838),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__5801 (
            .O(N__31835),
            .I(\current_shift_inst.control_input_cry_12 ));
    CascadeMux I__5800 (
            .O(N__31832),
            .I(N__31829));
    InMux I__5799 (
            .O(N__31829),
            .I(N__31826));
    LocalMux I__5798 (
            .O(N__31826),
            .I(N__31823));
    Odrv4 I__5797 (
            .O(N__31823),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ));
    InMux I__5796 (
            .O(N__31820),
            .I(\current_shift_inst.control_input_cry_13 ));
    CascadeMux I__5795 (
            .O(N__31817),
            .I(N__31814));
    InMux I__5794 (
            .O(N__31814),
            .I(N__31811));
    LocalMux I__5793 (
            .O(N__31811),
            .I(N__31808));
    Odrv4 I__5792 (
            .O(N__31808),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ));
    InMux I__5791 (
            .O(N__31805),
            .I(\current_shift_inst.control_input_cry_14 ));
    IoInMux I__5790 (
            .O(N__31802),
            .I(N__31799));
    LocalMux I__5789 (
            .O(N__31799),
            .I(N__31796));
    Span4Mux_s3_v I__5788 (
            .O(N__31796),
            .I(N__31793));
    Span4Mux_h I__5787 (
            .O(N__31793),
            .I(N__31790));
    Sp12to4 I__5786 (
            .O(N__31790),
            .I(N__31787));
    Span12Mux_v I__5785 (
            .O(N__31787),
            .I(N__31783));
    InMux I__5784 (
            .O(N__31786),
            .I(N__31780));
    Odrv12 I__5783 (
            .O(N__31783),
            .I(T45_c));
    LocalMux I__5782 (
            .O(N__31780),
            .I(T45_c));
    InMux I__5781 (
            .O(N__31775),
            .I(N__31772));
    LocalMux I__5780 (
            .O(N__31772),
            .I(\current_shift_inst.control_input_axb_0 ));
    CascadeMux I__5779 (
            .O(N__31769),
            .I(N__31764));
    InMux I__5778 (
            .O(N__31768),
            .I(N__31761));
    InMux I__5777 (
            .O(N__31767),
            .I(N__31758));
    InMux I__5776 (
            .O(N__31764),
            .I(N__31755));
    LocalMux I__5775 (
            .O(N__31761),
            .I(\current_shift_inst.N_1269_i ));
    LocalMux I__5774 (
            .O(N__31758),
            .I(\current_shift_inst.N_1269_i ));
    LocalMux I__5773 (
            .O(N__31755),
            .I(\current_shift_inst.N_1269_i ));
    InMux I__5772 (
            .O(N__31748),
            .I(N__31745));
    LocalMux I__5771 (
            .O(N__31745),
            .I(N__31742));
    Odrv4 I__5770 (
            .O(N__31742),
            .I(\current_shift_inst.control_input_1 ));
    InMux I__5769 (
            .O(N__31739),
            .I(N__31736));
    LocalMux I__5768 (
            .O(N__31736),
            .I(N__31733));
    Odrv4 I__5767 (
            .O(N__31733),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__5766 (
            .O(N__31730),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__5765 (
            .O(N__31727),
            .I(N__31724));
    LocalMux I__5764 (
            .O(N__31724),
            .I(N__31721));
    Odrv4 I__5763 (
            .O(N__31721),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__5762 (
            .O(N__31718),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__5761 (
            .O(N__31715),
            .I(N__31712));
    LocalMux I__5760 (
            .O(N__31712),
            .I(N__31709));
    Odrv4 I__5759 (
            .O(N__31709),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__5758 (
            .O(N__31706),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__5757 (
            .O(N__31703),
            .I(N__31700));
    LocalMux I__5756 (
            .O(N__31700),
            .I(N__31697));
    Odrv4 I__5755 (
            .O(N__31697),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__5754 (
            .O(N__31694),
            .I(\current_shift_inst.control_input_cry_3 ));
    CascadeMux I__5753 (
            .O(N__31691),
            .I(N__31688));
    InMux I__5752 (
            .O(N__31688),
            .I(N__31685));
    LocalMux I__5751 (
            .O(N__31685),
            .I(N__31682));
    Odrv4 I__5750 (
            .O(N__31682),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__5749 (
            .O(N__31679),
            .I(\current_shift_inst.control_input_cry_4 ));
    CascadeMux I__5748 (
            .O(N__31676),
            .I(N__31673));
    InMux I__5747 (
            .O(N__31673),
            .I(N__31670));
    LocalMux I__5746 (
            .O(N__31670),
            .I(N__31667));
    Odrv4 I__5745 (
            .O(N__31667),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__5744 (
            .O(N__31664),
            .I(\current_shift_inst.control_input_cry_5 ));
    CascadeMux I__5743 (
            .O(N__31661),
            .I(N__31658));
    InMux I__5742 (
            .O(N__31658),
            .I(N__31655));
    LocalMux I__5741 (
            .O(N__31655),
            .I(N__31652));
    Odrv4 I__5740 (
            .O(N__31652),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__5739 (
            .O(N__31649),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__5738 (
            .O(N__31646),
            .I(N__31642));
    InMux I__5737 (
            .O(N__31645),
            .I(N__31639));
    LocalMux I__5736 (
            .O(N__31642),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    LocalMux I__5735 (
            .O(N__31639),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    InMux I__5734 (
            .O(N__31634),
            .I(N__31630));
    InMux I__5733 (
            .O(N__31633),
            .I(N__31627));
    LocalMux I__5732 (
            .O(N__31630),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    LocalMux I__5731 (
            .O(N__31627),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    InMux I__5730 (
            .O(N__31622),
            .I(N__31619));
    LocalMux I__5729 (
            .O(N__31619),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ));
    CascadeMux I__5728 (
            .O(N__31616),
            .I(N__31611));
    CascadeMux I__5727 (
            .O(N__31615),
            .I(N__31608));
    InMux I__5726 (
            .O(N__31614),
            .I(N__31605));
    InMux I__5725 (
            .O(N__31611),
            .I(N__31599));
    InMux I__5724 (
            .O(N__31608),
            .I(N__31599));
    LocalMux I__5723 (
            .O(N__31605),
            .I(N__31596));
    InMux I__5722 (
            .O(N__31604),
            .I(N__31592));
    LocalMux I__5721 (
            .O(N__31599),
            .I(N__31587));
    Span4Mux_h I__5720 (
            .O(N__31596),
            .I(N__31587));
    InMux I__5719 (
            .O(N__31595),
            .I(N__31584));
    LocalMux I__5718 (
            .O(N__31592),
            .I(N__31581));
    Odrv4 I__5717 (
            .O(N__31587),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__5716 (
            .O(N__31584),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__5715 (
            .O(N__31581),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    InMux I__5714 (
            .O(N__31574),
            .I(N__31570));
    CascadeMux I__5713 (
            .O(N__31573),
            .I(N__31566));
    LocalMux I__5712 (
            .O(N__31570),
            .I(N__31562));
    InMux I__5711 (
            .O(N__31569),
            .I(N__31559));
    InMux I__5710 (
            .O(N__31566),
            .I(N__31554));
    InMux I__5709 (
            .O(N__31565),
            .I(N__31554));
    Span4Mux_v I__5708 (
            .O(N__31562),
            .I(N__31551));
    LocalMux I__5707 (
            .O(N__31559),
            .I(N__31548));
    LocalMux I__5706 (
            .O(N__31554),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__5705 (
            .O(N__31551),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__5704 (
            .O(N__31548),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    IoInMux I__5703 (
            .O(N__31541),
            .I(N__31516));
    InMux I__5702 (
            .O(N__31540),
            .I(N__31499));
    InMux I__5701 (
            .O(N__31539),
            .I(N__31499));
    InMux I__5700 (
            .O(N__31538),
            .I(N__31499));
    InMux I__5699 (
            .O(N__31537),
            .I(N__31499));
    InMux I__5698 (
            .O(N__31536),
            .I(N__31492));
    InMux I__5697 (
            .O(N__31535),
            .I(N__31492));
    InMux I__5696 (
            .O(N__31534),
            .I(N__31492));
    InMux I__5695 (
            .O(N__31533),
            .I(N__31483));
    InMux I__5694 (
            .O(N__31532),
            .I(N__31483));
    InMux I__5693 (
            .O(N__31531),
            .I(N__31483));
    InMux I__5692 (
            .O(N__31530),
            .I(N__31483));
    InMux I__5691 (
            .O(N__31529),
            .I(N__31476));
    InMux I__5690 (
            .O(N__31528),
            .I(N__31476));
    InMux I__5689 (
            .O(N__31527),
            .I(N__31476));
    InMux I__5688 (
            .O(N__31526),
            .I(N__31467));
    InMux I__5687 (
            .O(N__31525),
            .I(N__31467));
    InMux I__5686 (
            .O(N__31524),
            .I(N__31467));
    InMux I__5685 (
            .O(N__31523),
            .I(N__31467));
    InMux I__5684 (
            .O(N__31522),
            .I(N__31458));
    InMux I__5683 (
            .O(N__31521),
            .I(N__31458));
    InMux I__5682 (
            .O(N__31520),
            .I(N__31458));
    InMux I__5681 (
            .O(N__31519),
            .I(N__31458));
    LocalMux I__5680 (
            .O(N__31516),
            .I(N__31455));
    InMux I__5679 (
            .O(N__31515),
            .I(N__31446));
    InMux I__5678 (
            .O(N__31514),
            .I(N__31446));
    InMux I__5677 (
            .O(N__31513),
            .I(N__31446));
    InMux I__5676 (
            .O(N__31512),
            .I(N__31446));
    InMux I__5675 (
            .O(N__31511),
            .I(N__31437));
    InMux I__5674 (
            .O(N__31510),
            .I(N__31437));
    InMux I__5673 (
            .O(N__31509),
            .I(N__31437));
    InMux I__5672 (
            .O(N__31508),
            .I(N__31437));
    LocalMux I__5671 (
            .O(N__31499),
            .I(N__31430));
    LocalMux I__5670 (
            .O(N__31492),
            .I(N__31430));
    LocalMux I__5669 (
            .O(N__31483),
            .I(N__31430));
    LocalMux I__5668 (
            .O(N__31476),
            .I(N__31427));
    LocalMux I__5667 (
            .O(N__31467),
            .I(N__31424));
    LocalMux I__5666 (
            .O(N__31458),
            .I(N__31421));
    Span4Mux_s3_v I__5665 (
            .O(N__31455),
            .I(N__31418));
    LocalMux I__5664 (
            .O(N__31446),
            .I(N__31411));
    LocalMux I__5663 (
            .O(N__31437),
            .I(N__31411));
    Span4Mux_v I__5662 (
            .O(N__31430),
            .I(N__31411));
    Span4Mux_h I__5661 (
            .O(N__31427),
            .I(N__31406));
    Span4Mux_h I__5660 (
            .O(N__31424),
            .I(N__31406));
    Span4Mux_h I__5659 (
            .O(N__31421),
            .I(N__31403));
    Span4Mux_v I__5658 (
            .O(N__31418),
            .I(N__31400));
    Odrv4 I__5657 (
            .O(N__31411),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__5656 (
            .O(N__31406),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__5655 (
            .O(N__31403),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__5654 (
            .O(N__31400),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__5653 (
            .O(N__31391),
            .I(N__31386));
    InMux I__5652 (
            .O(N__31390),
            .I(N__31381));
    InMux I__5651 (
            .O(N__31389),
            .I(N__31381));
    LocalMux I__5650 (
            .O(N__31386),
            .I(N__31376));
    LocalMux I__5649 (
            .O(N__31381),
            .I(N__31373));
    InMux I__5648 (
            .O(N__31380),
            .I(N__31368));
    InMux I__5647 (
            .O(N__31379),
            .I(N__31368));
    Span4Mux_v I__5646 (
            .O(N__31376),
            .I(N__31365));
    Span4Mux_v I__5645 (
            .O(N__31373),
            .I(N__31362));
    LocalMux I__5644 (
            .O(N__31368),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    Odrv4 I__5643 (
            .O(N__31365),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    Odrv4 I__5642 (
            .O(N__31362),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__5641 (
            .O(N__31355),
            .I(N__31352));
    LocalMux I__5640 (
            .O(N__31352),
            .I(N__31347));
    InMux I__5639 (
            .O(N__31351),
            .I(N__31344));
    InMux I__5638 (
            .O(N__31350),
            .I(N__31341));
    Odrv12 I__5637 (
            .O(N__31347),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__5636 (
            .O(N__31344),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__5635 (
            .O(N__31341),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__5634 (
            .O(N__31334),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_ ));
    InMux I__5633 (
            .O(N__31331),
            .I(N__31328));
    LocalMux I__5632 (
            .O(N__31328),
            .I(N__31323));
    InMux I__5631 (
            .O(N__31327),
            .I(N__31320));
    InMux I__5630 (
            .O(N__31326),
            .I(N__31317));
    Span4Mux_v I__5629 (
            .O(N__31323),
            .I(N__31312));
    LocalMux I__5628 (
            .O(N__31320),
            .I(N__31312));
    LocalMux I__5627 (
            .O(N__31317),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__5626 (
            .O(N__31312),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__5625 (
            .O(N__31307),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ));
    InMux I__5624 (
            .O(N__31304),
            .I(N__31298));
    InMux I__5623 (
            .O(N__31303),
            .I(N__31298));
    LocalMux I__5622 (
            .O(N__31298),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__5621 (
            .O(N__31295),
            .I(N__31291));
    InMux I__5620 (
            .O(N__31294),
            .I(N__31287));
    LocalMux I__5619 (
            .O(N__31291),
            .I(N__31284));
    InMux I__5618 (
            .O(N__31290),
            .I(N__31281));
    LocalMux I__5617 (
            .O(N__31287),
            .I(N__31277));
    Span4Mux_v I__5616 (
            .O(N__31284),
            .I(N__31272));
    LocalMux I__5615 (
            .O(N__31281),
            .I(N__31272));
    InMux I__5614 (
            .O(N__31280),
            .I(N__31269));
    Span4Mux_v I__5613 (
            .O(N__31277),
            .I(N__31264));
    Span4Mux_h I__5612 (
            .O(N__31272),
            .I(N__31264));
    LocalMux I__5611 (
            .O(N__31269),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__5610 (
            .O(N__31264),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    CascadeMux I__5609 (
            .O(N__31259),
            .I(N__31256));
    InMux I__5608 (
            .O(N__31256),
            .I(N__31252));
    InMux I__5607 (
            .O(N__31255),
            .I(N__31249));
    LocalMux I__5606 (
            .O(N__31252),
            .I(N__31244));
    LocalMux I__5605 (
            .O(N__31249),
            .I(N__31244));
    Span4Mux_v I__5604 (
            .O(N__31244),
            .I(N__31238));
    InMux I__5603 (
            .O(N__31243),
            .I(N__31231));
    InMux I__5602 (
            .O(N__31242),
            .I(N__31231));
    InMux I__5601 (
            .O(N__31241),
            .I(N__31231));
    Odrv4 I__5600 (
            .O(N__31238),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__5599 (
            .O(N__31231),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    CascadeMux I__5598 (
            .O(N__31226),
            .I(N__31223));
    InMux I__5597 (
            .O(N__31223),
            .I(N__31220));
    LocalMux I__5596 (
            .O(N__31220),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    InMux I__5595 (
            .O(N__31217),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ));
    CascadeMux I__5594 (
            .O(N__31214),
            .I(N__31211));
    InMux I__5593 (
            .O(N__31211),
            .I(N__31208));
    LocalMux I__5592 (
            .O(N__31208),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt26 ));
    InMux I__5591 (
            .O(N__31205),
            .I(N__31202));
    LocalMux I__5590 (
            .O(N__31202),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ));
    InMux I__5589 (
            .O(N__31199),
            .I(N__31196));
    LocalMux I__5588 (
            .O(N__31196),
            .I(N__31193));
    Span4Mux_h I__5587 (
            .O(N__31193),
            .I(N__31189));
    InMux I__5586 (
            .O(N__31192),
            .I(N__31186));
    Odrv4 I__5585 (
            .O(N__31189),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    LocalMux I__5584 (
            .O(N__31186),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    CascadeMux I__5583 (
            .O(N__31181),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_));
    InMux I__5582 (
            .O(N__31178),
            .I(N__31175));
    LocalMux I__5581 (
            .O(N__31175),
            .I(N__31170));
    InMux I__5580 (
            .O(N__31174),
            .I(N__31165));
    InMux I__5579 (
            .O(N__31173),
            .I(N__31165));
    Span4Mux_v I__5578 (
            .O(N__31170),
            .I(N__31159));
    LocalMux I__5577 (
            .O(N__31165),
            .I(N__31159));
    InMux I__5576 (
            .O(N__31164),
            .I(N__31156));
    Span4Mux_h I__5575 (
            .O(N__31159),
            .I(N__31153));
    LocalMux I__5574 (
            .O(N__31156),
            .I(N__31150));
    Odrv4 I__5573 (
            .O(N__31153),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__5572 (
            .O(N__31150),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__5571 (
            .O(N__31145),
            .I(N__31139));
    InMux I__5570 (
            .O(N__31144),
            .I(N__31139));
    LocalMux I__5569 (
            .O(N__31139),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    InMux I__5568 (
            .O(N__31136),
            .I(N__31132));
    InMux I__5567 (
            .O(N__31135),
            .I(N__31129));
    LocalMux I__5566 (
            .O(N__31132),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    LocalMux I__5565 (
            .O(N__31129),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    CascadeMux I__5564 (
            .O(N__31124),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_));
    InMux I__5563 (
            .O(N__31121),
            .I(N__31116));
    InMux I__5562 (
            .O(N__31120),
            .I(N__31111));
    InMux I__5561 (
            .O(N__31119),
            .I(N__31111));
    LocalMux I__5560 (
            .O(N__31116),
            .I(N__31108));
    LocalMux I__5559 (
            .O(N__31111),
            .I(N__31105));
    Span4Mux_h I__5558 (
            .O(N__31108),
            .I(N__31101));
    Span4Mux_h I__5557 (
            .O(N__31105),
            .I(N__31098));
    InMux I__5556 (
            .O(N__31104),
            .I(N__31095));
    Odrv4 I__5555 (
            .O(N__31101),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv4 I__5554 (
            .O(N__31098),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    LocalMux I__5553 (
            .O(N__31095),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__5552 (
            .O(N__31088),
            .I(N__31082));
    InMux I__5551 (
            .O(N__31087),
            .I(N__31082));
    LocalMux I__5550 (
            .O(N__31082),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    CascadeMux I__5549 (
            .O(N__31079),
            .I(N__31076));
    InMux I__5548 (
            .O(N__31076),
            .I(N__31073));
    LocalMux I__5547 (
            .O(N__31073),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__5546 (
            .O(N__31070),
            .I(N__31067));
    LocalMux I__5545 (
            .O(N__31067),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__5544 (
            .O(N__31064),
            .I(N__31061));
    LocalMux I__5543 (
            .O(N__31061),
            .I(N__31058));
    Span4Mux_h I__5542 (
            .O(N__31058),
            .I(N__31055));
    Odrv4 I__5541 (
            .O(N__31055),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    CascadeMux I__5540 (
            .O(N__31052),
            .I(N__31049));
    InMux I__5539 (
            .O(N__31049),
            .I(N__31046));
    LocalMux I__5538 (
            .O(N__31046),
            .I(N__31043));
    Span4Mux_v I__5537 (
            .O(N__31043),
            .I(N__31040));
    Span4Mux_h I__5536 (
            .O(N__31040),
            .I(N__31037));
    Odrv4 I__5535 (
            .O(N__31037),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    InMux I__5534 (
            .O(N__31034),
            .I(N__31031));
    LocalMux I__5533 (
            .O(N__31031),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ));
    CascadeMux I__5532 (
            .O(N__31028),
            .I(N__31025));
    InMux I__5531 (
            .O(N__31025),
            .I(N__31022));
    LocalMux I__5530 (
            .O(N__31022),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt20 ));
    InMux I__5529 (
            .O(N__31019),
            .I(N__31016));
    LocalMux I__5528 (
            .O(N__31016),
            .I(N__31013));
    Odrv4 I__5527 (
            .O(N__31013),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ));
    CascadeMux I__5526 (
            .O(N__31010),
            .I(N__31007));
    InMux I__5525 (
            .O(N__31007),
            .I(N__31004));
    LocalMux I__5524 (
            .O(N__31004),
            .I(N__31001));
    Odrv12 I__5523 (
            .O(N__31001),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt22 ));
    InMux I__5522 (
            .O(N__30998),
            .I(N__30995));
    LocalMux I__5521 (
            .O(N__30995),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ));
    CascadeMux I__5520 (
            .O(N__30992),
            .I(N__30989));
    InMux I__5519 (
            .O(N__30989),
            .I(N__30986));
    LocalMux I__5518 (
            .O(N__30986),
            .I(N__30983));
    Odrv12 I__5517 (
            .O(N__30983),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt28 ));
    CascadeMux I__5516 (
            .O(N__30980),
            .I(N__30977));
    InMux I__5515 (
            .O(N__30977),
            .I(N__30974));
    LocalMux I__5514 (
            .O(N__30974),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__5513 (
            .O(N__30971),
            .I(N__30968));
    InMux I__5512 (
            .O(N__30968),
            .I(N__30965));
    LocalMux I__5511 (
            .O(N__30965),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__5510 (
            .O(N__30962),
            .I(N__30959));
    LocalMux I__5509 (
            .O(N__30959),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__5508 (
            .O(N__30956),
            .I(N__30953));
    InMux I__5507 (
            .O(N__30953),
            .I(N__30950));
    LocalMux I__5506 (
            .O(N__30950),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__5505 (
            .O(N__30947),
            .I(N__30944));
    LocalMux I__5504 (
            .O(N__30944),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__5503 (
            .O(N__30941),
            .I(N__30938));
    InMux I__5502 (
            .O(N__30938),
            .I(N__30935));
    LocalMux I__5501 (
            .O(N__30935),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__5500 (
            .O(N__30932),
            .I(N__30929));
    LocalMux I__5499 (
            .O(N__30929),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__5498 (
            .O(N__30926),
            .I(N__30923));
    InMux I__5497 (
            .O(N__30923),
            .I(N__30920));
    LocalMux I__5496 (
            .O(N__30920),
            .I(N__30917));
    Odrv4 I__5495 (
            .O(N__30917),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__5494 (
            .O(N__30914),
            .I(N__30911));
    LocalMux I__5493 (
            .O(N__30911),
            .I(N__30908));
    Odrv4 I__5492 (
            .O(N__30908),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__5491 (
            .O(N__30905),
            .I(N__30902));
    InMux I__5490 (
            .O(N__30902),
            .I(N__30899));
    LocalMux I__5489 (
            .O(N__30899),
            .I(N__30896));
    Odrv4 I__5488 (
            .O(N__30896),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__5487 (
            .O(N__30893),
            .I(N__30890));
    LocalMux I__5486 (
            .O(N__30890),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__5485 (
            .O(N__30887),
            .I(N__30884));
    LocalMux I__5484 (
            .O(N__30884),
            .I(N__30881));
    Odrv4 I__5483 (
            .O(N__30881),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__5482 (
            .O(N__30878),
            .I(N__30875));
    InMux I__5481 (
            .O(N__30875),
            .I(N__30872));
    LocalMux I__5480 (
            .O(N__30872),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__5479 (
            .O(N__30869),
            .I(N__30865));
    CascadeMux I__5478 (
            .O(N__30868),
            .I(N__30862));
    InMux I__5477 (
            .O(N__30865),
            .I(N__30857));
    InMux I__5476 (
            .O(N__30862),
            .I(N__30857));
    LocalMux I__5475 (
            .O(N__30857),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ));
    InMux I__5474 (
            .O(N__30854),
            .I(N__30848));
    InMux I__5473 (
            .O(N__30853),
            .I(N__30848));
    LocalMux I__5472 (
            .O(N__30848),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    InMux I__5471 (
            .O(N__30845),
            .I(N__30842));
    LocalMux I__5470 (
            .O(N__30842),
            .I(N__30839));
    Span4Mux_h I__5469 (
            .O(N__30839),
            .I(N__30835));
    InMux I__5468 (
            .O(N__30838),
            .I(N__30832));
    Span4Mux_v I__5467 (
            .O(N__30835),
            .I(N__30826));
    LocalMux I__5466 (
            .O(N__30832),
            .I(N__30826));
    InMux I__5465 (
            .O(N__30831),
            .I(N__30823));
    Span4Mux_h I__5464 (
            .O(N__30826),
            .I(N__30820));
    LocalMux I__5463 (
            .O(N__30823),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    Odrv4 I__5462 (
            .O(N__30820),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    InMux I__5461 (
            .O(N__30815),
            .I(N__30811));
    InMux I__5460 (
            .O(N__30814),
            .I(N__30808));
    LocalMux I__5459 (
            .O(N__30811),
            .I(N__30804));
    LocalMux I__5458 (
            .O(N__30808),
            .I(N__30801));
    CascadeMux I__5457 (
            .O(N__30807),
            .I(N__30797));
    Span4Mux_h I__5456 (
            .O(N__30804),
            .I(N__30792));
    Span4Mux_v I__5455 (
            .O(N__30801),
            .I(N__30792));
    InMux I__5454 (
            .O(N__30800),
            .I(N__30787));
    InMux I__5453 (
            .O(N__30797),
            .I(N__30787));
    Odrv4 I__5452 (
            .O(N__30792),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__5451 (
            .O(N__30787),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    CascadeMux I__5450 (
            .O(N__30782),
            .I(N__30779));
    InMux I__5449 (
            .O(N__30779),
            .I(N__30776));
    LocalMux I__5448 (
            .O(N__30776),
            .I(N__30773));
    Odrv4 I__5447 (
            .O(N__30773),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__5446 (
            .O(N__30770),
            .I(N__30767));
    LocalMux I__5445 (
            .O(N__30767),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__5444 (
            .O(N__30764),
            .I(N__30761));
    LocalMux I__5443 (
            .O(N__30761),
            .I(N__30758));
    Odrv12 I__5442 (
            .O(N__30758),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__5441 (
            .O(N__30755),
            .I(N__30752));
    InMux I__5440 (
            .O(N__30752),
            .I(N__30749));
    LocalMux I__5439 (
            .O(N__30749),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__5438 (
            .O(N__30746),
            .I(N__30743));
    LocalMux I__5437 (
            .O(N__30743),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__5436 (
            .O(N__30740),
            .I(N__30737));
    InMux I__5435 (
            .O(N__30737),
            .I(N__30734));
    LocalMux I__5434 (
            .O(N__30734),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__5433 (
            .O(N__30731),
            .I(N__30728));
    InMux I__5432 (
            .O(N__30728),
            .I(N__30725));
    LocalMux I__5431 (
            .O(N__30725),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__5430 (
            .O(N__30722),
            .I(N__30719));
    LocalMux I__5429 (
            .O(N__30719),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__5428 (
            .O(N__30716),
            .I(N__30713));
    LocalMux I__5427 (
            .O(N__30713),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__5426 (
            .O(N__30710),
            .I(N__30707));
    InMux I__5425 (
            .O(N__30707),
            .I(N__30704));
    LocalMux I__5424 (
            .O(N__30704),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__5423 (
            .O(N__30701),
            .I(N__30698));
    LocalMux I__5422 (
            .O(N__30698),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__5421 (
            .O(N__30695),
            .I(N__30692));
    InMux I__5420 (
            .O(N__30692),
            .I(N__30689));
    LocalMux I__5419 (
            .O(N__30689),
            .I(N__30686));
    Odrv4 I__5418 (
            .O(N__30686),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__5417 (
            .O(N__30683),
            .I(N__30680));
    InMux I__5416 (
            .O(N__30680),
            .I(N__30677));
    LocalMux I__5415 (
            .O(N__30677),
            .I(N__30674));
    Span4Mux_h I__5414 (
            .O(N__30674),
            .I(N__30671));
    Span4Mux_h I__5413 (
            .O(N__30671),
            .I(N__30668));
    Span4Mux_h I__5412 (
            .O(N__30668),
            .I(N__30665));
    Span4Mux_h I__5411 (
            .O(N__30665),
            .I(N__30662));
    Odrv4 I__5410 (
            .O(N__30662),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__5409 (
            .O(N__30659),
            .I(N__30656));
    LocalMux I__5408 (
            .O(N__30656),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ));
    InMux I__5407 (
            .O(N__30653),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    CascadeMux I__5406 (
            .O(N__30650),
            .I(N__30647));
    InMux I__5405 (
            .O(N__30647),
            .I(N__30644));
    LocalMux I__5404 (
            .O(N__30644),
            .I(N__30641));
    Span4Mux_v I__5403 (
            .O(N__30641),
            .I(N__30638));
    Sp12to4 I__5402 (
            .O(N__30638),
            .I(N__30635));
    Span12Mux_h I__5401 (
            .O(N__30635),
            .I(N__30632));
    Odrv12 I__5400 (
            .O(N__30632),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__5399 (
            .O(N__30629),
            .I(N__30626));
    LocalMux I__5398 (
            .O(N__30626),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ));
    InMux I__5397 (
            .O(N__30623),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    CascadeMux I__5396 (
            .O(N__30620),
            .I(N__30617));
    InMux I__5395 (
            .O(N__30617),
            .I(N__30614));
    LocalMux I__5394 (
            .O(N__30614),
            .I(N__30611));
    Span4Mux_v I__5393 (
            .O(N__30611),
            .I(N__30608));
    Sp12to4 I__5392 (
            .O(N__30608),
            .I(N__30605));
    Span12Mux_h I__5391 (
            .O(N__30605),
            .I(N__30602));
    Odrv12 I__5390 (
            .O(N__30602),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    InMux I__5389 (
            .O(N__30599),
            .I(N__30596));
    LocalMux I__5388 (
            .O(N__30596),
            .I(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ));
    InMux I__5387 (
            .O(N__30593),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    CascadeMux I__5386 (
            .O(N__30590),
            .I(N__30587));
    InMux I__5385 (
            .O(N__30587),
            .I(N__30584));
    LocalMux I__5384 (
            .O(N__30584),
            .I(N__30581));
    Span4Mux_v I__5383 (
            .O(N__30581),
            .I(N__30578));
    Span4Mux_h I__5382 (
            .O(N__30578),
            .I(N__30575));
    Sp12to4 I__5381 (
            .O(N__30575),
            .I(N__30572));
    Odrv12 I__5380 (
            .O(N__30572),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__5379 (
            .O(N__30569),
            .I(N__30566));
    LocalMux I__5378 (
            .O(N__30566),
            .I(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ));
    InMux I__5377 (
            .O(N__30563),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    CascadeMux I__5376 (
            .O(N__30560),
            .I(N__30557));
    InMux I__5375 (
            .O(N__30557),
            .I(N__30554));
    LocalMux I__5374 (
            .O(N__30554),
            .I(N__30551));
    Odrv12 I__5373 (
            .O(N__30551),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    InMux I__5372 (
            .O(N__30548),
            .I(N__30545));
    LocalMux I__5371 (
            .O(N__30545),
            .I(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ));
    InMux I__5370 (
            .O(N__30542),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__5369 (
            .O(N__30539),
            .I(N__30536));
    LocalMux I__5368 (
            .O(N__30536),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    InMux I__5367 (
            .O(N__30533),
            .I(bfn_10_28_0_));
    CascadeMux I__5366 (
            .O(N__30530),
            .I(N__30526));
    CascadeMux I__5365 (
            .O(N__30529),
            .I(N__30522));
    InMux I__5364 (
            .O(N__30526),
            .I(N__30516));
    InMux I__5363 (
            .O(N__30525),
            .I(N__30513));
    InMux I__5362 (
            .O(N__30522),
            .I(N__30510));
    CascadeMux I__5361 (
            .O(N__30521),
            .I(N__30507));
    CascadeMux I__5360 (
            .O(N__30520),
            .I(N__30504));
    InMux I__5359 (
            .O(N__30519),
            .I(N__30495));
    LocalMux I__5358 (
            .O(N__30516),
            .I(N__30492));
    LocalMux I__5357 (
            .O(N__30513),
            .I(N__30487));
    LocalMux I__5356 (
            .O(N__30510),
            .I(N__30487));
    InMux I__5355 (
            .O(N__30507),
            .I(N__30482));
    InMux I__5354 (
            .O(N__30504),
            .I(N__30482));
    InMux I__5353 (
            .O(N__30503),
            .I(N__30477));
    InMux I__5352 (
            .O(N__30502),
            .I(N__30477));
    InMux I__5351 (
            .O(N__30501),
            .I(N__30474));
    InMux I__5350 (
            .O(N__30500),
            .I(N__30471));
    InMux I__5349 (
            .O(N__30499),
            .I(N__30468));
    InMux I__5348 (
            .O(N__30498),
            .I(N__30465));
    LocalMux I__5347 (
            .O(N__30495),
            .I(N__30462));
    Span4Mux_v I__5346 (
            .O(N__30492),
            .I(N__30457));
    Span4Mux_v I__5345 (
            .O(N__30487),
            .I(N__30457));
    LocalMux I__5344 (
            .O(N__30482),
            .I(N__30454));
    LocalMux I__5343 (
            .O(N__30477),
            .I(N__30449));
    LocalMux I__5342 (
            .O(N__30474),
            .I(N__30449));
    LocalMux I__5341 (
            .O(N__30471),
            .I(N__30440));
    LocalMux I__5340 (
            .O(N__30468),
            .I(N__30440));
    LocalMux I__5339 (
            .O(N__30465),
            .I(N__30440));
    Span4Mux_s2_h I__5338 (
            .O(N__30462),
            .I(N__30440));
    Span4Mux_h I__5337 (
            .O(N__30457),
            .I(N__30437));
    Span4Mux_h I__5336 (
            .O(N__30454),
            .I(N__30432));
    Span4Mux_h I__5335 (
            .O(N__30449),
            .I(N__30432));
    Span4Mux_h I__5334 (
            .O(N__30440),
            .I(N__30429));
    Span4Mux_h I__5333 (
            .O(N__30437),
            .I(N__30426));
    Span4Mux_h I__5332 (
            .O(N__30432),
            .I(N__30423));
    Span4Mux_h I__5331 (
            .O(N__30429),
            .I(N__30420));
    Odrv4 I__5330 (
            .O(N__30426),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__5329 (
            .O(N__30423),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__5328 (
            .O(N__30420),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    InMux I__5327 (
            .O(N__30413),
            .I(N__30410));
    LocalMux I__5326 (
            .O(N__30410),
            .I(N__30407));
    Span4Mux_v I__5325 (
            .O(N__30407),
            .I(N__30404));
    Sp12to4 I__5324 (
            .O(N__30404),
            .I(N__30401));
    Span12Mux_h I__5323 (
            .O(N__30401),
            .I(N__30398));
    Odrv12 I__5322 (
            .O(N__30398),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    CascadeMux I__5321 (
            .O(N__30395),
            .I(N__30392));
    InMux I__5320 (
            .O(N__30392),
            .I(N__30389));
    LocalMux I__5319 (
            .O(N__30389),
            .I(N__30386));
    Span4Mux_h I__5318 (
            .O(N__30386),
            .I(N__30383));
    Span4Mux_h I__5317 (
            .O(N__30383),
            .I(N__30380));
    Span4Mux_h I__5316 (
            .O(N__30380),
            .I(N__30377));
    Odrv4 I__5315 (
            .O(N__30377),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    InMux I__5314 (
            .O(N__30374),
            .I(N__30371));
    LocalMux I__5313 (
            .O(N__30371),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ));
    InMux I__5312 (
            .O(N__30368),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__5311 (
            .O(N__30365),
            .I(N__30362));
    LocalMux I__5310 (
            .O(N__30362),
            .I(N__30359));
    Span4Mux_v I__5309 (
            .O(N__30359),
            .I(N__30356));
    Sp12to4 I__5308 (
            .O(N__30356),
            .I(N__30353));
    Span12Mux_h I__5307 (
            .O(N__30353),
            .I(N__30350));
    Odrv12 I__5306 (
            .O(N__30350),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__5305 (
            .O(N__30347),
            .I(N__30344));
    InMux I__5304 (
            .O(N__30344),
            .I(N__30341));
    LocalMux I__5303 (
            .O(N__30341),
            .I(N__30338));
    Span4Mux_v I__5302 (
            .O(N__30338),
            .I(N__30335));
    Sp12to4 I__5301 (
            .O(N__30335),
            .I(N__30332));
    Odrv12 I__5300 (
            .O(N__30332),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    InMux I__5299 (
            .O(N__30329),
            .I(N__30326));
    LocalMux I__5298 (
            .O(N__30326),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ));
    InMux I__5297 (
            .O(N__30323),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__5296 (
            .O(N__30320),
            .I(N__30317));
    LocalMux I__5295 (
            .O(N__30317),
            .I(N__30314));
    Span4Mux_v I__5294 (
            .O(N__30314),
            .I(N__30311));
    Sp12to4 I__5293 (
            .O(N__30311),
            .I(N__30308));
    Span12Mux_h I__5292 (
            .O(N__30308),
            .I(N__30305));
    Odrv12 I__5291 (
            .O(N__30305),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    CascadeMux I__5290 (
            .O(N__30302),
            .I(N__30299));
    InMux I__5289 (
            .O(N__30299),
            .I(N__30296));
    LocalMux I__5288 (
            .O(N__30296),
            .I(N__30293));
    Sp12to4 I__5287 (
            .O(N__30293),
            .I(N__30290));
    Span12Mux_s5_v I__5286 (
            .O(N__30290),
            .I(N__30287));
    Odrv12 I__5285 (
            .O(N__30287),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    InMux I__5284 (
            .O(N__30284),
            .I(N__30281));
    LocalMux I__5283 (
            .O(N__30281),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ));
    InMux I__5282 (
            .O(N__30278),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__5281 (
            .O(N__30275),
            .I(N__30272));
    LocalMux I__5280 (
            .O(N__30272),
            .I(N__30269));
    Span12Mux_s7_v I__5279 (
            .O(N__30269),
            .I(N__30266));
    Span12Mux_h I__5278 (
            .O(N__30266),
            .I(N__30263));
    Odrv12 I__5277 (
            .O(N__30263),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    CascadeMux I__5276 (
            .O(N__30260),
            .I(N__30257));
    InMux I__5275 (
            .O(N__30257),
            .I(N__30254));
    LocalMux I__5274 (
            .O(N__30254),
            .I(N__30251));
    Sp12to4 I__5273 (
            .O(N__30251),
            .I(N__30248));
    Span12Mux_s5_v I__5272 (
            .O(N__30248),
            .I(N__30245));
    Odrv12 I__5271 (
            .O(N__30245),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    InMux I__5270 (
            .O(N__30242),
            .I(N__30239));
    LocalMux I__5269 (
            .O(N__30239),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ));
    InMux I__5268 (
            .O(N__30236),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__5267 (
            .O(N__30233),
            .I(N__30230));
    LocalMux I__5266 (
            .O(N__30230),
            .I(N__30227));
    Span4Mux_v I__5265 (
            .O(N__30227),
            .I(N__30224));
    Sp12to4 I__5264 (
            .O(N__30224),
            .I(N__30221));
    Odrv12 I__5263 (
            .O(N__30221),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    CascadeMux I__5262 (
            .O(N__30218),
            .I(N__30215));
    InMux I__5261 (
            .O(N__30215),
            .I(N__30212));
    LocalMux I__5260 (
            .O(N__30212),
            .I(N__30209));
    Span4Mux_v I__5259 (
            .O(N__30209),
            .I(N__30206));
    Sp12to4 I__5258 (
            .O(N__30206),
            .I(N__30203));
    Span12Mux_h I__5257 (
            .O(N__30203),
            .I(N__30200));
    Odrv12 I__5256 (
            .O(N__30200),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    InMux I__5255 (
            .O(N__30197),
            .I(N__30194));
    LocalMux I__5254 (
            .O(N__30194),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ));
    InMux I__5253 (
            .O(N__30191),
            .I(bfn_10_27_0_));
    InMux I__5252 (
            .O(N__30188),
            .I(N__30185));
    LocalMux I__5251 (
            .O(N__30185),
            .I(N__30182));
    Span4Mux_h I__5250 (
            .O(N__30182),
            .I(N__30179));
    Span4Mux_h I__5249 (
            .O(N__30179),
            .I(N__30176));
    Span4Mux_h I__5248 (
            .O(N__30176),
            .I(N__30173));
    Odrv4 I__5247 (
            .O(N__30173),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    CascadeMux I__5246 (
            .O(N__30170),
            .I(N__30167));
    InMux I__5245 (
            .O(N__30167),
            .I(N__30164));
    LocalMux I__5244 (
            .O(N__30164),
            .I(N__30161));
    Span4Mux_v I__5243 (
            .O(N__30161),
            .I(N__30158));
    Span4Mux_h I__5242 (
            .O(N__30158),
            .I(N__30155));
    Span4Mux_h I__5241 (
            .O(N__30155),
            .I(N__30152));
    Span4Mux_h I__5240 (
            .O(N__30152),
            .I(N__30149));
    Odrv4 I__5239 (
            .O(N__30149),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    InMux I__5238 (
            .O(N__30146),
            .I(N__30143));
    LocalMux I__5237 (
            .O(N__30143),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ));
    InMux I__5236 (
            .O(N__30140),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    CascadeMux I__5235 (
            .O(N__30137),
            .I(N__30134));
    InMux I__5234 (
            .O(N__30134),
            .I(N__30131));
    LocalMux I__5233 (
            .O(N__30131),
            .I(N__30128));
    Span4Mux_v I__5232 (
            .O(N__30128),
            .I(N__30125));
    Sp12to4 I__5231 (
            .O(N__30125),
            .I(N__30122));
    Span12Mux_h I__5230 (
            .O(N__30122),
            .I(N__30119));
    Odrv12 I__5229 (
            .O(N__30119),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__5228 (
            .O(N__30116),
            .I(N__30113));
    LocalMux I__5227 (
            .O(N__30113),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ));
    InMux I__5226 (
            .O(N__30110),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    InMux I__5225 (
            .O(N__30107),
            .I(N__30104));
    LocalMux I__5224 (
            .O(N__30104),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ));
    InMux I__5223 (
            .O(N__30101),
            .I(N__30098));
    LocalMux I__5222 (
            .O(N__30098),
            .I(N__30095));
    Span4Mux_v I__5221 (
            .O(N__30095),
            .I(N__30092));
    Sp12to4 I__5220 (
            .O(N__30092),
            .I(N__30089));
    Span12Mux_h I__5219 (
            .O(N__30089),
            .I(N__30086));
    Odrv12 I__5218 (
            .O(N__30086),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__5217 (
            .O(N__30083),
            .I(N__30080));
    InMux I__5216 (
            .O(N__30080),
            .I(N__30077));
    LocalMux I__5215 (
            .O(N__30077),
            .I(N__30074));
    Span4Mux_h I__5214 (
            .O(N__30074),
            .I(N__30071));
    Span4Mux_h I__5213 (
            .O(N__30071),
            .I(N__30068));
    Span4Mux_h I__5212 (
            .O(N__30068),
            .I(N__30065));
    Odrv4 I__5211 (
            .O(N__30065),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__5210 (
            .O(N__30062),
            .I(N__30059));
    LocalMux I__5209 (
            .O(N__30059),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    InMux I__5208 (
            .O(N__30056),
            .I(N__30053));
    LocalMux I__5207 (
            .O(N__30053),
            .I(N__30050));
    Span4Mux_v I__5206 (
            .O(N__30050),
            .I(N__30047));
    Sp12to4 I__5205 (
            .O(N__30047),
            .I(N__30044));
    Span12Mux_h I__5204 (
            .O(N__30044),
            .I(N__30041));
    Odrv12 I__5203 (
            .O(N__30041),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__5202 (
            .O(N__30038),
            .I(N__30035));
    InMux I__5201 (
            .O(N__30035),
            .I(N__30032));
    LocalMux I__5200 (
            .O(N__30032),
            .I(N__30029));
    Span4Mux_h I__5199 (
            .O(N__30029),
            .I(N__30026));
    Span4Mux_h I__5198 (
            .O(N__30026),
            .I(N__30023));
    Span4Mux_h I__5197 (
            .O(N__30023),
            .I(N__30020));
    Odrv4 I__5196 (
            .O(N__30020),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    CascadeMux I__5195 (
            .O(N__30017),
            .I(N__30014));
    InMux I__5194 (
            .O(N__30014),
            .I(N__30011));
    LocalMux I__5193 (
            .O(N__30011),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ));
    InMux I__5192 (
            .O(N__30008),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__5191 (
            .O(N__30005),
            .I(N__30002));
    LocalMux I__5190 (
            .O(N__30002),
            .I(N__29999));
    Span4Mux_v I__5189 (
            .O(N__29999),
            .I(N__29996));
    Sp12to4 I__5188 (
            .O(N__29996),
            .I(N__29993));
    Span12Mux_h I__5187 (
            .O(N__29993),
            .I(N__29990));
    Odrv12 I__5186 (
            .O(N__29990),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__5185 (
            .O(N__29987),
            .I(N__29984));
    InMux I__5184 (
            .O(N__29984),
            .I(N__29981));
    LocalMux I__5183 (
            .O(N__29981),
            .I(N__29978));
    Span4Mux_h I__5182 (
            .O(N__29978),
            .I(N__29975));
    Span4Mux_h I__5181 (
            .O(N__29975),
            .I(N__29972));
    Span4Mux_h I__5180 (
            .O(N__29972),
            .I(N__29969));
    Odrv4 I__5179 (
            .O(N__29969),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    InMux I__5178 (
            .O(N__29966),
            .I(N__29963));
    LocalMux I__5177 (
            .O(N__29963),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ));
    InMux I__5176 (
            .O(N__29960),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__5175 (
            .O(N__29957),
            .I(N__29954));
    LocalMux I__5174 (
            .O(N__29954),
            .I(N__29951));
    Span12Mux_h I__5173 (
            .O(N__29951),
            .I(N__29948));
    Span12Mux_h I__5172 (
            .O(N__29948),
            .I(N__29945));
    Odrv12 I__5171 (
            .O(N__29945),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__5170 (
            .O(N__29942),
            .I(N__29939));
    InMux I__5169 (
            .O(N__29939),
            .I(N__29936));
    LocalMux I__5168 (
            .O(N__29936),
            .I(N__29933));
    Span4Mux_h I__5167 (
            .O(N__29933),
            .I(N__29930));
    Span4Mux_h I__5166 (
            .O(N__29930),
            .I(N__29927));
    Span4Mux_h I__5165 (
            .O(N__29927),
            .I(N__29924));
    Odrv4 I__5164 (
            .O(N__29924),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    CascadeMux I__5163 (
            .O(N__29921),
            .I(N__29918));
    InMux I__5162 (
            .O(N__29918),
            .I(N__29915));
    LocalMux I__5161 (
            .O(N__29915),
            .I(N__29912));
    Odrv4 I__5160 (
            .O(N__29912),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ));
    InMux I__5159 (
            .O(N__29909),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    CascadeMux I__5158 (
            .O(N__29906),
            .I(N__29903));
    InMux I__5157 (
            .O(N__29903),
            .I(N__29900));
    LocalMux I__5156 (
            .O(N__29900),
            .I(N__29897));
    Odrv4 I__5155 (
            .O(N__29897),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    InMux I__5154 (
            .O(N__29894),
            .I(N__29888));
    InMux I__5153 (
            .O(N__29893),
            .I(N__29888));
    LocalMux I__5152 (
            .O(N__29888),
            .I(N__29884));
    InMux I__5151 (
            .O(N__29887),
            .I(N__29881));
    Span4Mux_h I__5150 (
            .O(N__29884),
            .I(N__29878));
    LocalMux I__5149 (
            .O(N__29881),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__5148 (
            .O(N__29878),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__5147 (
            .O(N__29873),
            .I(N__29870));
    InMux I__5146 (
            .O(N__29870),
            .I(N__29864));
    InMux I__5145 (
            .O(N__29869),
            .I(N__29864));
    LocalMux I__5144 (
            .O(N__29864),
            .I(N__29860));
    InMux I__5143 (
            .O(N__29863),
            .I(N__29857));
    Span4Mux_h I__5142 (
            .O(N__29860),
            .I(N__29854));
    LocalMux I__5141 (
            .O(N__29857),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__5140 (
            .O(N__29854),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__5139 (
            .O(N__29849),
            .I(N__29846));
    LocalMux I__5138 (
            .O(N__29846),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    InMux I__5137 (
            .O(N__29843),
            .I(N__29837));
    InMux I__5136 (
            .O(N__29842),
            .I(N__29837));
    LocalMux I__5135 (
            .O(N__29837),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__5134 (
            .O(N__29834),
            .I(N__29831));
    InMux I__5133 (
            .O(N__29831),
            .I(N__29825));
    InMux I__5132 (
            .O(N__29830),
            .I(N__29825));
    LocalMux I__5131 (
            .O(N__29825),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    InMux I__5130 (
            .O(N__29822),
            .I(N__29819));
    LocalMux I__5129 (
            .O(N__29819),
            .I(N__29814));
    InMux I__5128 (
            .O(N__29818),
            .I(N__29809));
    InMux I__5127 (
            .O(N__29817),
            .I(N__29809));
    Span4Mux_v I__5126 (
            .O(N__29814),
            .I(N__29804));
    LocalMux I__5125 (
            .O(N__29809),
            .I(N__29804));
    Span4Mux_v I__5124 (
            .O(N__29804),
            .I(N__29800));
    InMux I__5123 (
            .O(N__29803),
            .I(N__29797));
    Odrv4 I__5122 (
            .O(N__29800),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    LocalMux I__5121 (
            .O(N__29797),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    InMux I__5120 (
            .O(N__29792),
            .I(N__29789));
    LocalMux I__5119 (
            .O(N__29789),
            .I(N__29785));
    InMux I__5118 (
            .O(N__29788),
            .I(N__29782));
    Odrv12 I__5117 (
            .O(N__29785),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    LocalMux I__5116 (
            .O(N__29782),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    CascadeMux I__5115 (
            .O(N__29777),
            .I(N__29774));
    InMux I__5114 (
            .O(N__29774),
            .I(N__29771));
    LocalMux I__5113 (
            .O(N__29771),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    CEMux I__5112 (
            .O(N__29768),
            .I(N__29735));
    CEMux I__5111 (
            .O(N__29767),
            .I(N__29735));
    CEMux I__5110 (
            .O(N__29766),
            .I(N__29735));
    CEMux I__5109 (
            .O(N__29765),
            .I(N__29735));
    CEMux I__5108 (
            .O(N__29764),
            .I(N__29735));
    CEMux I__5107 (
            .O(N__29763),
            .I(N__29735));
    CEMux I__5106 (
            .O(N__29762),
            .I(N__29735));
    CEMux I__5105 (
            .O(N__29761),
            .I(N__29735));
    CEMux I__5104 (
            .O(N__29760),
            .I(N__29735));
    CEMux I__5103 (
            .O(N__29759),
            .I(N__29735));
    CEMux I__5102 (
            .O(N__29758),
            .I(N__29735));
    GlobalMux I__5101 (
            .O(N__29735),
            .I(N__29732));
    gio2CtrlBuf I__5100 (
            .O(N__29732),
            .I(\phase_controller_inst2.stoper_tr.un1_start_g ));
    CascadeMux I__5099 (
            .O(N__29729),
            .I(\current_shift_inst.control_input_axb_0_cascade_ ));
    InMux I__5098 (
            .O(N__29726),
            .I(N__29722));
    InMux I__5097 (
            .O(N__29725),
            .I(N__29719));
    LocalMux I__5096 (
            .O(N__29722),
            .I(N__29716));
    LocalMux I__5095 (
            .O(N__29719),
            .I(N__29713));
    Span4Mux_s2_h I__5094 (
            .O(N__29716),
            .I(N__29710));
    Span4Mux_v I__5093 (
            .O(N__29713),
            .I(N__29707));
    Span4Mux_h I__5092 (
            .O(N__29710),
            .I(N__29704));
    Span4Mux_h I__5091 (
            .O(N__29707),
            .I(N__29701));
    Span4Mux_h I__5090 (
            .O(N__29704),
            .I(N__29698));
    Odrv4 I__5089 (
            .O(N__29701),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    Odrv4 I__5088 (
            .O(N__29698),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__5087 (
            .O(N__29693),
            .I(N__29690));
    LocalMux I__5086 (
            .O(N__29690),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    InMux I__5085 (
            .O(N__29687),
            .I(N__29684));
    LocalMux I__5084 (
            .O(N__29684),
            .I(N__29681));
    Span4Mux_h I__5083 (
            .O(N__29681),
            .I(N__29675));
    InMux I__5082 (
            .O(N__29680),
            .I(N__29668));
    InMux I__5081 (
            .O(N__29679),
            .I(N__29668));
    InMux I__5080 (
            .O(N__29678),
            .I(N__29668));
    Odrv4 I__5079 (
            .O(N__29675),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    LocalMux I__5078 (
            .O(N__29668),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__5077 (
            .O(N__29663),
            .I(N__29660));
    LocalMux I__5076 (
            .O(N__29660),
            .I(N__29657));
    Span4Mux_v I__5075 (
            .O(N__29657),
            .I(N__29653));
    InMux I__5074 (
            .O(N__29656),
            .I(N__29650));
    Odrv4 I__5073 (
            .O(N__29653),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    LocalMux I__5072 (
            .O(N__29650),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    InMux I__5071 (
            .O(N__29645),
            .I(N__29642));
    LocalMux I__5070 (
            .O(N__29642),
            .I(N__29637));
    InMux I__5069 (
            .O(N__29641),
            .I(N__29632));
    InMux I__5068 (
            .O(N__29640),
            .I(N__29632));
    Span4Mux_v I__5067 (
            .O(N__29637),
            .I(N__29628));
    LocalMux I__5066 (
            .O(N__29632),
            .I(N__29625));
    InMux I__5065 (
            .O(N__29631),
            .I(N__29622));
    Odrv4 I__5064 (
            .O(N__29628),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv12 I__5063 (
            .O(N__29625),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    LocalMux I__5062 (
            .O(N__29622),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__5061 (
            .O(N__29615),
            .I(N__29612));
    LocalMux I__5060 (
            .O(N__29612),
            .I(N__29608));
    InMux I__5059 (
            .O(N__29611),
            .I(N__29605));
    Odrv12 I__5058 (
            .O(N__29608),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    LocalMux I__5057 (
            .O(N__29605),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    InMux I__5056 (
            .O(N__29600),
            .I(N__29597));
    LocalMux I__5055 (
            .O(N__29597),
            .I(N__29594));
    Span4Mux_h I__5054 (
            .O(N__29594),
            .I(N__29589));
    InMux I__5053 (
            .O(N__29593),
            .I(N__29584));
    InMux I__5052 (
            .O(N__29592),
            .I(N__29584));
    Span4Mux_v I__5051 (
            .O(N__29589),
            .I(N__29579));
    LocalMux I__5050 (
            .O(N__29584),
            .I(N__29579));
    Span4Mux_h I__5049 (
            .O(N__29579),
            .I(N__29575));
    InMux I__5048 (
            .O(N__29578),
            .I(N__29572));
    Odrv4 I__5047 (
            .O(N__29575),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    LocalMux I__5046 (
            .O(N__29572),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    InMux I__5045 (
            .O(N__29567),
            .I(N__29564));
    LocalMux I__5044 (
            .O(N__29564),
            .I(N__29560));
    InMux I__5043 (
            .O(N__29563),
            .I(N__29557));
    Odrv12 I__5042 (
            .O(N__29560),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    LocalMux I__5041 (
            .O(N__29557),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    CascadeMux I__5040 (
            .O(N__29552),
            .I(N__29549));
    InMux I__5039 (
            .O(N__29549),
            .I(N__29546));
    LocalMux I__5038 (
            .O(N__29546),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    InMux I__5037 (
            .O(N__29543),
            .I(N__29540));
    LocalMux I__5036 (
            .O(N__29540),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__5035 (
            .O(N__29537),
            .I(N__29534));
    InMux I__5034 (
            .O(N__29534),
            .I(N__29531));
    LocalMux I__5033 (
            .O(N__29531),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt20 ));
    InMux I__5032 (
            .O(N__29528),
            .I(N__29522));
    InMux I__5031 (
            .O(N__29527),
            .I(N__29522));
    LocalMux I__5030 (
            .O(N__29522),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ));
    InMux I__5029 (
            .O(N__29519),
            .I(N__29512));
    InMux I__5028 (
            .O(N__29518),
            .I(N__29512));
    InMux I__5027 (
            .O(N__29517),
            .I(N__29509));
    LocalMux I__5026 (
            .O(N__29512),
            .I(N__29506));
    LocalMux I__5025 (
            .O(N__29509),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__5024 (
            .O(N__29506),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    CascadeMux I__5023 (
            .O(N__29501),
            .I(N__29497));
    InMux I__5022 (
            .O(N__29500),
            .I(N__29491));
    InMux I__5021 (
            .O(N__29497),
            .I(N__29491));
    InMux I__5020 (
            .O(N__29496),
            .I(N__29488));
    LocalMux I__5019 (
            .O(N__29491),
            .I(N__29485));
    LocalMux I__5018 (
            .O(N__29488),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__5017 (
            .O(N__29485),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    CascadeMux I__5016 (
            .O(N__29480),
            .I(N__29476));
    InMux I__5015 (
            .O(N__29479),
            .I(N__29471));
    InMux I__5014 (
            .O(N__29476),
            .I(N__29471));
    LocalMux I__5013 (
            .O(N__29471),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    InMux I__5012 (
            .O(N__29468),
            .I(N__29465));
    LocalMux I__5011 (
            .O(N__29465),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ));
    InMux I__5010 (
            .O(N__29462),
            .I(N__29459));
    LocalMux I__5009 (
            .O(N__29459),
            .I(N__29455));
    InMux I__5008 (
            .O(N__29458),
            .I(N__29451));
    Span4Mux_v I__5007 (
            .O(N__29455),
            .I(N__29448));
    InMux I__5006 (
            .O(N__29454),
            .I(N__29445));
    LocalMux I__5005 (
            .O(N__29451),
            .I(N__29442));
    Span4Mux_v I__5004 (
            .O(N__29448),
            .I(N__29436));
    LocalMux I__5003 (
            .O(N__29445),
            .I(N__29436));
    Span4Mux_h I__5002 (
            .O(N__29442),
            .I(N__29433));
    InMux I__5001 (
            .O(N__29441),
            .I(N__29430));
    Odrv4 I__5000 (
            .O(N__29436),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__4999 (
            .O(N__29433),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    LocalMux I__4998 (
            .O(N__29430),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__4997 (
            .O(N__29423),
            .I(N__29420));
    LocalMux I__4996 (
            .O(N__29420),
            .I(N__29416));
    InMux I__4995 (
            .O(N__29419),
            .I(N__29412));
    Span4Mux_v I__4994 (
            .O(N__29416),
            .I(N__29409));
    InMux I__4993 (
            .O(N__29415),
            .I(N__29406));
    LocalMux I__4992 (
            .O(N__29412),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    Odrv4 I__4991 (
            .O(N__29409),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    LocalMux I__4990 (
            .O(N__29406),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    InMux I__4989 (
            .O(N__29399),
            .I(N__29396));
    LocalMux I__4988 (
            .O(N__29396),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__4987 (
            .O(N__29393),
            .I(N__29390));
    InMux I__4986 (
            .O(N__29390),
            .I(N__29387));
    LocalMux I__4985 (
            .O(N__29387),
            .I(N__29384));
    Span4Mux_v I__4984 (
            .O(N__29384),
            .I(N__29381));
    Odrv4 I__4983 (
            .O(N__29381),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    InMux I__4982 (
            .O(N__29378),
            .I(N__29372));
    InMux I__4981 (
            .O(N__29377),
            .I(N__29372));
    LocalMux I__4980 (
            .O(N__29372),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    InMux I__4979 (
            .O(N__29369),
            .I(N__29363));
    InMux I__4978 (
            .O(N__29368),
            .I(N__29363));
    LocalMux I__4977 (
            .O(N__29363),
            .I(N__29359));
    InMux I__4976 (
            .O(N__29362),
            .I(N__29356));
    Span4Mux_h I__4975 (
            .O(N__29359),
            .I(N__29353));
    LocalMux I__4974 (
            .O(N__29356),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__4973 (
            .O(N__29353),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    CascadeMux I__4972 (
            .O(N__29348),
            .I(N__29344));
    InMux I__4971 (
            .O(N__29347),
            .I(N__29339));
    InMux I__4970 (
            .O(N__29344),
            .I(N__29339));
    LocalMux I__4969 (
            .O(N__29339),
            .I(N__29335));
    InMux I__4968 (
            .O(N__29338),
            .I(N__29332));
    Span12Mux_h I__4967 (
            .O(N__29335),
            .I(N__29329));
    LocalMux I__4966 (
            .O(N__29332),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv12 I__4965 (
            .O(N__29329),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__4964 (
            .O(N__29324),
            .I(N__29321));
    LocalMux I__4963 (
            .O(N__29321),
            .I(N__29318));
    Span4Mux_v I__4962 (
            .O(N__29318),
            .I(N__29315));
    Odrv4 I__4961 (
            .O(N__29315),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    InMux I__4960 (
            .O(N__29312),
            .I(N__29309));
    LocalMux I__4959 (
            .O(N__29309),
            .I(N__29304));
    InMux I__4958 (
            .O(N__29308),
            .I(N__29301));
    InMux I__4957 (
            .O(N__29307),
            .I(N__29298));
    Span4Mux_v I__4956 (
            .O(N__29304),
            .I(N__29293));
    LocalMux I__4955 (
            .O(N__29301),
            .I(N__29293));
    LocalMux I__4954 (
            .O(N__29298),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    Odrv4 I__4953 (
            .O(N__29293),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    InMux I__4952 (
            .O(N__29288),
            .I(N__29283));
    InMux I__4951 (
            .O(N__29287),
            .I(N__29280));
    CascadeMux I__4950 (
            .O(N__29286),
            .I(N__29277));
    LocalMux I__4949 (
            .O(N__29283),
            .I(N__29274));
    LocalMux I__4948 (
            .O(N__29280),
            .I(N__29271));
    InMux I__4947 (
            .O(N__29277),
            .I(N__29267));
    Span4Mux_h I__4946 (
            .O(N__29274),
            .I(N__29264));
    Span4Mux_h I__4945 (
            .O(N__29271),
            .I(N__29261));
    InMux I__4944 (
            .O(N__29270),
            .I(N__29258));
    LocalMux I__4943 (
            .O(N__29267),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__4942 (
            .O(N__29264),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__4941 (
            .O(N__29261),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    LocalMux I__4940 (
            .O(N__29258),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    CascadeMux I__4939 (
            .O(N__29249),
            .I(N__29246));
    InMux I__4938 (
            .O(N__29246),
            .I(N__29240));
    InMux I__4937 (
            .O(N__29245),
            .I(N__29240));
    LocalMux I__4936 (
            .O(N__29240),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__4935 (
            .O(N__29237),
            .I(N__29234));
    LocalMux I__4934 (
            .O(N__29234),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    InMux I__4933 (
            .O(N__29231),
            .I(N__29228));
    LocalMux I__4932 (
            .O(N__29228),
            .I(N__29225));
    Span4Mux_h I__4931 (
            .O(N__29225),
            .I(N__29221));
    InMux I__4930 (
            .O(N__29224),
            .I(N__29218));
    Span4Mux_v I__4929 (
            .O(N__29221),
            .I(N__29212));
    LocalMux I__4928 (
            .O(N__29218),
            .I(N__29212));
    InMux I__4927 (
            .O(N__29217),
            .I(N__29209));
    Span4Mux_h I__4926 (
            .O(N__29212),
            .I(N__29206));
    LocalMux I__4925 (
            .O(N__29209),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    Odrv4 I__4924 (
            .O(N__29206),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    InMux I__4923 (
            .O(N__29201),
            .I(N__29198));
    LocalMux I__4922 (
            .O(N__29198),
            .I(N__29194));
    InMux I__4921 (
            .O(N__29197),
            .I(N__29191));
    Span4Mux_v I__4920 (
            .O(N__29194),
            .I(N__29184));
    LocalMux I__4919 (
            .O(N__29191),
            .I(N__29184));
    InMux I__4918 (
            .O(N__29190),
            .I(N__29179));
    InMux I__4917 (
            .O(N__29189),
            .I(N__29179));
    Odrv4 I__4916 (
            .O(N__29184),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__4915 (
            .O(N__29179),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__4914 (
            .O(N__29174),
            .I(N__29171));
    LocalMux I__4913 (
            .O(N__29171),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    InMux I__4912 (
            .O(N__29168),
            .I(N__29165));
    LocalMux I__4911 (
            .O(N__29165),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    InMux I__4910 (
            .O(N__29162),
            .I(N__29156));
    InMux I__4909 (
            .O(N__29161),
            .I(N__29156));
    LocalMux I__4908 (
            .O(N__29156),
            .I(N__29153));
    Span4Mux_h I__4907 (
            .O(N__29153),
            .I(N__29150));
    Odrv4 I__4906 (
            .O(N__29150),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ));
    CascadeMux I__4905 (
            .O(N__29147),
            .I(N__29144));
    InMux I__4904 (
            .O(N__29144),
            .I(N__29141));
    LocalMux I__4903 (
            .O(N__29141),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__4902 (
            .O(N__29138),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_));
    CascadeMux I__4901 (
            .O(N__29135),
            .I(elapsed_time_ns_1_RNI2COBB_0_15_cascade_));
    InMux I__4900 (
            .O(N__29132),
            .I(N__29126));
    InMux I__4899 (
            .O(N__29131),
            .I(N__29126));
    LocalMux I__4898 (
            .O(N__29126),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ));
    CascadeMux I__4897 (
            .O(N__29123),
            .I(N__29119));
    InMux I__4896 (
            .O(N__29122),
            .I(N__29114));
    InMux I__4895 (
            .O(N__29119),
            .I(N__29114));
    LocalMux I__4894 (
            .O(N__29114),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    InMux I__4893 (
            .O(N__29111),
            .I(N__29108));
    LocalMux I__4892 (
            .O(N__29108),
            .I(N__29102));
    InMux I__4891 (
            .O(N__29107),
            .I(N__29099));
    InMux I__4890 (
            .O(N__29106),
            .I(N__29096));
    InMux I__4889 (
            .O(N__29105),
            .I(N__29093));
    Span4Mux_v I__4888 (
            .O(N__29102),
            .I(N__29090));
    LocalMux I__4887 (
            .O(N__29099),
            .I(N__29085));
    LocalMux I__4886 (
            .O(N__29096),
            .I(N__29085));
    LocalMux I__4885 (
            .O(N__29093),
            .I(N__29082));
    Odrv4 I__4884 (
            .O(N__29090),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv12 I__4883 (
            .O(N__29085),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv4 I__4882 (
            .O(N__29082),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__4881 (
            .O(N__29075),
            .I(N__29071));
    InMux I__4880 (
            .O(N__29074),
            .I(N__29067));
    LocalMux I__4879 (
            .O(N__29071),
            .I(N__29064));
    InMux I__4878 (
            .O(N__29070),
            .I(N__29061));
    LocalMux I__4877 (
            .O(N__29067),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    Odrv12 I__4876 (
            .O(N__29064),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    LocalMux I__4875 (
            .O(N__29061),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    InMux I__4874 (
            .O(N__29054),
            .I(N__29048));
    InMux I__4873 (
            .O(N__29053),
            .I(N__29048));
    LocalMux I__4872 (
            .O(N__29048),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ));
    CascadeMux I__4871 (
            .O(N__29045),
            .I(N__29041));
    CascadeMux I__4870 (
            .O(N__29044),
            .I(N__29038));
    InMux I__4869 (
            .O(N__29041),
            .I(N__29033));
    InMux I__4868 (
            .O(N__29038),
            .I(N__29033));
    LocalMux I__4867 (
            .O(N__29033),
            .I(N__29030));
    Odrv4 I__4866 (
            .O(N__29030),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ));
    InMux I__4865 (
            .O(N__29027),
            .I(N__29022));
    InMux I__4864 (
            .O(N__29026),
            .I(N__29019));
    InMux I__4863 (
            .O(N__29025),
            .I(N__29016));
    LocalMux I__4862 (
            .O(N__29022),
            .I(N__29011));
    LocalMux I__4861 (
            .O(N__29019),
            .I(N__29011));
    LocalMux I__4860 (
            .O(N__29016),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    Odrv4 I__4859 (
            .O(N__29011),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    CascadeMux I__4858 (
            .O(N__29006),
            .I(N__29002));
    InMux I__4857 (
            .O(N__29005),
            .I(N__28998));
    InMux I__4856 (
            .O(N__29002),
            .I(N__28995));
    InMux I__4855 (
            .O(N__29001),
            .I(N__28991));
    LocalMux I__4854 (
            .O(N__28998),
            .I(N__28986));
    LocalMux I__4853 (
            .O(N__28995),
            .I(N__28986));
    InMux I__4852 (
            .O(N__28994),
            .I(N__28983));
    LocalMux I__4851 (
            .O(N__28991),
            .I(N__28980));
    Span4Mux_v I__4850 (
            .O(N__28986),
            .I(N__28977));
    LocalMux I__4849 (
            .O(N__28983),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv12 I__4848 (
            .O(N__28980),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__4847 (
            .O(N__28977),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__4846 (
            .O(N__28970),
            .I(N__28967));
    LocalMux I__4845 (
            .O(N__28967),
            .I(N__28963));
    InMux I__4844 (
            .O(N__28966),
            .I(N__28959));
    Span4Mux_v I__4843 (
            .O(N__28963),
            .I(N__28956));
    InMux I__4842 (
            .O(N__28962),
            .I(N__28953));
    LocalMux I__4841 (
            .O(N__28959),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    Odrv4 I__4840 (
            .O(N__28956),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    LocalMux I__4839 (
            .O(N__28953),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    InMux I__4838 (
            .O(N__28946),
            .I(N__28942));
    InMux I__4837 (
            .O(N__28945),
            .I(N__28939));
    LocalMux I__4836 (
            .O(N__28942),
            .I(N__28935));
    LocalMux I__4835 (
            .O(N__28939),
            .I(N__28932));
    InMux I__4834 (
            .O(N__28938),
            .I(N__28929));
    Span4Mux_h I__4833 (
            .O(N__28935),
            .I(N__28925));
    Span4Mux_h I__4832 (
            .O(N__28932),
            .I(N__28922));
    LocalMux I__4831 (
            .O(N__28929),
            .I(N__28919));
    InMux I__4830 (
            .O(N__28928),
            .I(N__28916));
    Odrv4 I__4829 (
            .O(N__28925),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    Odrv4 I__4828 (
            .O(N__28922),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    Odrv12 I__4827 (
            .O(N__28919),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    LocalMux I__4826 (
            .O(N__28916),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__4825 (
            .O(N__28907),
            .I(N__28903));
    InMux I__4824 (
            .O(N__28906),
            .I(N__28899));
    LocalMux I__4823 (
            .O(N__28903),
            .I(N__28896));
    InMux I__4822 (
            .O(N__28902),
            .I(N__28893));
    LocalMux I__4821 (
            .O(N__28899),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv4 I__4820 (
            .O(N__28896),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    LocalMux I__4819 (
            .O(N__28893),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    InMux I__4818 (
            .O(N__28886),
            .I(N__28881));
    InMux I__4817 (
            .O(N__28885),
            .I(N__28878));
    InMux I__4816 (
            .O(N__28884),
            .I(N__28874));
    LocalMux I__4815 (
            .O(N__28881),
            .I(N__28871));
    LocalMux I__4814 (
            .O(N__28878),
            .I(N__28868));
    InMux I__4813 (
            .O(N__28877),
            .I(N__28865));
    LocalMux I__4812 (
            .O(N__28874),
            .I(N__28862));
    Span4Mux_h I__4811 (
            .O(N__28871),
            .I(N__28855));
    Span4Mux_h I__4810 (
            .O(N__28868),
            .I(N__28855));
    LocalMux I__4809 (
            .O(N__28865),
            .I(N__28855));
    Span4Mux_h I__4808 (
            .O(N__28862),
            .I(N__28852));
    Span4Mux_v I__4807 (
            .O(N__28855),
            .I(N__28849));
    Odrv4 I__4806 (
            .O(N__28852),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__4805 (
            .O(N__28849),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__4804 (
            .O(N__28844),
            .I(N__28841));
    LocalMux I__4803 (
            .O(N__28841),
            .I(N__28837));
    InMux I__4802 (
            .O(N__28840),
            .I(N__28834));
    Odrv4 I__4801 (
            .O(N__28837),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    LocalMux I__4800 (
            .O(N__28834),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    InMux I__4799 (
            .O(N__28829),
            .I(N__28824));
    InMux I__4798 (
            .O(N__28828),
            .I(N__28819));
    InMux I__4797 (
            .O(N__28827),
            .I(N__28819));
    LocalMux I__4796 (
            .O(N__28824),
            .I(N__28815));
    LocalMux I__4795 (
            .O(N__28819),
            .I(N__28812));
    InMux I__4794 (
            .O(N__28818),
            .I(N__28809));
    Odrv4 I__4793 (
            .O(N__28815),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    Odrv4 I__4792 (
            .O(N__28812),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    LocalMux I__4791 (
            .O(N__28809),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    CascadeMux I__4790 (
            .O(N__28802),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11_cascade_));
    InMux I__4789 (
            .O(N__28799),
            .I(N__28796));
    LocalMux I__4788 (
            .O(N__28796),
            .I(N__28792));
    InMux I__4787 (
            .O(N__28795),
            .I(N__28789));
    Odrv4 I__4786 (
            .O(N__28792),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    LocalMux I__4785 (
            .O(N__28789),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    InMux I__4784 (
            .O(N__28784),
            .I(N__28777));
    InMux I__4783 (
            .O(N__28783),
            .I(N__28777));
    InMux I__4782 (
            .O(N__28782),
            .I(N__28774));
    LocalMux I__4781 (
            .O(N__28777),
            .I(N__28771));
    LocalMux I__4780 (
            .O(N__28774),
            .I(N__28767));
    Span4Mux_h I__4779 (
            .O(N__28771),
            .I(N__28764));
    InMux I__4778 (
            .O(N__28770),
            .I(N__28761));
    Odrv4 I__4777 (
            .O(N__28767),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    Odrv4 I__4776 (
            .O(N__28764),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__4775 (
            .O(N__28761),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    CascadeMux I__4774 (
            .O(N__28754),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_));
    CascadeMux I__4773 (
            .O(N__28751),
            .I(elapsed_time_ns_1_RNILK91B_0_9_cascade_));
    InMux I__4772 (
            .O(N__28748),
            .I(N__28744));
    InMux I__4771 (
            .O(N__28747),
            .I(N__28741));
    LocalMux I__4770 (
            .O(N__28744),
            .I(N__28736));
    LocalMux I__4769 (
            .O(N__28741),
            .I(N__28733));
    InMux I__4768 (
            .O(N__28740),
            .I(N__28728));
    InMux I__4767 (
            .O(N__28739),
            .I(N__28728));
    Odrv4 I__4766 (
            .O(N__28736),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    Odrv4 I__4765 (
            .O(N__28733),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    LocalMux I__4764 (
            .O(N__28728),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__4763 (
            .O(N__28721),
            .I(N__28716));
    InMux I__4762 (
            .O(N__28720),
            .I(N__28713));
    InMux I__4761 (
            .O(N__28719),
            .I(N__28710));
    LocalMux I__4760 (
            .O(N__28716),
            .I(N__28705));
    LocalMux I__4759 (
            .O(N__28713),
            .I(N__28705));
    LocalMux I__4758 (
            .O(N__28710),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    Odrv12 I__4757 (
            .O(N__28705),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    InMux I__4756 (
            .O(N__28700),
            .I(N__28695));
    InMux I__4755 (
            .O(N__28699),
            .I(N__28692));
    InMux I__4754 (
            .O(N__28698),
            .I(N__28689));
    LocalMux I__4753 (
            .O(N__28695),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__4752 (
            .O(N__28692),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__4751 (
            .O(N__28689),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    InMux I__4750 (
            .O(N__28682),
            .I(N__28676));
    InMux I__4749 (
            .O(N__28681),
            .I(N__28673));
    InMux I__4748 (
            .O(N__28680),
            .I(N__28670));
    CascadeMux I__4747 (
            .O(N__28679),
            .I(N__28667));
    LocalMux I__4746 (
            .O(N__28676),
            .I(N__28664));
    LocalMux I__4745 (
            .O(N__28673),
            .I(N__28659));
    LocalMux I__4744 (
            .O(N__28670),
            .I(N__28659));
    InMux I__4743 (
            .O(N__28667),
            .I(N__28656));
    Span4Mux_v I__4742 (
            .O(N__28664),
            .I(N__28653));
    Span4Mux_h I__4741 (
            .O(N__28659),
            .I(N__28650));
    LocalMux I__4740 (
            .O(N__28656),
            .I(N__28647));
    Odrv4 I__4739 (
            .O(N__28653),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__4738 (
            .O(N__28650),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__4737 (
            .O(N__28647),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__4736 (
            .O(N__28640),
            .I(N__28635));
    InMux I__4735 (
            .O(N__28639),
            .I(N__28632));
    InMux I__4734 (
            .O(N__28638),
            .I(N__28629));
    LocalMux I__4733 (
            .O(N__28635),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    LocalMux I__4732 (
            .O(N__28632),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    LocalMux I__4731 (
            .O(N__28629),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    CascadeMux I__4730 (
            .O(N__28622),
            .I(N__28619));
    InMux I__4729 (
            .O(N__28619),
            .I(N__28614));
    InMux I__4728 (
            .O(N__28618),
            .I(N__28611));
    InMux I__4727 (
            .O(N__28617),
            .I(N__28608));
    LocalMux I__4726 (
            .O(N__28614),
            .I(N__28604));
    LocalMux I__4725 (
            .O(N__28611),
            .I(N__28599));
    LocalMux I__4724 (
            .O(N__28608),
            .I(N__28599));
    CascadeMux I__4723 (
            .O(N__28607),
            .I(N__28596));
    Span4Mux_v I__4722 (
            .O(N__28604),
            .I(N__28593));
    Span4Mux_h I__4721 (
            .O(N__28599),
            .I(N__28590));
    InMux I__4720 (
            .O(N__28596),
            .I(N__28587));
    Odrv4 I__4719 (
            .O(N__28593),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    Odrv4 I__4718 (
            .O(N__28590),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    LocalMux I__4717 (
            .O(N__28587),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__4716 (
            .O(N__28580),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__4715 (
            .O(N__28577),
            .I(N__28574));
    LocalMux I__4714 (
            .O(N__28574),
            .I(N__28571));
    Span4Mux_h I__4713 (
            .O(N__28571),
            .I(N__28568));
    Odrv4 I__4712 (
            .O(N__28568),
            .I(il_min_comp1_c));
    InMux I__4711 (
            .O(N__28565),
            .I(N__28562));
    LocalMux I__4710 (
            .O(N__28562),
            .I(il_min_comp1_D1));
    InMux I__4709 (
            .O(N__28559),
            .I(N__28556));
    LocalMux I__4708 (
            .O(N__28556),
            .I(N__28553));
    Span4Mux_v I__4707 (
            .O(N__28553),
            .I(N__28549));
    InMux I__4706 (
            .O(N__28552),
            .I(N__28546));
    Sp12to4 I__4705 (
            .O(N__28549),
            .I(N__28541));
    LocalMux I__4704 (
            .O(N__28546),
            .I(N__28541));
    Odrv12 I__4703 (
            .O(N__28541),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    InMux I__4702 (
            .O(N__28538),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    CascadeMux I__4701 (
            .O(N__28535),
            .I(N__28532));
    InMux I__4700 (
            .O(N__28532),
            .I(N__28529));
    LocalMux I__4699 (
            .O(N__28529),
            .I(N__28526));
    Span4Mux_v I__4698 (
            .O(N__28526),
            .I(N__28522));
    InMux I__4697 (
            .O(N__28525),
            .I(N__28519));
    Sp12to4 I__4696 (
            .O(N__28522),
            .I(N__28514));
    LocalMux I__4695 (
            .O(N__28519),
            .I(N__28514));
    Odrv12 I__4694 (
            .O(N__28514),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    InMux I__4693 (
            .O(N__28511),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__4692 (
            .O(N__28508),
            .I(N__28505));
    LocalMux I__4691 (
            .O(N__28505),
            .I(N__28502));
    Span4Mux_h I__4690 (
            .O(N__28502),
            .I(N__28499));
    Span4Mux_h I__4689 (
            .O(N__28499),
            .I(N__28496));
    Odrv4 I__4688 (
            .O(N__28496),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ));
    InMux I__4687 (
            .O(N__28493),
            .I(bfn_9_27_0_));
    InMux I__4686 (
            .O(N__28490),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ));
    InMux I__4685 (
            .O(N__28487),
            .I(N__28484));
    LocalMux I__4684 (
            .O(N__28484),
            .I(N__28481));
    Odrv4 I__4683 (
            .O(N__28481),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_31 ));
    InMux I__4682 (
            .O(N__28478),
            .I(N__28475));
    LocalMux I__4681 (
            .O(N__28475),
            .I(N__28472));
    Odrv12 I__4680 (
            .O(N__28472),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ));
    InMux I__4679 (
            .O(N__28469),
            .I(N__28457));
    InMux I__4678 (
            .O(N__28468),
            .I(N__28457));
    InMux I__4677 (
            .O(N__28467),
            .I(N__28457));
    InMux I__4676 (
            .O(N__28466),
            .I(N__28454));
    InMux I__4675 (
            .O(N__28465),
            .I(N__28445));
    InMux I__4674 (
            .O(N__28464),
            .I(N__28445));
    LocalMux I__4673 (
            .O(N__28457),
            .I(N__28442));
    LocalMux I__4672 (
            .O(N__28454),
            .I(N__28439));
    InMux I__4671 (
            .O(N__28453),
            .I(N__28430));
    InMux I__4670 (
            .O(N__28452),
            .I(N__28430));
    InMux I__4669 (
            .O(N__28451),
            .I(N__28430));
    InMux I__4668 (
            .O(N__28450),
            .I(N__28430));
    LocalMux I__4667 (
            .O(N__28445),
            .I(N__28427));
    Span4Mux_h I__4666 (
            .O(N__28442),
            .I(N__28422));
    Span4Mux_h I__4665 (
            .O(N__28439),
            .I(N__28422));
    LocalMux I__4664 (
            .O(N__28430),
            .I(N__28419));
    Span4Mux_h I__4663 (
            .O(N__28427),
            .I(N__28416));
    Span4Mux_h I__4662 (
            .O(N__28422),
            .I(N__28413));
    Span4Mux_h I__4661 (
            .O(N__28419),
            .I(N__28410));
    Odrv4 I__4660 (
            .O(N__28416),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__4659 (
            .O(N__28413),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__4658 (
            .O(N__28410),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__4657 (
            .O(N__28403),
            .I(N__28400));
    LocalMux I__4656 (
            .O(N__28400),
            .I(N__28397));
    Span4Mux_v I__4655 (
            .O(N__28397),
            .I(N__28394));
    Span4Mux_h I__4654 (
            .O(N__28394),
            .I(N__28390));
    InMux I__4653 (
            .O(N__28393),
            .I(N__28387));
    Span4Mux_h I__4652 (
            .O(N__28390),
            .I(N__28384));
    LocalMux I__4651 (
            .O(N__28387),
            .I(\pwm_generator_inst.un3_threshold ));
    Odrv4 I__4650 (
            .O(N__28384),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__4649 (
            .O(N__28379),
            .I(N__28376));
    LocalMux I__4648 (
            .O(N__28376),
            .I(N__28373));
    Span4Mux_v I__4647 (
            .O(N__28373),
            .I(N__28370));
    Sp12to4 I__4646 (
            .O(N__28370),
            .I(N__28367));
    Odrv12 I__4645 (
            .O(N__28367),
            .I(\pwm_generator_inst.O_12 ));
    CascadeMux I__4644 (
            .O(N__28364),
            .I(N__28361));
    InMux I__4643 (
            .O(N__28361),
            .I(N__28358));
    LocalMux I__4642 (
            .O(N__28358),
            .I(N__28354));
    InMux I__4641 (
            .O(N__28357),
            .I(N__28351));
    Sp12to4 I__4640 (
            .O(N__28354),
            .I(N__28348));
    LocalMux I__4639 (
            .O(N__28351),
            .I(N__28345));
    Span12Mux_v I__4638 (
            .O(N__28348),
            .I(N__28340));
    Span12Mux_s4_h I__4637 (
            .O(N__28345),
            .I(N__28340));
    Odrv12 I__4636 (
            .O(N__28340),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    InMux I__4635 (
            .O(N__28337),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__4634 (
            .O(N__28334),
            .I(N__28331));
    LocalMux I__4633 (
            .O(N__28331),
            .I(N__28328));
    Span4Mux_v I__4632 (
            .O(N__28328),
            .I(N__28325));
    Sp12to4 I__4631 (
            .O(N__28325),
            .I(N__28322));
    Odrv12 I__4630 (
            .O(N__28322),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__4629 (
            .O(N__28319),
            .I(N__28315));
    InMux I__4628 (
            .O(N__28318),
            .I(N__28312));
    LocalMux I__4627 (
            .O(N__28315),
            .I(N__28309));
    LocalMux I__4626 (
            .O(N__28312),
            .I(N__28306));
    Span12Mux_v I__4625 (
            .O(N__28309),
            .I(N__28301));
    Span12Mux_s3_h I__4624 (
            .O(N__28306),
            .I(N__28301));
    Odrv12 I__4623 (
            .O(N__28301),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    InMux I__4622 (
            .O(N__28298),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__4621 (
            .O(N__28295),
            .I(N__28292));
    LocalMux I__4620 (
            .O(N__28292),
            .I(N__28289));
    Span4Mux_v I__4619 (
            .O(N__28289),
            .I(N__28286));
    Sp12to4 I__4618 (
            .O(N__28286),
            .I(N__28283));
    Odrv12 I__4617 (
            .O(N__28283),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__4616 (
            .O(N__28280),
            .I(N__28277));
    LocalMux I__4615 (
            .O(N__28277),
            .I(N__28274));
    Span4Mux_v I__4614 (
            .O(N__28274),
            .I(N__28270));
    InMux I__4613 (
            .O(N__28273),
            .I(N__28267));
    Sp12to4 I__4612 (
            .O(N__28270),
            .I(N__28262));
    LocalMux I__4611 (
            .O(N__28267),
            .I(N__28262));
    Odrv12 I__4610 (
            .O(N__28262),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    InMux I__4609 (
            .O(N__28259),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__4608 (
            .O(N__28256),
            .I(N__28252));
    InMux I__4607 (
            .O(N__28255),
            .I(N__28249));
    LocalMux I__4606 (
            .O(N__28252),
            .I(N__28244));
    LocalMux I__4605 (
            .O(N__28249),
            .I(N__28244));
    Span4Mux_h I__4604 (
            .O(N__28244),
            .I(N__28241));
    Span4Mux_h I__4603 (
            .O(N__28241),
            .I(N__28238));
    Odrv4 I__4602 (
            .O(N__28238),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    InMux I__4601 (
            .O(N__28235),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    InMux I__4600 (
            .O(N__28232),
            .I(N__28229));
    LocalMux I__4599 (
            .O(N__28229),
            .I(N__28226));
    Span4Mux_v I__4598 (
            .O(N__28226),
            .I(N__28222));
    InMux I__4597 (
            .O(N__28225),
            .I(N__28219));
    Sp12to4 I__4596 (
            .O(N__28222),
            .I(N__28214));
    LocalMux I__4595 (
            .O(N__28219),
            .I(N__28214));
    Odrv12 I__4594 (
            .O(N__28214),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    InMux I__4593 (
            .O(N__28211),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__4592 (
            .O(N__28208),
            .I(N__28205));
    LocalMux I__4591 (
            .O(N__28205),
            .I(N__28202));
    Span4Mux_v I__4590 (
            .O(N__28202),
            .I(N__28198));
    InMux I__4589 (
            .O(N__28201),
            .I(N__28195));
    Span4Mux_h I__4588 (
            .O(N__28198),
            .I(N__28192));
    LocalMux I__4587 (
            .O(N__28195),
            .I(N__28189));
    Span4Mux_v I__4586 (
            .O(N__28192),
            .I(N__28186));
    Span4Mux_h I__4585 (
            .O(N__28189),
            .I(N__28181));
    Span4Mux_h I__4584 (
            .O(N__28186),
            .I(N__28181));
    Odrv4 I__4583 (
            .O(N__28181),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    InMux I__4582 (
            .O(N__28178),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ));
    InMux I__4581 (
            .O(N__28175),
            .I(N__28172));
    LocalMux I__4580 (
            .O(N__28172),
            .I(N__28168));
    InMux I__4579 (
            .O(N__28171),
            .I(N__28165));
    Span4Mux_v I__4578 (
            .O(N__28168),
            .I(N__28162));
    LocalMux I__4577 (
            .O(N__28165),
            .I(N__28159));
    Sp12to4 I__4576 (
            .O(N__28162),
            .I(N__28156));
    Span4Mux_h I__4575 (
            .O(N__28159),
            .I(N__28153));
    Span12Mux_s9_h I__4574 (
            .O(N__28156),
            .I(N__28150));
    Odrv4 I__4573 (
            .O(N__28153),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    Odrv12 I__4572 (
            .O(N__28150),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    InMux I__4571 (
            .O(N__28145),
            .I(bfn_9_18_0_));
    InMux I__4570 (
            .O(N__28142),
            .I(N__28138));
    InMux I__4569 (
            .O(N__28141),
            .I(N__28135));
    LocalMux I__4568 (
            .O(N__28138),
            .I(N__28132));
    LocalMux I__4567 (
            .O(N__28135),
            .I(N__28129));
    Span4Mux_h I__4566 (
            .O(N__28132),
            .I(N__28126));
    Span12Mux_s9_h I__4565 (
            .O(N__28129),
            .I(N__28123));
    Odrv4 I__4564 (
            .O(N__28126),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    Odrv12 I__4563 (
            .O(N__28123),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    InMux I__4562 (
            .O(N__28118),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ));
    InMux I__4561 (
            .O(N__28115),
            .I(N__28112));
    LocalMux I__4560 (
            .O(N__28112),
            .I(N__28108));
    InMux I__4559 (
            .O(N__28111),
            .I(N__28105));
    Span4Mux_v I__4558 (
            .O(N__28108),
            .I(N__28102));
    LocalMux I__4557 (
            .O(N__28105),
            .I(N__28099));
    Sp12to4 I__4556 (
            .O(N__28102),
            .I(N__28096));
    Span4Mux_v I__4555 (
            .O(N__28099),
            .I(N__28093));
    Span12Mux_s9_h I__4554 (
            .O(N__28096),
            .I(N__28090));
    Odrv4 I__4553 (
            .O(N__28093),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    Odrv12 I__4552 (
            .O(N__28090),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    InMux I__4551 (
            .O(N__28085),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ));
    InMux I__4550 (
            .O(N__28082),
            .I(N__28079));
    LocalMux I__4549 (
            .O(N__28079),
            .I(N__28076));
    Span4Mux_s2_h I__4548 (
            .O(N__28076),
            .I(N__28072));
    InMux I__4547 (
            .O(N__28075),
            .I(N__28069));
    Sp12to4 I__4546 (
            .O(N__28072),
            .I(N__28066));
    LocalMux I__4545 (
            .O(N__28069),
            .I(N__28061));
    Span12Mux_v I__4544 (
            .O(N__28066),
            .I(N__28061));
    Odrv12 I__4543 (
            .O(N__28061),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    InMux I__4542 (
            .O(N__28058),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ));
    InMux I__4541 (
            .O(N__28055),
            .I(N__28052));
    LocalMux I__4540 (
            .O(N__28052),
            .I(N__28049));
    Span4Mux_v I__4539 (
            .O(N__28049),
            .I(N__28045));
    InMux I__4538 (
            .O(N__28048),
            .I(N__28042));
    Sp12to4 I__4537 (
            .O(N__28045),
            .I(N__28039));
    LocalMux I__4536 (
            .O(N__28042),
            .I(N__28036));
    Span12Mux_s9_h I__4535 (
            .O(N__28039),
            .I(N__28033));
    Odrv12 I__4534 (
            .O(N__28036),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    Odrv12 I__4533 (
            .O(N__28033),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    InMux I__4532 (
            .O(N__28028),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ));
    InMux I__4531 (
            .O(N__28025),
            .I(N__28021));
    InMux I__4530 (
            .O(N__28024),
            .I(N__28018));
    LocalMux I__4529 (
            .O(N__28021),
            .I(N__28015));
    LocalMux I__4528 (
            .O(N__28018),
            .I(N__28012));
    Span4Mux_v I__4527 (
            .O(N__28015),
            .I(N__28009));
    Span12Mux_v I__4526 (
            .O(N__28012),
            .I(N__28006));
    Odrv4 I__4525 (
            .O(N__28009),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    Odrv12 I__4524 (
            .O(N__28006),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    InMux I__4523 (
            .O(N__28001),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ));
    InMux I__4522 (
            .O(N__27998),
            .I(N__27995));
    LocalMux I__4521 (
            .O(N__27995),
            .I(N__27992));
    Span4Mux_v I__4520 (
            .O(N__27992),
            .I(N__27988));
    InMux I__4519 (
            .O(N__27991),
            .I(N__27985));
    Span4Mux_v I__4518 (
            .O(N__27988),
            .I(N__27982));
    LocalMux I__4517 (
            .O(N__27985),
            .I(N__27979));
    Span4Mux_v I__4516 (
            .O(N__27982),
            .I(N__27976));
    Span4Mux_h I__4515 (
            .O(N__27979),
            .I(N__27973));
    Sp12to4 I__4514 (
            .O(N__27976),
            .I(N__27970));
    Odrv4 I__4513 (
            .O(N__27973),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    Odrv12 I__4512 (
            .O(N__27970),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    InMux I__4511 (
            .O(N__27965),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ));
    InMux I__4510 (
            .O(N__27962),
            .I(N__27959));
    LocalMux I__4509 (
            .O(N__27959),
            .I(N__27956));
    Span4Mux_v I__4508 (
            .O(N__27956),
            .I(N__27952));
    InMux I__4507 (
            .O(N__27955),
            .I(N__27949));
    Span4Mux_v I__4506 (
            .O(N__27952),
            .I(N__27946));
    LocalMux I__4505 (
            .O(N__27949),
            .I(N__27943));
    Span4Mux_h I__4504 (
            .O(N__27946),
            .I(N__27940));
    Span4Mux_h I__4503 (
            .O(N__27943),
            .I(N__27935));
    Span4Mux_h I__4502 (
            .O(N__27940),
            .I(N__27935));
    Odrv4 I__4501 (
            .O(N__27935),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    InMux I__4500 (
            .O(N__27932),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ));
    InMux I__4499 (
            .O(N__27929),
            .I(N__27926));
    LocalMux I__4498 (
            .O(N__27926),
            .I(N__27923));
    Span4Mux_v I__4497 (
            .O(N__27923),
            .I(N__27919));
    InMux I__4496 (
            .O(N__27922),
            .I(N__27916));
    Sp12to4 I__4495 (
            .O(N__27919),
            .I(N__27913));
    LocalMux I__4494 (
            .O(N__27916),
            .I(N__27910));
    Span12Mux_s9_h I__4493 (
            .O(N__27913),
            .I(N__27907));
    Odrv12 I__4492 (
            .O(N__27910),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv12 I__4491 (
            .O(N__27907),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    InMux I__4490 (
            .O(N__27902),
            .I(bfn_9_17_0_));
    InMux I__4489 (
            .O(N__27899),
            .I(N__27896));
    LocalMux I__4488 (
            .O(N__27896),
            .I(N__27893));
    Span4Mux_v I__4487 (
            .O(N__27893),
            .I(N__27889));
    InMux I__4486 (
            .O(N__27892),
            .I(N__27886));
    Span4Mux_v I__4485 (
            .O(N__27889),
            .I(N__27883));
    LocalMux I__4484 (
            .O(N__27886),
            .I(N__27880));
    Span4Mux_h I__4483 (
            .O(N__27883),
            .I(N__27877));
    Span4Mux_h I__4482 (
            .O(N__27880),
            .I(N__27874));
    Span4Mux_h I__4481 (
            .O(N__27877),
            .I(N__27871));
    Odrv4 I__4480 (
            .O(N__27874),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    Odrv4 I__4479 (
            .O(N__27871),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    InMux I__4478 (
            .O(N__27866),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ));
    InMux I__4477 (
            .O(N__27863),
            .I(N__27860));
    LocalMux I__4476 (
            .O(N__27860),
            .I(N__27856));
    InMux I__4475 (
            .O(N__27859),
            .I(N__27853));
    Span4Mux_h I__4474 (
            .O(N__27856),
            .I(N__27850));
    LocalMux I__4473 (
            .O(N__27853),
            .I(N__27847));
    Span4Mux_h I__4472 (
            .O(N__27850),
            .I(N__27844));
    Span12Mux_s9_h I__4471 (
            .O(N__27847),
            .I(N__27841));
    Odrv4 I__4470 (
            .O(N__27844),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    Odrv12 I__4469 (
            .O(N__27841),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    InMux I__4468 (
            .O(N__27836),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ));
    InMux I__4467 (
            .O(N__27833),
            .I(N__27830));
    LocalMux I__4466 (
            .O(N__27830),
            .I(N__27827));
    Span4Mux_v I__4465 (
            .O(N__27827),
            .I(N__27823));
    InMux I__4464 (
            .O(N__27826),
            .I(N__27820));
    Span4Mux_h I__4463 (
            .O(N__27823),
            .I(N__27817));
    LocalMux I__4462 (
            .O(N__27820),
            .I(N__27814));
    Span4Mux_v I__4461 (
            .O(N__27817),
            .I(N__27811));
    Span4Mux_h I__4460 (
            .O(N__27814),
            .I(N__27806));
    Span4Mux_h I__4459 (
            .O(N__27811),
            .I(N__27806));
    Odrv4 I__4458 (
            .O(N__27806),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    InMux I__4457 (
            .O(N__27803),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ));
    InMux I__4456 (
            .O(N__27800),
            .I(N__27796));
    InMux I__4455 (
            .O(N__27799),
            .I(N__27793));
    LocalMux I__4454 (
            .O(N__27796),
            .I(N__27790));
    LocalMux I__4453 (
            .O(N__27793),
            .I(N__27787));
    Span4Mux_v I__4452 (
            .O(N__27790),
            .I(N__27784));
    Span4Mux_h I__4451 (
            .O(N__27787),
            .I(N__27781));
    Sp12to4 I__4450 (
            .O(N__27784),
            .I(N__27778));
    Span4Mux_h I__4449 (
            .O(N__27781),
            .I(N__27775));
    Span12Mux_s9_h I__4448 (
            .O(N__27778),
            .I(N__27772));
    Odrv4 I__4447 (
            .O(N__27775),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    Odrv12 I__4446 (
            .O(N__27772),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    InMux I__4445 (
            .O(N__27767),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ));
    InMux I__4444 (
            .O(N__27764),
            .I(N__27760));
    InMux I__4443 (
            .O(N__27763),
            .I(N__27757));
    LocalMux I__4442 (
            .O(N__27760),
            .I(N__27754));
    LocalMux I__4441 (
            .O(N__27757),
            .I(N__27751));
    Span4Mux_v I__4440 (
            .O(N__27754),
            .I(N__27748));
    Span12Mux_v I__4439 (
            .O(N__27751),
            .I(N__27745));
    Odrv4 I__4438 (
            .O(N__27748),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    Odrv12 I__4437 (
            .O(N__27745),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    InMux I__4436 (
            .O(N__27740),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ));
    InMux I__4435 (
            .O(N__27737),
            .I(N__27734));
    LocalMux I__4434 (
            .O(N__27734),
            .I(N__27730));
    InMux I__4433 (
            .O(N__27733),
            .I(N__27727));
    Span4Mux_v I__4432 (
            .O(N__27730),
            .I(N__27724));
    LocalMux I__4431 (
            .O(N__27727),
            .I(N__27721));
    Span4Mux_v I__4430 (
            .O(N__27724),
            .I(N__27718));
    Span4Mux_v I__4429 (
            .O(N__27721),
            .I(N__27713));
    Span4Mux_h I__4428 (
            .O(N__27718),
            .I(N__27713));
    Span4Mux_h I__4427 (
            .O(N__27713),
            .I(N__27710));
    Odrv4 I__4426 (
            .O(N__27710),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    InMux I__4425 (
            .O(N__27707),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ));
    InMux I__4424 (
            .O(N__27704),
            .I(N__27701));
    LocalMux I__4423 (
            .O(N__27701),
            .I(N__27697));
    InMux I__4422 (
            .O(N__27700),
            .I(N__27694));
    Span4Mux_v I__4421 (
            .O(N__27697),
            .I(N__27691));
    LocalMux I__4420 (
            .O(N__27694),
            .I(N__27686));
    Sp12to4 I__4419 (
            .O(N__27691),
            .I(N__27686));
    Odrv12 I__4418 (
            .O(N__27686),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__4417 (
            .O(N__27683),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__4416 (
            .O(N__27680),
            .I(N__27677));
    LocalMux I__4415 (
            .O(N__27677),
            .I(N__27674));
    Span4Mux_s2_h I__4414 (
            .O(N__27674),
            .I(N__27670));
    InMux I__4413 (
            .O(N__27673),
            .I(N__27667));
    Span4Mux_h I__4412 (
            .O(N__27670),
            .I(N__27664));
    LocalMux I__4411 (
            .O(N__27667),
            .I(N__27661));
    Span4Mux_h I__4410 (
            .O(N__27664),
            .I(N__27658));
    Odrv12 I__4409 (
            .O(N__27661),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__4408 (
            .O(N__27658),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__4407 (
            .O(N__27653),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__4406 (
            .O(N__27650),
            .I(N__27646));
    InMux I__4405 (
            .O(N__27649),
            .I(N__27643));
    LocalMux I__4404 (
            .O(N__27646),
            .I(N__27640));
    LocalMux I__4403 (
            .O(N__27643),
            .I(N__27637));
    Span12Mux_s9_h I__4402 (
            .O(N__27640),
            .I(N__27634));
    Odrv12 I__4401 (
            .O(N__27637),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv12 I__4400 (
            .O(N__27634),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__4399 (
            .O(N__27629),
            .I(bfn_9_16_0_));
    InMux I__4398 (
            .O(N__27626),
            .I(N__27623));
    LocalMux I__4397 (
            .O(N__27623),
            .I(N__27619));
    InMux I__4396 (
            .O(N__27622),
            .I(N__27616));
    Span4Mux_s1_h I__4395 (
            .O(N__27619),
            .I(N__27613));
    LocalMux I__4394 (
            .O(N__27616),
            .I(N__27610));
    Span4Mux_h I__4393 (
            .O(N__27613),
            .I(N__27607));
    Span4Mux_h I__4392 (
            .O(N__27610),
            .I(N__27604));
    Span4Mux_h I__4391 (
            .O(N__27607),
            .I(N__27601));
    Odrv4 I__4390 (
            .O(N__27604),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv4 I__4389 (
            .O(N__27601),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__4388 (
            .O(N__27596),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__4387 (
            .O(N__27593),
            .I(N__27589));
    InMux I__4386 (
            .O(N__27592),
            .I(N__27586));
    LocalMux I__4385 (
            .O(N__27589),
            .I(N__27583));
    LocalMux I__4384 (
            .O(N__27586),
            .I(N__27580));
    Span4Mux_s2_h I__4383 (
            .O(N__27583),
            .I(N__27577));
    Span4Mux_h I__4382 (
            .O(N__27580),
            .I(N__27574));
    Span4Mux_h I__4381 (
            .O(N__27577),
            .I(N__27571));
    Span4Mux_h I__4380 (
            .O(N__27574),
            .I(N__27568));
    Span4Mux_h I__4379 (
            .O(N__27571),
            .I(N__27565));
    Odrv4 I__4378 (
            .O(N__27568),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv4 I__4377 (
            .O(N__27565),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__4376 (
            .O(N__27560),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__4375 (
            .O(N__27557),
            .I(N__27554));
    LocalMux I__4374 (
            .O(N__27554),
            .I(N__27551));
    Span4Mux_s2_h I__4373 (
            .O(N__27551),
            .I(N__27547));
    InMux I__4372 (
            .O(N__27550),
            .I(N__27544));
    Span4Mux_h I__4371 (
            .O(N__27547),
            .I(N__27541));
    LocalMux I__4370 (
            .O(N__27544),
            .I(N__27538));
    Span4Mux_h I__4369 (
            .O(N__27541),
            .I(N__27535));
    Odrv12 I__4368 (
            .O(N__27538),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv4 I__4367 (
            .O(N__27535),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__4366 (
            .O(N__27530),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__4365 (
            .O(N__27527),
            .I(N__27524));
    LocalMux I__4364 (
            .O(N__27524),
            .I(N__27521));
    Span4Mux_s1_h I__4363 (
            .O(N__27521),
            .I(N__27517));
    InMux I__4362 (
            .O(N__27520),
            .I(N__27514));
    Span4Mux_h I__4361 (
            .O(N__27517),
            .I(N__27511));
    LocalMux I__4360 (
            .O(N__27514),
            .I(N__27508));
    Span4Mux_h I__4359 (
            .O(N__27511),
            .I(N__27505));
    Odrv12 I__4358 (
            .O(N__27508),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__4357 (
            .O(N__27505),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__4356 (
            .O(N__27500),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__4355 (
            .O(N__27497),
            .I(N__27494));
    LocalMux I__4354 (
            .O(N__27494),
            .I(N__27490));
    InMux I__4353 (
            .O(N__27493),
            .I(N__27487));
    Span4Mux_v I__4352 (
            .O(N__27490),
            .I(N__27484));
    LocalMux I__4351 (
            .O(N__27487),
            .I(N__27481));
    Sp12to4 I__4350 (
            .O(N__27484),
            .I(N__27476));
    Span12Mux_v I__4349 (
            .O(N__27481),
            .I(N__27476));
    Odrv12 I__4348 (
            .O(N__27476),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__4347 (
            .O(N__27473),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__4346 (
            .O(N__27470),
            .I(N__27467));
    LocalMux I__4345 (
            .O(N__27467),
            .I(N__27463));
    InMux I__4344 (
            .O(N__27466),
            .I(N__27460));
    Span4Mux_s2_h I__4343 (
            .O(N__27463),
            .I(N__27457));
    LocalMux I__4342 (
            .O(N__27460),
            .I(N__27454));
    Span4Mux_v I__4341 (
            .O(N__27457),
            .I(N__27451));
    Span4Mux_v I__4340 (
            .O(N__27454),
            .I(N__27446));
    Span4Mux_h I__4339 (
            .O(N__27451),
            .I(N__27446));
    Odrv4 I__4338 (
            .O(N__27446),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__4337 (
            .O(N__27443),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__4336 (
            .O(N__27440),
            .I(N__27437));
    LocalMux I__4335 (
            .O(N__27437),
            .I(N__27434));
    Odrv4 I__4334 (
            .O(N__27434),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    CascadeMux I__4333 (
            .O(N__27431),
            .I(N__27428));
    InMux I__4332 (
            .O(N__27428),
            .I(N__27425));
    LocalMux I__4331 (
            .O(N__27425),
            .I(N__27422));
    Span4Mux_v I__4330 (
            .O(N__27422),
            .I(N__27419));
    Odrv4 I__4329 (
            .O(N__27419),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    InMux I__4328 (
            .O(N__27416),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ));
    InMux I__4327 (
            .O(N__27413),
            .I(N__27410));
    LocalMux I__4326 (
            .O(N__27410),
            .I(N__27405));
    InMux I__4325 (
            .O(N__27409),
            .I(N__27400));
    InMux I__4324 (
            .O(N__27408),
            .I(N__27400));
    Span4Mux_h I__4323 (
            .O(N__27405),
            .I(N__27397));
    LocalMux I__4322 (
            .O(N__27400),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__4321 (
            .O(N__27397),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__4320 (
            .O(N__27392),
            .I(N__27389));
    LocalMux I__4319 (
            .O(N__27389),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__4318 (
            .O(N__27386),
            .I(N__27382));
    InMux I__4317 (
            .O(N__27385),
            .I(N__27379));
    LocalMux I__4316 (
            .O(N__27382),
            .I(N__27376));
    LocalMux I__4315 (
            .O(N__27379),
            .I(N__27373));
    Span4Mux_h I__4314 (
            .O(N__27376),
            .I(N__27370));
    Span12Mux_s9_h I__4313 (
            .O(N__27373),
            .I(N__27367));
    Odrv4 I__4312 (
            .O(N__27370),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    Odrv12 I__4311 (
            .O(N__27367),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__4310 (
            .O(N__27362),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__4309 (
            .O(N__27359),
            .I(N__27356));
    LocalMux I__4308 (
            .O(N__27356),
            .I(N__27353));
    Span4Mux_s1_h I__4307 (
            .O(N__27353),
            .I(N__27349));
    InMux I__4306 (
            .O(N__27352),
            .I(N__27346));
    Span4Mux_h I__4305 (
            .O(N__27349),
            .I(N__27343));
    LocalMux I__4304 (
            .O(N__27346),
            .I(N__27340));
    Span4Mux_h I__4303 (
            .O(N__27343),
            .I(N__27337));
    Odrv12 I__4302 (
            .O(N__27340),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv4 I__4301 (
            .O(N__27337),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__4300 (
            .O(N__27332),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__4299 (
            .O(N__27329),
            .I(N__27325));
    InMux I__4298 (
            .O(N__27328),
            .I(N__27322));
    LocalMux I__4297 (
            .O(N__27325),
            .I(N__27319));
    LocalMux I__4296 (
            .O(N__27322),
            .I(N__27316));
    Span4Mux_s1_h I__4295 (
            .O(N__27319),
            .I(N__27313));
    Span4Mux_v I__4294 (
            .O(N__27316),
            .I(N__27308));
    Span4Mux_h I__4293 (
            .O(N__27313),
            .I(N__27308));
    Span4Mux_h I__4292 (
            .O(N__27308),
            .I(N__27305));
    Odrv4 I__4291 (
            .O(N__27305),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__4290 (
            .O(N__27302),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__4289 (
            .O(N__27299),
            .I(N__27296));
    LocalMux I__4288 (
            .O(N__27296),
            .I(N__27292));
    InMux I__4287 (
            .O(N__27295),
            .I(N__27289));
    Span4Mux_v I__4286 (
            .O(N__27292),
            .I(N__27286));
    LocalMux I__4285 (
            .O(N__27289),
            .I(N__27281));
    Sp12to4 I__4284 (
            .O(N__27286),
            .I(N__27281));
    Odrv12 I__4283 (
            .O(N__27281),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__4282 (
            .O(N__27278),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__4281 (
            .O(N__27275),
            .I(N__27272));
    LocalMux I__4280 (
            .O(N__27272),
            .I(N__27268));
    InMux I__4279 (
            .O(N__27271),
            .I(N__27265));
    Span4Mux_v I__4278 (
            .O(N__27268),
            .I(N__27262));
    LocalMux I__4277 (
            .O(N__27265),
            .I(N__27259));
    Sp12to4 I__4276 (
            .O(N__27262),
            .I(N__27254));
    Span12Mux_v I__4275 (
            .O(N__27259),
            .I(N__27254));
    Odrv12 I__4274 (
            .O(N__27254),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__4273 (
            .O(N__27251),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__4272 (
            .O(N__27248),
            .I(N__27244));
    InMux I__4271 (
            .O(N__27247),
            .I(N__27241));
    LocalMux I__4270 (
            .O(N__27244),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__4269 (
            .O(N__27241),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__4268 (
            .O(N__27236),
            .I(N__27233));
    LocalMux I__4267 (
            .O(N__27233),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__4266 (
            .O(N__27230),
            .I(N__27227));
    LocalMux I__4265 (
            .O(N__27227),
            .I(N__27224));
    Odrv12 I__4264 (
            .O(N__27224),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ));
    CascadeMux I__4263 (
            .O(N__27221),
            .I(N__27218));
    InMux I__4262 (
            .O(N__27218),
            .I(N__27215));
    LocalMux I__4261 (
            .O(N__27215),
            .I(N__27212));
    Odrv12 I__4260 (
            .O(N__27212),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt22 ));
    InMux I__4259 (
            .O(N__27209),
            .I(N__27206));
    LocalMux I__4258 (
            .O(N__27206),
            .I(N__27203));
    Odrv12 I__4257 (
            .O(N__27203),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ));
    CascadeMux I__4256 (
            .O(N__27200),
            .I(N__27197));
    InMux I__4255 (
            .O(N__27197),
            .I(N__27194));
    LocalMux I__4254 (
            .O(N__27194),
            .I(N__27191));
    Span4Mux_v I__4253 (
            .O(N__27191),
            .I(N__27188));
    Odrv4 I__4252 (
            .O(N__27188),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt24 ));
    InMux I__4251 (
            .O(N__27185),
            .I(N__27182));
    LocalMux I__4250 (
            .O(N__27182),
            .I(N__27179));
    Odrv4 I__4249 (
            .O(N__27179),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt26 ));
    CascadeMux I__4248 (
            .O(N__27176),
            .I(N__27173));
    InMux I__4247 (
            .O(N__27173),
            .I(N__27170));
    LocalMux I__4246 (
            .O(N__27170),
            .I(N__27167));
    Odrv4 I__4245 (
            .O(N__27167),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ));
    InMux I__4244 (
            .O(N__27164),
            .I(N__27161));
    LocalMux I__4243 (
            .O(N__27161),
            .I(N__27158));
    Span4Mux_h I__4242 (
            .O(N__27158),
            .I(N__27155));
    Odrv4 I__4241 (
            .O(N__27155),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt28 ));
    CascadeMux I__4240 (
            .O(N__27152),
            .I(N__27149));
    InMux I__4239 (
            .O(N__27149),
            .I(N__27146));
    LocalMux I__4238 (
            .O(N__27146),
            .I(N__27143));
    Span4Mux_h I__4237 (
            .O(N__27143),
            .I(N__27140));
    Odrv4 I__4236 (
            .O(N__27140),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ));
    InMux I__4235 (
            .O(N__27137),
            .I(N__27134));
    LocalMux I__4234 (
            .O(N__27134),
            .I(N__27131));
    Odrv4 I__4233 (
            .O(N__27131),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    InMux I__4232 (
            .O(N__27128),
            .I(N__27124));
    InMux I__4231 (
            .O(N__27127),
            .I(N__27121));
    LocalMux I__4230 (
            .O(N__27124),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__4229 (
            .O(N__27121),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__4228 (
            .O(N__27116),
            .I(N__27113));
    InMux I__4227 (
            .O(N__27113),
            .I(N__27110));
    LocalMux I__4226 (
            .O(N__27110),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    InMux I__4225 (
            .O(N__27107),
            .I(N__27103));
    InMux I__4224 (
            .O(N__27106),
            .I(N__27100));
    LocalMux I__4223 (
            .O(N__27103),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__4222 (
            .O(N__27100),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__4221 (
            .O(N__27095),
            .I(N__27092));
    LocalMux I__4220 (
            .O(N__27092),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__4219 (
            .O(N__27089),
            .I(N__27085));
    InMux I__4218 (
            .O(N__27088),
            .I(N__27082));
    LocalMux I__4217 (
            .O(N__27085),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__4216 (
            .O(N__27082),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__4215 (
            .O(N__27077),
            .I(N__27074));
    LocalMux I__4214 (
            .O(N__27074),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__4213 (
            .O(N__27071),
            .I(N__27068));
    LocalMux I__4212 (
            .O(N__27068),
            .I(N__27065));
    Odrv4 I__4211 (
            .O(N__27065),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    InMux I__4210 (
            .O(N__27062),
            .I(N__27059));
    LocalMux I__4209 (
            .O(N__27059),
            .I(N__27055));
    InMux I__4208 (
            .O(N__27058),
            .I(N__27052));
    Span4Mux_v I__4207 (
            .O(N__27055),
            .I(N__27049));
    LocalMux I__4206 (
            .O(N__27052),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__4205 (
            .O(N__27049),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    CascadeMux I__4204 (
            .O(N__27044),
            .I(N__27041));
    InMux I__4203 (
            .O(N__27041),
            .I(N__27038));
    LocalMux I__4202 (
            .O(N__27038),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__4201 (
            .O(N__27035),
            .I(N__27032));
    LocalMux I__4200 (
            .O(N__27032),
            .I(N__27029));
    Odrv4 I__4199 (
            .O(N__27029),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    InMux I__4198 (
            .O(N__27026),
            .I(N__27022));
    InMux I__4197 (
            .O(N__27025),
            .I(N__27019));
    LocalMux I__4196 (
            .O(N__27022),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__4195 (
            .O(N__27019),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    CascadeMux I__4194 (
            .O(N__27014),
            .I(N__27011));
    InMux I__4193 (
            .O(N__27011),
            .I(N__27008));
    LocalMux I__4192 (
            .O(N__27008),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__4191 (
            .O(N__27005),
            .I(N__27002));
    InMux I__4190 (
            .O(N__27002),
            .I(N__26999));
    LocalMux I__4189 (
            .O(N__26999),
            .I(N__26996));
    Odrv12 I__4188 (
            .O(N__26996),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    InMux I__4187 (
            .O(N__26993),
            .I(N__26989));
    InMux I__4186 (
            .O(N__26992),
            .I(N__26986));
    LocalMux I__4185 (
            .O(N__26989),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__4184 (
            .O(N__26986),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__4183 (
            .O(N__26981),
            .I(N__26978));
    LocalMux I__4182 (
            .O(N__26978),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__4181 (
            .O(N__26975),
            .I(N__26971));
    InMux I__4180 (
            .O(N__26974),
            .I(N__26968));
    LocalMux I__4179 (
            .O(N__26971),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__4178 (
            .O(N__26968),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__4177 (
            .O(N__26963),
            .I(N__26960));
    InMux I__4176 (
            .O(N__26960),
            .I(N__26957));
    LocalMux I__4175 (
            .O(N__26957),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__4174 (
            .O(N__26954),
            .I(N__26951));
    InMux I__4173 (
            .O(N__26951),
            .I(N__26948));
    LocalMux I__4172 (
            .O(N__26948),
            .I(N__26945));
    Odrv4 I__4171 (
            .O(N__26945),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    InMux I__4170 (
            .O(N__26942),
            .I(N__26938));
    InMux I__4169 (
            .O(N__26941),
            .I(N__26935));
    LocalMux I__4168 (
            .O(N__26938),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__4167 (
            .O(N__26935),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__4166 (
            .O(N__26930),
            .I(N__26927));
    LocalMux I__4165 (
            .O(N__26927),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__4164 (
            .O(N__26924),
            .I(N__26917));
    InMux I__4163 (
            .O(N__26923),
            .I(N__26917));
    InMux I__4162 (
            .O(N__26922),
            .I(N__26914));
    LocalMux I__4161 (
            .O(N__26917),
            .I(N__26911));
    LocalMux I__4160 (
            .O(N__26914),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__4159 (
            .O(N__26911),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    CascadeMux I__4158 (
            .O(N__26906),
            .I(N__26902));
    InMux I__4157 (
            .O(N__26905),
            .I(N__26897));
    InMux I__4156 (
            .O(N__26902),
            .I(N__26897));
    LocalMux I__4155 (
            .O(N__26897),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ));
    CascadeMux I__4154 (
            .O(N__26894),
            .I(N__26890));
    InMux I__4153 (
            .O(N__26893),
            .I(N__26885));
    InMux I__4152 (
            .O(N__26890),
            .I(N__26885));
    LocalMux I__4151 (
            .O(N__26885),
            .I(N__26881));
    InMux I__4150 (
            .O(N__26884),
            .I(N__26878));
    Span4Mux_h I__4149 (
            .O(N__26881),
            .I(N__26875));
    LocalMux I__4148 (
            .O(N__26878),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__4147 (
            .O(N__26875),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__4146 (
            .O(N__26870),
            .I(N__26864));
    InMux I__4145 (
            .O(N__26869),
            .I(N__26864));
    LocalMux I__4144 (
            .O(N__26864),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ));
    CascadeMux I__4143 (
            .O(N__26861),
            .I(N__26858));
    InMux I__4142 (
            .O(N__26858),
            .I(N__26855));
    LocalMux I__4141 (
            .O(N__26855),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    InMux I__4140 (
            .O(N__26852),
            .I(N__26848));
    InMux I__4139 (
            .O(N__26851),
            .I(N__26845));
    LocalMux I__4138 (
            .O(N__26848),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__4137 (
            .O(N__26845),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    CascadeMux I__4136 (
            .O(N__26840),
            .I(N__26837));
    InMux I__4135 (
            .O(N__26837),
            .I(N__26834));
    LocalMux I__4134 (
            .O(N__26834),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    InMux I__4133 (
            .O(N__26831),
            .I(N__26827));
    InMux I__4132 (
            .O(N__26830),
            .I(N__26824));
    LocalMux I__4131 (
            .O(N__26827),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__4130 (
            .O(N__26824),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__4129 (
            .O(N__26819),
            .I(N__26816));
    InMux I__4128 (
            .O(N__26816),
            .I(N__26813));
    LocalMux I__4127 (
            .O(N__26813),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__4126 (
            .O(N__26810),
            .I(N__26806));
    InMux I__4125 (
            .O(N__26809),
            .I(N__26803));
    LocalMux I__4124 (
            .O(N__26806),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__4123 (
            .O(N__26803),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    CascadeMux I__4122 (
            .O(N__26798),
            .I(N__26795));
    InMux I__4121 (
            .O(N__26795),
            .I(N__26792));
    LocalMux I__4120 (
            .O(N__26792),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__4119 (
            .O(N__26789),
            .I(N__26786));
    InMux I__4118 (
            .O(N__26786),
            .I(N__26783));
    LocalMux I__4117 (
            .O(N__26783),
            .I(N__26780));
    Odrv12 I__4116 (
            .O(N__26780),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    InMux I__4115 (
            .O(N__26777),
            .I(N__26773));
    InMux I__4114 (
            .O(N__26776),
            .I(N__26770));
    LocalMux I__4113 (
            .O(N__26773),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__4112 (
            .O(N__26770),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__4111 (
            .O(N__26765),
            .I(N__26762));
    LocalMux I__4110 (
            .O(N__26762),
            .I(N__26759));
    Odrv4 I__4109 (
            .O(N__26759),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__4108 (
            .O(N__26756),
            .I(N__26752));
    InMux I__4107 (
            .O(N__26755),
            .I(N__26749));
    LocalMux I__4106 (
            .O(N__26752),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__4105 (
            .O(N__26749),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__4104 (
            .O(N__26744),
            .I(N__26741));
    InMux I__4103 (
            .O(N__26741),
            .I(N__26738));
    LocalMux I__4102 (
            .O(N__26738),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__4101 (
            .O(N__26735),
            .I(N__26731));
    InMux I__4100 (
            .O(N__26734),
            .I(N__26728));
    LocalMux I__4099 (
            .O(N__26731),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    LocalMux I__4098 (
            .O(N__26728),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    InMux I__4097 (
            .O(N__26723),
            .I(N__26719));
    InMux I__4096 (
            .O(N__26722),
            .I(N__26714));
    LocalMux I__4095 (
            .O(N__26719),
            .I(N__26711));
    InMux I__4094 (
            .O(N__26718),
            .I(N__26706));
    InMux I__4093 (
            .O(N__26717),
            .I(N__26706));
    LocalMux I__4092 (
            .O(N__26714),
            .I(N__26703));
    Odrv4 I__4091 (
            .O(N__26711),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    LocalMux I__4090 (
            .O(N__26706),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    Odrv4 I__4089 (
            .O(N__26703),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    InMux I__4088 (
            .O(N__26696),
            .I(N__26693));
    LocalMux I__4087 (
            .O(N__26693),
            .I(N__26687));
    InMux I__4086 (
            .O(N__26692),
            .I(N__26682));
    InMux I__4085 (
            .O(N__26691),
            .I(N__26682));
    InMux I__4084 (
            .O(N__26690),
            .I(N__26679));
    Odrv4 I__4083 (
            .O(N__26687),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    LocalMux I__4082 (
            .O(N__26682),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    LocalMux I__4081 (
            .O(N__26679),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__4080 (
            .O(N__26672),
            .I(N__26668));
    InMux I__4079 (
            .O(N__26671),
            .I(N__26665));
    LocalMux I__4078 (
            .O(N__26668),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    LocalMux I__4077 (
            .O(N__26665),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    InMux I__4076 (
            .O(N__26660),
            .I(N__26654));
    InMux I__4075 (
            .O(N__26659),
            .I(N__26654));
    LocalMux I__4074 (
            .O(N__26654),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ));
    InMux I__4073 (
            .O(N__26651),
            .I(N__26644));
    InMux I__4072 (
            .O(N__26650),
            .I(N__26644));
    InMux I__4071 (
            .O(N__26649),
            .I(N__26641));
    LocalMux I__4070 (
            .O(N__26644),
            .I(N__26638));
    LocalMux I__4069 (
            .O(N__26641),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__4068 (
            .O(N__26638),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    CascadeMux I__4067 (
            .O(N__26633),
            .I(N__26630));
    InMux I__4066 (
            .O(N__26630),
            .I(N__26623));
    InMux I__4065 (
            .O(N__26629),
            .I(N__26623));
    InMux I__4064 (
            .O(N__26628),
            .I(N__26620));
    LocalMux I__4063 (
            .O(N__26623),
            .I(N__26617));
    LocalMux I__4062 (
            .O(N__26620),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__4061 (
            .O(N__26617),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    CascadeMux I__4060 (
            .O(N__26612),
            .I(N__26609));
    InMux I__4059 (
            .O(N__26609),
            .I(N__26603));
    InMux I__4058 (
            .O(N__26608),
            .I(N__26603));
    LocalMux I__4057 (
            .O(N__26603),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    CascadeMux I__4056 (
            .O(N__26600),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_));
    InMux I__4055 (
            .O(N__26597),
            .I(N__26591));
    InMux I__4054 (
            .O(N__26596),
            .I(N__26591));
    LocalMux I__4053 (
            .O(N__26591),
            .I(N__26588));
    Odrv4 I__4052 (
            .O(N__26588),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__4051 (
            .O(N__26585),
            .I(N__26579));
    InMux I__4050 (
            .O(N__26584),
            .I(N__26579));
    LocalMux I__4049 (
            .O(N__26579),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__4048 (
            .O(N__26576),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_));
    CascadeMux I__4047 (
            .O(N__26573),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ));
    InMux I__4046 (
            .O(N__26570),
            .I(N__26567));
    LocalMux I__4045 (
            .O(N__26567),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ));
    InMux I__4044 (
            .O(N__26564),
            .I(N__26561));
    LocalMux I__4043 (
            .O(N__26561),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ));
    CascadeMux I__4042 (
            .O(N__26558),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_ ));
    InMux I__4041 (
            .O(N__26555),
            .I(N__26552));
    LocalMux I__4040 (
            .O(N__26552),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    InMux I__4039 (
            .O(N__26549),
            .I(N__26546));
    LocalMux I__4038 (
            .O(N__26546),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ));
    InMux I__4037 (
            .O(N__26543),
            .I(N__26540));
    LocalMux I__4036 (
            .O(N__26540),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ));
    InMux I__4035 (
            .O(N__26537),
            .I(N__26534));
    LocalMux I__4034 (
            .O(N__26534),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ));
    CascadeMux I__4033 (
            .O(N__26531),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21_cascade_));
    InMux I__4032 (
            .O(N__26528),
            .I(N__26522));
    InMux I__4031 (
            .O(N__26527),
            .I(N__26522));
    LocalMux I__4030 (
            .O(N__26522),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ));
    CascadeMux I__4029 (
            .O(N__26519),
            .I(N__26515));
    InMux I__4028 (
            .O(N__26518),
            .I(N__26510));
    InMux I__4027 (
            .O(N__26515),
            .I(N__26510));
    LocalMux I__4026 (
            .O(N__26510),
            .I(N__26507));
    Span4Mux_h I__4025 (
            .O(N__26507),
            .I(N__26503));
    InMux I__4024 (
            .O(N__26506),
            .I(N__26500));
    Span4Mux_v I__4023 (
            .O(N__26503),
            .I(N__26497));
    LocalMux I__4022 (
            .O(N__26500),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__4021 (
            .O(N__26497),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__4020 (
            .O(N__26492),
            .I(N__26486));
    InMux I__4019 (
            .O(N__26491),
            .I(N__26486));
    LocalMux I__4018 (
            .O(N__26486),
            .I(N__26482));
    InMux I__4017 (
            .O(N__26485),
            .I(N__26479));
    Span4Mux_v I__4016 (
            .O(N__26482),
            .I(N__26476));
    LocalMux I__4015 (
            .O(N__26479),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__4014 (
            .O(N__26476),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    CascadeMux I__4013 (
            .O(N__26471),
            .I(N__26467));
    InMux I__4012 (
            .O(N__26470),
            .I(N__26462));
    InMux I__4011 (
            .O(N__26467),
            .I(N__26462));
    LocalMux I__4010 (
            .O(N__26462),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ));
    InMux I__4009 (
            .O(N__26459),
            .I(N__26456));
    LocalMux I__4008 (
            .O(N__26456),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ));
    CascadeMux I__4007 (
            .O(N__26453),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ));
    CascadeMux I__4006 (
            .O(N__26450),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    InMux I__4005 (
            .O(N__26447),
            .I(N__26443));
    InMux I__4004 (
            .O(N__26446),
            .I(N__26440));
    LocalMux I__4003 (
            .O(N__26443),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    LocalMux I__4002 (
            .O(N__26440),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__4001 (
            .O(N__26435),
            .I(N__26432));
    LocalMux I__4000 (
            .O(N__26432),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    InMux I__3999 (
            .O(N__26429),
            .I(N__26426));
    LocalMux I__3998 (
            .O(N__26426),
            .I(N__26422));
    InMux I__3997 (
            .O(N__26425),
            .I(N__26419));
    Span4Mux_v I__3996 (
            .O(N__26422),
            .I(N__26416));
    LocalMux I__3995 (
            .O(N__26419),
            .I(N__26413));
    Odrv4 I__3994 (
            .O(N__26416),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ));
    Odrv12 I__3993 (
            .O(N__26413),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ));
    InMux I__3992 (
            .O(N__26408),
            .I(N__26402));
    InMux I__3991 (
            .O(N__26407),
            .I(N__26399));
    InMux I__3990 (
            .O(N__26406),
            .I(N__26396));
    InMux I__3989 (
            .O(N__26405),
            .I(N__26393));
    LocalMux I__3988 (
            .O(N__26402),
            .I(N__26390));
    LocalMux I__3987 (
            .O(N__26399),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__3986 (
            .O(N__26396),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__3985 (
            .O(N__26393),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv12 I__3984 (
            .O(N__26390),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    CEMux I__3983 (
            .O(N__26381),
            .I(N__26376));
    CEMux I__3982 (
            .O(N__26380),
            .I(N__26373));
    CEMux I__3981 (
            .O(N__26379),
            .I(N__26368));
    LocalMux I__3980 (
            .O(N__26376),
            .I(N__26365));
    LocalMux I__3979 (
            .O(N__26373),
            .I(N__26362));
    CEMux I__3978 (
            .O(N__26372),
            .I(N__26359));
    CEMux I__3977 (
            .O(N__26371),
            .I(N__26356));
    LocalMux I__3976 (
            .O(N__26368),
            .I(N__26353));
    Span4Mux_v I__3975 (
            .O(N__26365),
            .I(N__26346));
    Span4Mux_v I__3974 (
            .O(N__26362),
            .I(N__26346));
    LocalMux I__3973 (
            .O(N__26359),
            .I(N__26346));
    LocalMux I__3972 (
            .O(N__26356),
            .I(N__26343));
    Span4Mux_v I__3971 (
            .O(N__26353),
            .I(N__26340));
    Span4Mux_v I__3970 (
            .O(N__26346),
            .I(N__26337));
    Odrv12 I__3969 (
            .O(N__26343),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv4 I__3968 (
            .O(N__26340),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv4 I__3967 (
            .O(N__26337),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    InMux I__3966 (
            .O(N__26330),
            .I(N__26324));
    InMux I__3965 (
            .O(N__26329),
            .I(N__26319));
    InMux I__3964 (
            .O(N__26328),
            .I(N__26319));
    InMux I__3963 (
            .O(N__26327),
            .I(N__26316));
    LocalMux I__3962 (
            .O(N__26324),
            .I(N__26313));
    LocalMux I__3961 (
            .O(N__26319),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__3960 (
            .O(N__26316),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__3959 (
            .O(N__26313),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    CascadeMux I__3958 (
            .O(N__26306),
            .I(N__26303));
    InMux I__3957 (
            .O(N__26303),
            .I(N__26299));
    InMux I__3956 (
            .O(N__26302),
            .I(N__26295));
    LocalMux I__3955 (
            .O(N__26299),
            .I(N__26292));
    InMux I__3954 (
            .O(N__26298),
            .I(N__26289));
    LocalMux I__3953 (
            .O(N__26295),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__3952 (
            .O(N__26292),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__3951 (
            .O(N__26289),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    ClkMux I__3950 (
            .O(N__26282),
            .I(N__26279));
    GlobalMux I__3949 (
            .O(N__26279),
            .I(N__26276));
    gio2CtrlBuf I__3948 (
            .O(N__26276),
            .I(delay_tr_input_c_g));
    InMux I__3947 (
            .O(N__26273),
            .I(N__26270));
    LocalMux I__3946 (
            .O(N__26270),
            .I(N__26265));
    CascadeMux I__3945 (
            .O(N__26269),
            .I(N__26261));
    CascadeMux I__3944 (
            .O(N__26268),
            .I(N__26258));
    Span12Mux_s5_v I__3943 (
            .O(N__26265),
            .I(N__26255));
    InMux I__3942 (
            .O(N__26264),
            .I(N__26252));
    InMux I__3941 (
            .O(N__26261),
            .I(N__26247));
    InMux I__3940 (
            .O(N__26258),
            .I(N__26247));
    Span12Mux_v I__3939 (
            .O(N__26255),
            .I(N__26244));
    LocalMux I__3938 (
            .O(N__26252),
            .I(N__26241));
    LocalMux I__3937 (
            .O(N__26247),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv12 I__3936 (
            .O(N__26244),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__3935 (
            .O(N__26241),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    IoInMux I__3934 (
            .O(N__26234),
            .I(N__26231));
    LocalMux I__3933 (
            .O(N__26231),
            .I(N__26228));
    Odrv4 I__3932 (
            .O(N__26228),
            .I(s3_phy_c));
    InMux I__3931 (
            .O(N__26225),
            .I(N__26222));
    LocalMux I__3930 (
            .O(N__26222),
            .I(N__26219));
    Span4Mux_v I__3929 (
            .O(N__26219),
            .I(N__26214));
    InMux I__3928 (
            .O(N__26218),
            .I(N__26211));
    CascadeMux I__3927 (
            .O(N__26217),
            .I(N__26208));
    Span4Mux_v I__3926 (
            .O(N__26214),
            .I(N__26204));
    LocalMux I__3925 (
            .O(N__26211),
            .I(N__26201));
    InMux I__3924 (
            .O(N__26208),
            .I(N__26198));
    InMux I__3923 (
            .O(N__26207),
            .I(N__26195));
    Span4Mux_v I__3922 (
            .O(N__26204),
            .I(N__26192));
    Span4Mux_h I__3921 (
            .O(N__26201),
            .I(N__26189));
    LocalMux I__3920 (
            .O(N__26198),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__3919 (
            .O(N__26195),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__3918 (
            .O(N__26192),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__3917 (
            .O(N__26189),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    IoInMux I__3916 (
            .O(N__26180),
            .I(N__26177));
    LocalMux I__3915 (
            .O(N__26177),
            .I(N__26174));
    Odrv4 I__3914 (
            .O(N__26174),
            .I(s4_phy_c));
    IoInMux I__3913 (
            .O(N__26171),
            .I(N__26168));
    LocalMux I__3912 (
            .O(N__26168),
            .I(GB_BUFFER_clock_output_0_THRU_CO));
    InMux I__3911 (
            .O(N__26165),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__3910 (
            .O(N__26162),
            .I(bfn_8_14_0_));
    CascadeMux I__3909 (
            .O(N__26159),
            .I(N__26154));
    InMux I__3908 (
            .O(N__26158),
            .I(N__26151));
    InMux I__3907 (
            .O(N__26157),
            .I(N__26146));
    InMux I__3906 (
            .O(N__26154),
            .I(N__26146));
    LocalMux I__3905 (
            .O(N__26151),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__3904 (
            .O(N__26146),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__3903 (
            .O(N__26141),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__3902 (
            .O(N__26138),
            .I(N__26133));
    InMux I__3901 (
            .O(N__26137),
            .I(N__26128));
    InMux I__3900 (
            .O(N__26136),
            .I(N__26128));
    LocalMux I__3899 (
            .O(N__26133),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__3898 (
            .O(N__26128),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__3897 (
            .O(N__26123),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__3896 (
            .O(N__26120),
            .I(N__26115));
    InMux I__3895 (
            .O(N__26119),
            .I(N__26110));
    InMux I__3894 (
            .O(N__26118),
            .I(N__26110));
    LocalMux I__3893 (
            .O(N__26115),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    LocalMux I__3892 (
            .O(N__26110),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__3891 (
            .O(N__26105),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    CascadeMux I__3890 (
            .O(N__26102),
            .I(N__26097));
    InMux I__3889 (
            .O(N__26101),
            .I(N__26094));
    InMux I__3888 (
            .O(N__26100),
            .I(N__26089));
    InMux I__3887 (
            .O(N__26097),
            .I(N__26089));
    LocalMux I__3886 (
            .O(N__26094),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__3885 (
            .O(N__26089),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__3884 (
            .O(N__26084),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__3883 (
            .O(N__26081),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__3882 (
            .O(N__26078),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__3881 (
            .O(N__26075),
            .I(N__26070));
    InMux I__3880 (
            .O(N__26074),
            .I(N__26067));
    InMux I__3879 (
            .O(N__26073),
            .I(N__26064));
    LocalMux I__3878 (
            .O(N__26070),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__3877 (
            .O(N__26067),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__3876 (
            .O(N__26064),
            .I(\phase_controller_inst2.tr_time_passed ));
    InMux I__3875 (
            .O(N__26057),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__3874 (
            .O(N__26054),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__3873 (
            .O(N__26051),
            .I(bfn_8_13_0_));
    InMux I__3872 (
            .O(N__26048),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__3871 (
            .O(N__26045),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__3870 (
            .O(N__26042),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__3869 (
            .O(N__26039),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__3868 (
            .O(N__26036),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__3867 (
            .O(N__26033),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__3866 (
            .O(N__26030),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__3865 (
            .O(N__26027),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__3864 (
            .O(N__26024),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__3863 (
            .O(N__26021),
            .I(bfn_8_12_0_));
    InMux I__3862 (
            .O(N__26018),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__3861 (
            .O(N__26015),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__3860 (
            .O(N__26012),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__3859 (
            .O(N__26009),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__3858 (
            .O(N__26006),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__3857 (
            .O(N__26003),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__3856 (
            .O(N__26000),
            .I(N__25996));
    InMux I__3855 (
            .O(N__25999),
            .I(N__25993));
    LocalMux I__3854 (
            .O(N__25996),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__3853 (
            .O(N__25993),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__3852 (
            .O(N__25988),
            .I(N__25985));
    InMux I__3851 (
            .O(N__25985),
            .I(N__25980));
    InMux I__3850 (
            .O(N__25984),
            .I(N__25977));
    InMux I__3849 (
            .O(N__25983),
            .I(N__25974));
    LocalMux I__3848 (
            .O(N__25980),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__3847 (
            .O(N__25977),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__3846 (
            .O(N__25974),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__3845 (
            .O(N__25967),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__3844 (
            .O(N__25964),
            .I(N__25960));
    InMux I__3843 (
            .O(N__25963),
            .I(N__25957));
    LocalMux I__3842 (
            .O(N__25960),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__3841 (
            .O(N__25957),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__3840 (
            .O(N__25952),
            .I(N__25949));
    InMux I__3839 (
            .O(N__25949),
            .I(N__25944));
    InMux I__3838 (
            .O(N__25948),
            .I(N__25941));
    InMux I__3837 (
            .O(N__25947),
            .I(N__25938));
    LocalMux I__3836 (
            .O(N__25944),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__3835 (
            .O(N__25941),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__3834 (
            .O(N__25938),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__3833 (
            .O(N__25931),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__3832 (
            .O(N__25928),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__3831 (
            .O(N__25925),
            .I(N__25922));
    InMux I__3830 (
            .O(N__25922),
            .I(N__25919));
    LocalMux I__3829 (
            .O(N__25919),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    InMux I__3828 (
            .O(N__25916),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__3827 (
            .O(N__25913),
            .I(N__25910));
    InMux I__3826 (
            .O(N__25910),
            .I(N__25907));
    LocalMux I__3825 (
            .O(N__25907),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ));
    InMux I__3824 (
            .O(N__25904),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__3823 (
            .O(N__25901),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__3822 (
            .O(N__25898),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    CascadeMux I__3821 (
            .O(N__25895),
            .I(N__25892));
    InMux I__3820 (
            .O(N__25892),
            .I(N__25887));
    InMux I__3819 (
            .O(N__25891),
            .I(N__25884));
    InMux I__3818 (
            .O(N__25890),
            .I(N__25881));
    LocalMux I__3817 (
            .O(N__25887),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__3816 (
            .O(N__25884),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__3815 (
            .O(N__25881),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__3814 (
            .O(N__25874),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__3813 (
            .O(N__25871),
            .I(N__25868));
    InMux I__3812 (
            .O(N__25868),
            .I(N__25863));
    InMux I__3811 (
            .O(N__25867),
            .I(N__25860));
    InMux I__3810 (
            .O(N__25866),
            .I(N__25857));
    LocalMux I__3809 (
            .O(N__25863),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__3808 (
            .O(N__25860),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__3807 (
            .O(N__25857),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__3806 (
            .O(N__25850),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__3805 (
            .O(N__25847),
            .I(N__25844));
    InMux I__3804 (
            .O(N__25844),
            .I(N__25839));
    InMux I__3803 (
            .O(N__25843),
            .I(N__25836));
    InMux I__3802 (
            .O(N__25842),
            .I(N__25833));
    LocalMux I__3801 (
            .O(N__25839),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__3800 (
            .O(N__25836),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__3799 (
            .O(N__25833),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__3798 (
            .O(N__25826),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__3797 (
            .O(N__25823),
            .I(N__25820));
    InMux I__3796 (
            .O(N__25820),
            .I(N__25815));
    InMux I__3795 (
            .O(N__25819),
            .I(N__25812));
    InMux I__3794 (
            .O(N__25818),
            .I(N__25809));
    LocalMux I__3793 (
            .O(N__25815),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__3792 (
            .O(N__25812),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__3791 (
            .O(N__25809),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__3790 (
            .O(N__25802),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__3789 (
            .O(N__25799),
            .I(N__25796));
    InMux I__3788 (
            .O(N__25796),
            .I(N__25791));
    InMux I__3787 (
            .O(N__25795),
            .I(N__25788));
    InMux I__3786 (
            .O(N__25794),
            .I(N__25785));
    LocalMux I__3785 (
            .O(N__25791),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__3784 (
            .O(N__25788),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__3783 (
            .O(N__25785),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__3782 (
            .O(N__25778),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__3781 (
            .O(N__25775),
            .I(N__25772));
    InMux I__3780 (
            .O(N__25772),
            .I(N__25767));
    InMux I__3779 (
            .O(N__25771),
            .I(N__25764));
    InMux I__3778 (
            .O(N__25770),
            .I(N__25761));
    LocalMux I__3777 (
            .O(N__25767),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__3776 (
            .O(N__25764),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__3775 (
            .O(N__25761),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__3774 (
            .O(N__25754),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__3773 (
            .O(N__25751),
            .I(N__25748));
    InMux I__3772 (
            .O(N__25748),
            .I(N__25743));
    InMux I__3771 (
            .O(N__25747),
            .I(N__25740));
    InMux I__3770 (
            .O(N__25746),
            .I(N__25737));
    LocalMux I__3769 (
            .O(N__25743),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__3768 (
            .O(N__25740),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__3767 (
            .O(N__25737),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__3766 (
            .O(N__25730),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__3765 (
            .O(N__25727),
            .I(N__25724));
    InMux I__3764 (
            .O(N__25724),
            .I(N__25719));
    InMux I__3763 (
            .O(N__25723),
            .I(N__25716));
    InMux I__3762 (
            .O(N__25722),
            .I(N__25713));
    LocalMux I__3761 (
            .O(N__25719),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__3760 (
            .O(N__25716),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__3759 (
            .O(N__25713),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__3758 (
            .O(N__25706),
            .I(bfn_8_10_0_));
    CascadeMux I__3757 (
            .O(N__25703),
            .I(N__25700));
    InMux I__3756 (
            .O(N__25700),
            .I(N__25695));
    InMux I__3755 (
            .O(N__25699),
            .I(N__25692));
    InMux I__3754 (
            .O(N__25698),
            .I(N__25689));
    LocalMux I__3753 (
            .O(N__25695),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__3752 (
            .O(N__25692),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__3751 (
            .O(N__25689),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    CascadeMux I__3750 (
            .O(N__25682),
            .I(N__25679));
    InMux I__3749 (
            .O(N__25679),
            .I(N__25674));
    InMux I__3748 (
            .O(N__25678),
            .I(N__25671));
    InMux I__3747 (
            .O(N__25677),
            .I(N__25668));
    LocalMux I__3746 (
            .O(N__25674),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__3745 (
            .O(N__25671),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__3744 (
            .O(N__25668),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__3743 (
            .O(N__25661),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__3742 (
            .O(N__25658),
            .I(N__25655));
    InMux I__3741 (
            .O(N__25655),
            .I(N__25650));
    InMux I__3740 (
            .O(N__25654),
            .I(N__25647));
    InMux I__3739 (
            .O(N__25653),
            .I(N__25644));
    LocalMux I__3738 (
            .O(N__25650),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__3737 (
            .O(N__25647),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__3736 (
            .O(N__25644),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__3735 (
            .O(N__25637),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__3734 (
            .O(N__25634),
            .I(N__25631));
    InMux I__3733 (
            .O(N__25631),
            .I(N__25626));
    InMux I__3732 (
            .O(N__25630),
            .I(N__25623));
    InMux I__3731 (
            .O(N__25629),
            .I(N__25620));
    LocalMux I__3730 (
            .O(N__25626),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__3729 (
            .O(N__25623),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__3728 (
            .O(N__25620),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__3727 (
            .O(N__25613),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__3726 (
            .O(N__25610),
            .I(N__25607));
    InMux I__3725 (
            .O(N__25607),
            .I(N__25602));
    InMux I__3724 (
            .O(N__25606),
            .I(N__25599));
    InMux I__3723 (
            .O(N__25605),
            .I(N__25596));
    LocalMux I__3722 (
            .O(N__25602),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__3721 (
            .O(N__25599),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__3720 (
            .O(N__25596),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__3719 (
            .O(N__25589),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__3718 (
            .O(N__25586),
            .I(N__25583));
    InMux I__3717 (
            .O(N__25583),
            .I(N__25578));
    InMux I__3716 (
            .O(N__25582),
            .I(N__25575));
    InMux I__3715 (
            .O(N__25581),
            .I(N__25572));
    LocalMux I__3714 (
            .O(N__25578),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__3713 (
            .O(N__25575),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__3712 (
            .O(N__25572),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__3711 (
            .O(N__25565),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__3710 (
            .O(N__25562),
            .I(N__25559));
    InMux I__3709 (
            .O(N__25559),
            .I(N__25554));
    InMux I__3708 (
            .O(N__25558),
            .I(N__25551));
    InMux I__3707 (
            .O(N__25557),
            .I(N__25548));
    LocalMux I__3706 (
            .O(N__25554),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__3705 (
            .O(N__25551),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__3704 (
            .O(N__25548),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__3703 (
            .O(N__25541),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__3702 (
            .O(N__25538),
            .I(N__25535));
    InMux I__3701 (
            .O(N__25535),
            .I(N__25530));
    InMux I__3700 (
            .O(N__25534),
            .I(N__25527));
    InMux I__3699 (
            .O(N__25533),
            .I(N__25524));
    LocalMux I__3698 (
            .O(N__25530),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__3697 (
            .O(N__25527),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__3696 (
            .O(N__25524),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__3695 (
            .O(N__25517),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__3694 (
            .O(N__25514),
            .I(N__25511));
    InMux I__3693 (
            .O(N__25511),
            .I(N__25506));
    InMux I__3692 (
            .O(N__25510),
            .I(N__25503));
    InMux I__3691 (
            .O(N__25509),
            .I(N__25500));
    LocalMux I__3690 (
            .O(N__25506),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__3689 (
            .O(N__25503),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__3688 (
            .O(N__25500),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__3687 (
            .O(N__25493),
            .I(bfn_8_9_0_));
    CascadeMux I__3686 (
            .O(N__25490),
            .I(N__25486));
    InMux I__3685 (
            .O(N__25489),
            .I(N__25482));
    InMux I__3684 (
            .O(N__25486),
            .I(N__25479));
    InMux I__3683 (
            .O(N__25485),
            .I(N__25476));
    LocalMux I__3682 (
            .O(N__25482),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__3681 (
            .O(N__25479),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__3680 (
            .O(N__25476),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    CascadeMux I__3679 (
            .O(N__25469),
            .I(N__25465));
    InMux I__3678 (
            .O(N__25468),
            .I(N__25461));
    InMux I__3677 (
            .O(N__25465),
            .I(N__25458));
    InMux I__3676 (
            .O(N__25464),
            .I(N__25455));
    LocalMux I__3675 (
            .O(N__25461),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__3674 (
            .O(N__25458),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__3673 (
            .O(N__25455),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__3672 (
            .O(N__25448),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__3671 (
            .O(N__25445),
            .I(N__25442));
    InMux I__3670 (
            .O(N__25442),
            .I(N__25437));
    InMux I__3669 (
            .O(N__25441),
            .I(N__25434));
    InMux I__3668 (
            .O(N__25440),
            .I(N__25431));
    LocalMux I__3667 (
            .O(N__25437),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__3666 (
            .O(N__25434),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__3665 (
            .O(N__25431),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__3664 (
            .O(N__25424),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__3663 (
            .O(N__25421),
            .I(N__25418));
    InMux I__3662 (
            .O(N__25418),
            .I(N__25413));
    InMux I__3661 (
            .O(N__25417),
            .I(N__25410));
    InMux I__3660 (
            .O(N__25416),
            .I(N__25407));
    LocalMux I__3659 (
            .O(N__25413),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__3658 (
            .O(N__25410),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__3657 (
            .O(N__25407),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__3656 (
            .O(N__25400),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__3655 (
            .O(N__25397),
            .I(N__25394));
    InMux I__3654 (
            .O(N__25394),
            .I(N__25389));
    InMux I__3653 (
            .O(N__25393),
            .I(N__25386));
    InMux I__3652 (
            .O(N__25392),
            .I(N__25383));
    LocalMux I__3651 (
            .O(N__25389),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__3650 (
            .O(N__25386),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__3649 (
            .O(N__25383),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__3648 (
            .O(N__25376),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__3647 (
            .O(N__25373),
            .I(N__25370));
    InMux I__3646 (
            .O(N__25370),
            .I(N__25365));
    InMux I__3645 (
            .O(N__25369),
            .I(N__25362));
    InMux I__3644 (
            .O(N__25368),
            .I(N__25359));
    LocalMux I__3643 (
            .O(N__25365),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__3642 (
            .O(N__25362),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__3641 (
            .O(N__25359),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__3640 (
            .O(N__25352),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__3639 (
            .O(N__25349),
            .I(N__25346));
    InMux I__3638 (
            .O(N__25346),
            .I(N__25341));
    InMux I__3637 (
            .O(N__25345),
            .I(N__25338));
    InMux I__3636 (
            .O(N__25344),
            .I(N__25335));
    LocalMux I__3635 (
            .O(N__25341),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__3634 (
            .O(N__25338),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__3633 (
            .O(N__25335),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__3632 (
            .O(N__25328),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__3631 (
            .O(N__25325),
            .I(N__25322));
    InMux I__3630 (
            .O(N__25322),
            .I(N__25317));
    InMux I__3629 (
            .O(N__25321),
            .I(N__25314));
    InMux I__3628 (
            .O(N__25320),
            .I(N__25311));
    LocalMux I__3627 (
            .O(N__25317),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__3626 (
            .O(N__25314),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__3625 (
            .O(N__25311),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__3624 (
            .O(N__25304),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__3623 (
            .O(N__25301),
            .I(N__25298));
    InMux I__3622 (
            .O(N__25298),
            .I(N__25293));
    InMux I__3621 (
            .O(N__25297),
            .I(N__25290));
    InMux I__3620 (
            .O(N__25296),
            .I(N__25287));
    LocalMux I__3619 (
            .O(N__25293),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__3618 (
            .O(N__25290),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__3617 (
            .O(N__25287),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__3616 (
            .O(N__25280),
            .I(bfn_8_8_0_));
    InMux I__3615 (
            .O(N__25277),
            .I(N__25272));
    InMux I__3614 (
            .O(N__25276),
            .I(N__25269));
    InMux I__3613 (
            .O(N__25275),
            .I(N__25266));
    LocalMux I__3612 (
            .O(N__25272),
            .I(N__25259));
    LocalMux I__3611 (
            .O(N__25269),
            .I(N__25259));
    LocalMux I__3610 (
            .O(N__25266),
            .I(N__25259));
    Span12Mux_v I__3609 (
            .O(N__25259),
            .I(N__25256));
    Odrv12 I__3608 (
            .O(N__25256),
            .I(il_min_comp2_c));
    InMux I__3607 (
            .O(N__25253),
            .I(N__25249));
    InMux I__3606 (
            .O(N__25252),
            .I(N__25246));
    LocalMux I__3605 (
            .O(N__25249),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__3604 (
            .O(N__25246),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    CascadeMux I__3603 (
            .O(N__25241),
            .I(N__25238));
    InMux I__3602 (
            .O(N__25238),
            .I(N__25232));
    InMux I__3601 (
            .O(N__25237),
            .I(N__25232));
    LocalMux I__3600 (
            .O(N__25232),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ));
    CascadeMux I__3599 (
            .O(N__25229),
            .I(N__25225));
    InMux I__3598 (
            .O(N__25228),
            .I(N__25220));
    InMux I__3597 (
            .O(N__25225),
            .I(N__25220));
    LocalMux I__3596 (
            .O(N__25220),
            .I(N__25217));
    Span4Mux_v I__3595 (
            .O(N__25217),
            .I(N__25214));
    Span4Mux_v I__3594 (
            .O(N__25214),
            .I(N__25211));
    Odrv4 I__3593 (
            .O(N__25211),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    InMux I__3592 (
            .O(N__25208),
            .I(N__25202));
    InMux I__3591 (
            .O(N__25207),
            .I(N__25202));
    LocalMux I__3590 (
            .O(N__25202),
            .I(N__25199));
    Span4Mux_h I__3589 (
            .O(N__25199),
            .I(N__25196));
    Odrv4 I__3588 (
            .O(N__25196),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    InMux I__3587 (
            .O(N__25193),
            .I(N__25190));
    LocalMux I__3586 (
            .O(N__25190),
            .I(N__25187));
    Span4Mux_h I__3585 (
            .O(N__25187),
            .I(N__25182));
    InMux I__3584 (
            .O(N__25186),
            .I(N__25177));
    InMux I__3583 (
            .O(N__25185),
            .I(N__25177));
    Span4Mux_v I__3582 (
            .O(N__25182),
            .I(N__25174));
    LocalMux I__3581 (
            .O(N__25177),
            .I(N__25171));
    Sp12to4 I__3580 (
            .O(N__25174),
            .I(N__25166));
    Span12Mux_h I__3579 (
            .O(N__25171),
            .I(N__25166));
    Span12Mux_v I__3578 (
            .O(N__25166),
            .I(N__25163));
    Odrv12 I__3577 (
            .O(N__25163),
            .I(il_max_comp2_c));
    CEMux I__3576 (
            .O(N__25160),
            .I(N__25157));
    LocalMux I__3575 (
            .O(N__25157),
            .I(N__25153));
    CEMux I__3574 (
            .O(N__25156),
            .I(N__25150));
    Span4Mux_h I__3573 (
            .O(N__25153),
            .I(N__25143));
    LocalMux I__3572 (
            .O(N__25150),
            .I(N__25143));
    CEMux I__3571 (
            .O(N__25149),
            .I(N__25140));
    CEMux I__3570 (
            .O(N__25148),
            .I(N__25137));
    Span4Mux_v I__3569 (
            .O(N__25143),
            .I(N__25134));
    LocalMux I__3568 (
            .O(N__25140),
            .I(N__25129));
    LocalMux I__3567 (
            .O(N__25137),
            .I(N__25129));
    Span4Mux_h I__3566 (
            .O(N__25134),
            .I(N__25124));
    Span4Mux_v I__3565 (
            .O(N__25129),
            .I(N__25124));
    Odrv4 I__3564 (
            .O(N__25124),
            .I(\delay_measurement_inst.delay_tr_timer.N_201_i ));
    InMux I__3563 (
            .O(N__25121),
            .I(N__25115));
    InMux I__3562 (
            .O(N__25120),
            .I(N__25115));
    LocalMux I__3561 (
            .O(N__25115),
            .I(N__25112));
    Odrv4 I__3560 (
            .O(N__25112),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    InMux I__3559 (
            .O(N__25109),
            .I(N__25103));
    InMux I__3558 (
            .O(N__25108),
            .I(N__25103));
    LocalMux I__3557 (
            .O(N__25103),
            .I(N__25092));
    InMux I__3556 (
            .O(N__25102),
            .I(N__25083));
    InMux I__3555 (
            .O(N__25101),
            .I(N__25083));
    InMux I__3554 (
            .O(N__25100),
            .I(N__25083));
    InMux I__3553 (
            .O(N__25099),
            .I(N__25083));
    InMux I__3552 (
            .O(N__25098),
            .I(N__25054));
    InMux I__3551 (
            .O(N__25097),
            .I(N__25054));
    InMux I__3550 (
            .O(N__25096),
            .I(N__25054));
    InMux I__3549 (
            .O(N__25095),
            .I(N__25054));
    Span4Mux_v I__3548 (
            .O(N__25092),
            .I(N__25049));
    LocalMux I__3547 (
            .O(N__25083),
            .I(N__25049));
    InMux I__3546 (
            .O(N__25082),
            .I(N__25040));
    InMux I__3545 (
            .O(N__25081),
            .I(N__25040));
    InMux I__3544 (
            .O(N__25080),
            .I(N__25040));
    InMux I__3543 (
            .O(N__25079),
            .I(N__25040));
    InMux I__3542 (
            .O(N__25078),
            .I(N__25031));
    InMux I__3541 (
            .O(N__25077),
            .I(N__25031));
    InMux I__3540 (
            .O(N__25076),
            .I(N__25031));
    InMux I__3539 (
            .O(N__25075),
            .I(N__25031));
    InMux I__3538 (
            .O(N__25074),
            .I(N__25022));
    InMux I__3537 (
            .O(N__25073),
            .I(N__25022));
    InMux I__3536 (
            .O(N__25072),
            .I(N__25022));
    InMux I__3535 (
            .O(N__25071),
            .I(N__25022));
    InMux I__3534 (
            .O(N__25070),
            .I(N__25013));
    InMux I__3533 (
            .O(N__25069),
            .I(N__25013));
    InMux I__3532 (
            .O(N__25068),
            .I(N__25013));
    InMux I__3531 (
            .O(N__25067),
            .I(N__25013));
    InMux I__3530 (
            .O(N__25066),
            .I(N__25004));
    InMux I__3529 (
            .O(N__25065),
            .I(N__25004));
    InMux I__3528 (
            .O(N__25064),
            .I(N__25004));
    InMux I__3527 (
            .O(N__25063),
            .I(N__25004));
    LocalMux I__3526 (
            .O(N__25054),
            .I(N__24997));
    Span4Mux_h I__3525 (
            .O(N__25049),
            .I(N__24997));
    LocalMux I__3524 (
            .O(N__25040),
            .I(N__24997));
    LocalMux I__3523 (
            .O(N__25031),
            .I(N__24988));
    LocalMux I__3522 (
            .O(N__25022),
            .I(N__24988));
    LocalMux I__3521 (
            .O(N__25013),
            .I(N__24988));
    LocalMux I__3520 (
            .O(N__25004),
            .I(N__24988));
    Odrv4 I__3519 (
            .O(N__24997),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv12 I__3518 (
            .O(N__24988),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__3517 (
            .O(N__24983),
            .I(N__24980));
    LocalMux I__3516 (
            .O(N__24980),
            .I(\phase_controller_inst2.start_timer_tr_RNO_0_0 ));
    CascadeMux I__3515 (
            .O(N__24977),
            .I(N__24971));
    InMux I__3514 (
            .O(N__24976),
            .I(N__24968));
    InMux I__3513 (
            .O(N__24975),
            .I(N__24963));
    InMux I__3512 (
            .O(N__24974),
            .I(N__24963));
    InMux I__3511 (
            .O(N__24971),
            .I(N__24960));
    LocalMux I__3510 (
            .O(N__24968),
            .I(N__24957));
    LocalMux I__3509 (
            .O(N__24963),
            .I(\phase_controller_inst2.hc_time_passed ));
    LocalMux I__3508 (
            .O(N__24960),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__3507 (
            .O(N__24957),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__3506 (
            .O(N__24950),
            .I(N__24946));
    InMux I__3505 (
            .O(N__24949),
            .I(N__24942));
    LocalMux I__3504 (
            .O(N__24946),
            .I(N__24939));
    InMux I__3503 (
            .O(N__24945),
            .I(N__24936));
    LocalMux I__3502 (
            .O(N__24942),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    Odrv4 I__3501 (
            .O(N__24939),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__3500 (
            .O(N__24936),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__3499 (
            .O(N__24929),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__3498 (
            .O(N__24926),
            .I(bfn_7_10_0_));
    InMux I__3497 (
            .O(N__24923),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__3496 (
            .O(N__24920),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__3495 (
            .O(N__24917),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__3494 (
            .O(N__24914),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__3493 (
            .O(N__24911),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__3492 (
            .O(N__24908),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__3491 (
            .O(N__24905),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__3490 (
            .O(N__24902),
            .I(bfn_7_9_0_));
    InMux I__3489 (
            .O(N__24899),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__3488 (
            .O(N__24896),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__3487 (
            .O(N__24893),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__3486 (
            .O(N__24890),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__3485 (
            .O(N__24887),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__3484 (
            .O(N__24884),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__3483 (
            .O(N__24881),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__3482 (
            .O(N__24878),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__3481 (
            .O(N__24875),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__3480 (
            .O(N__24872),
            .I(bfn_7_8_0_));
    InMux I__3479 (
            .O(N__24869),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__3478 (
            .O(N__24866),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__3477 (
            .O(N__24863),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__3476 (
            .O(N__24860),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__3475 (
            .O(N__24857),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__3474 (
            .O(N__24854),
            .I(N__24849));
    InMux I__3473 (
            .O(N__24853),
            .I(N__24846));
    InMux I__3472 (
            .O(N__24852),
            .I(N__24843));
    LocalMux I__3471 (
            .O(N__24849),
            .I(N__24840));
    LocalMux I__3470 (
            .O(N__24846),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__3469 (
            .O(N__24843),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv12 I__3468 (
            .O(N__24840),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__3467 (
            .O(N__24833),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__3466 (
            .O(N__24830),
            .I(N__24825));
    InMux I__3465 (
            .O(N__24829),
            .I(N__24822));
    InMux I__3464 (
            .O(N__24828),
            .I(N__24819));
    LocalMux I__3463 (
            .O(N__24825),
            .I(N__24816));
    LocalMux I__3462 (
            .O(N__24822),
            .I(N__24813));
    LocalMux I__3461 (
            .O(N__24819),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__3460 (
            .O(N__24816),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__3459 (
            .O(N__24813),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__3458 (
            .O(N__24806),
            .I(bfn_5_27_0_));
    InMux I__3457 (
            .O(N__24803),
            .I(N__24785));
    InMux I__3456 (
            .O(N__24802),
            .I(N__24785));
    InMux I__3455 (
            .O(N__24801),
            .I(N__24785));
    InMux I__3454 (
            .O(N__24800),
            .I(N__24785));
    InMux I__3453 (
            .O(N__24799),
            .I(N__24780));
    InMux I__3452 (
            .O(N__24798),
            .I(N__24780));
    InMux I__3451 (
            .O(N__24797),
            .I(N__24771));
    InMux I__3450 (
            .O(N__24796),
            .I(N__24771));
    InMux I__3449 (
            .O(N__24795),
            .I(N__24771));
    InMux I__3448 (
            .O(N__24794),
            .I(N__24771));
    LocalMux I__3447 (
            .O(N__24785),
            .I(N__24766));
    LocalMux I__3446 (
            .O(N__24780),
            .I(N__24766));
    LocalMux I__3445 (
            .O(N__24771),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__3444 (
            .O(N__24766),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__3443 (
            .O(N__24761),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__3442 (
            .O(N__24758),
            .I(N__24753));
    InMux I__3441 (
            .O(N__24757),
            .I(N__24750));
    InMux I__3440 (
            .O(N__24756),
            .I(N__24747));
    LocalMux I__3439 (
            .O(N__24753),
            .I(N__24744));
    LocalMux I__3438 (
            .O(N__24750),
            .I(N__24741));
    LocalMux I__3437 (
            .O(N__24747),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__3436 (
            .O(N__24744),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__3435 (
            .O(N__24741),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__3434 (
            .O(N__24734),
            .I(bfn_7_7_0_));
    InMux I__3433 (
            .O(N__24731),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__3432 (
            .O(N__24728),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__3431 (
            .O(N__24725),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__3430 (
            .O(N__24722),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    CascadeMux I__3429 (
            .O(N__24719),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__3428 (
            .O(N__24716),
            .I(N__24713));
    LocalMux I__3427 (
            .O(N__24713),
            .I(\pwm_generator_inst.un1_counterlt9 ));
    InMux I__3426 (
            .O(N__24710),
            .I(N__24706));
    InMux I__3425 (
            .O(N__24709),
            .I(N__24702));
    LocalMux I__3424 (
            .O(N__24706),
            .I(N__24699));
    InMux I__3423 (
            .O(N__24705),
            .I(N__24696));
    LocalMux I__3422 (
            .O(N__24702),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__3421 (
            .O(N__24699),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__3420 (
            .O(N__24696),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__3419 (
            .O(N__24689),
            .I(bfn_5_26_0_));
    InMux I__3418 (
            .O(N__24686),
            .I(N__24681));
    InMux I__3417 (
            .O(N__24685),
            .I(N__24678));
    InMux I__3416 (
            .O(N__24684),
            .I(N__24675));
    LocalMux I__3415 (
            .O(N__24681),
            .I(N__24672));
    LocalMux I__3414 (
            .O(N__24678),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__3413 (
            .O(N__24675),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__3412 (
            .O(N__24672),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__3411 (
            .O(N__24665),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__3410 (
            .O(N__24662),
            .I(N__24658));
    InMux I__3409 (
            .O(N__24661),
            .I(N__24654));
    LocalMux I__3408 (
            .O(N__24658),
            .I(N__24651));
    InMux I__3407 (
            .O(N__24657),
            .I(N__24648));
    LocalMux I__3406 (
            .O(N__24654),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__3405 (
            .O(N__24651),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__3404 (
            .O(N__24648),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__3403 (
            .O(N__24641),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__3402 (
            .O(N__24638),
            .I(N__24633));
    InMux I__3401 (
            .O(N__24637),
            .I(N__24630));
    InMux I__3400 (
            .O(N__24636),
            .I(N__24627));
    LocalMux I__3399 (
            .O(N__24633),
            .I(N__24624));
    LocalMux I__3398 (
            .O(N__24630),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__3397 (
            .O(N__24627),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__3396 (
            .O(N__24624),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__3395 (
            .O(N__24617),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__3394 (
            .O(N__24614),
            .I(N__24609));
    InMux I__3393 (
            .O(N__24613),
            .I(N__24606));
    InMux I__3392 (
            .O(N__24612),
            .I(N__24603));
    LocalMux I__3391 (
            .O(N__24609),
            .I(N__24600));
    LocalMux I__3390 (
            .O(N__24606),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__3389 (
            .O(N__24603),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__3388 (
            .O(N__24600),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__3387 (
            .O(N__24593),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__3386 (
            .O(N__24590),
            .I(N__24585));
    InMux I__3385 (
            .O(N__24589),
            .I(N__24582));
    InMux I__3384 (
            .O(N__24588),
            .I(N__24579));
    LocalMux I__3383 (
            .O(N__24585),
            .I(N__24576));
    LocalMux I__3382 (
            .O(N__24582),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__3381 (
            .O(N__24579),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__3380 (
            .O(N__24576),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__3379 (
            .O(N__24569),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__3378 (
            .O(N__24566),
            .I(N__24561));
    InMux I__3377 (
            .O(N__24565),
            .I(N__24558));
    InMux I__3376 (
            .O(N__24564),
            .I(N__24555));
    LocalMux I__3375 (
            .O(N__24561),
            .I(N__24552));
    LocalMux I__3374 (
            .O(N__24558),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__3373 (
            .O(N__24555),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv12 I__3372 (
            .O(N__24552),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__3371 (
            .O(N__24545),
            .I(\pwm_generator_inst.counter_cry_5 ));
    CascadeMux I__3370 (
            .O(N__24542),
            .I(N__24539));
    InMux I__3369 (
            .O(N__24539),
            .I(N__24536));
    LocalMux I__3368 (
            .O(N__24536),
            .I(\pwm_generator_inst.un14_counter_6 ));
    InMux I__3367 (
            .O(N__24533),
            .I(N__24530));
    LocalMux I__3366 (
            .O(N__24530),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__3365 (
            .O(N__24527),
            .I(N__24524));
    LocalMux I__3364 (
            .O(N__24524),
            .I(\pwm_generator_inst.un14_counter_7 ));
    CascadeMux I__3363 (
            .O(N__24521),
            .I(N__24518));
    InMux I__3362 (
            .O(N__24518),
            .I(N__24515));
    LocalMux I__3361 (
            .O(N__24515),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__3360 (
            .O(N__24512),
            .I(N__24509));
    InMux I__3359 (
            .O(N__24509),
            .I(N__24506));
    LocalMux I__3358 (
            .O(N__24506),
            .I(\pwm_generator_inst.un14_counter_8 ));
    InMux I__3357 (
            .O(N__24503),
            .I(N__24500));
    LocalMux I__3356 (
            .O(N__24500),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__3355 (
            .O(N__24497),
            .I(N__24494));
    InMux I__3354 (
            .O(N__24494),
            .I(N__24491));
    LocalMux I__3353 (
            .O(N__24491),
            .I(N__24488));
    Odrv4 I__3352 (
            .O(N__24488),
            .I(\pwm_generator_inst.threshold_9 ));
    InMux I__3351 (
            .O(N__24485),
            .I(N__24482));
    LocalMux I__3350 (
            .O(N__24482),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__3349 (
            .O(N__24479),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__3348 (
            .O(N__24476),
            .I(N__24473));
    LocalMux I__3347 (
            .O(N__24473),
            .I(N__24470));
    Span4Mux_s1_v I__3346 (
            .O(N__24470),
            .I(N__24467));
    Span4Mux_h I__3345 (
            .O(N__24467),
            .I(N__24464));
    Sp12to4 I__3344 (
            .O(N__24464),
            .I(N__24461));
    Span12Mux_h I__3343 (
            .O(N__24461),
            .I(N__24458));
    Span12Mux_v I__3342 (
            .O(N__24458),
            .I(N__24455));
    Odrv12 I__3341 (
            .O(N__24455),
            .I(pwm_output_c));
    InMux I__3340 (
            .O(N__24452),
            .I(N__24449));
    LocalMux I__3339 (
            .O(N__24449),
            .I(N__24446));
    Span4Mux_s3_v I__3338 (
            .O(N__24446),
            .I(N__24443));
    Span4Mux_h I__3337 (
            .O(N__24443),
            .I(N__24440));
    Odrv4 I__3336 (
            .O(N__24440),
            .I(N_38_i_i));
    CascadeMux I__3335 (
            .O(N__24437),
            .I(\pwm_generator_inst.un1_counterlto9_2_cascade_ ));
    InMux I__3334 (
            .O(N__24434),
            .I(N__24431));
    LocalMux I__3333 (
            .O(N__24431),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__3332 (
            .O(N__24428),
            .I(N__24425));
    LocalMux I__3331 (
            .O(N__24425),
            .I(N__24422));
    Odrv12 I__3330 (
            .O(N__24422),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    CascadeMux I__3329 (
            .O(N__24419),
            .I(N__24416));
    InMux I__3328 (
            .O(N__24416),
            .I(N__24413));
    LocalMux I__3327 (
            .O(N__24413),
            .I(\pwm_generator_inst.threshold_0 ));
    InMux I__3326 (
            .O(N__24410),
            .I(N__24407));
    LocalMux I__3325 (
            .O(N__24407),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__3324 (
            .O(N__24404),
            .I(N__24401));
    InMux I__3323 (
            .O(N__24401),
            .I(N__24398));
    LocalMux I__3322 (
            .O(N__24398),
            .I(\pwm_generator_inst.un14_counter_1 ));
    InMux I__3321 (
            .O(N__24395),
            .I(N__24392));
    LocalMux I__3320 (
            .O(N__24392),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__3319 (
            .O(N__24389),
            .I(N__24386));
    InMux I__3318 (
            .O(N__24386),
            .I(N__24383));
    LocalMux I__3317 (
            .O(N__24383),
            .I(\pwm_generator_inst.threshold_2 ));
    InMux I__3316 (
            .O(N__24380),
            .I(N__24377));
    LocalMux I__3315 (
            .O(N__24377),
            .I(N__24374));
    Odrv4 I__3314 (
            .O(N__24374),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__3313 (
            .O(N__24371),
            .I(N__24368));
    InMux I__3312 (
            .O(N__24368),
            .I(N__24365));
    LocalMux I__3311 (
            .O(N__24365),
            .I(\pwm_generator_inst.threshold_3 ));
    InMux I__3310 (
            .O(N__24362),
            .I(N__24359));
    LocalMux I__3309 (
            .O(N__24359),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__3308 (
            .O(N__24356),
            .I(N__24353));
    LocalMux I__3307 (
            .O(N__24353),
            .I(\pwm_generator_inst.threshold_4 ));
    CascadeMux I__3306 (
            .O(N__24350),
            .I(N__24347));
    InMux I__3305 (
            .O(N__24347),
            .I(N__24344));
    LocalMux I__3304 (
            .O(N__24344),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__3303 (
            .O(N__24341),
            .I(N__24338));
    InMux I__3302 (
            .O(N__24338),
            .I(N__24335));
    LocalMux I__3301 (
            .O(N__24335),
            .I(\pwm_generator_inst.threshold_5 ));
    InMux I__3300 (
            .O(N__24332),
            .I(N__24329));
    LocalMux I__3299 (
            .O(N__24329),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__3298 (
            .O(N__24326),
            .I(N__24323));
    LocalMux I__3297 (
            .O(N__24323),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    CascadeMux I__3296 (
            .O(N__24320),
            .I(N__24317));
    InMux I__3295 (
            .O(N__24317),
            .I(N__24314));
    LocalMux I__3294 (
            .O(N__24314),
            .I(N__24311));
    Odrv4 I__3293 (
            .O(N__24311),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ));
    InMux I__3292 (
            .O(N__24308),
            .I(N__24305));
    LocalMux I__3291 (
            .O(N__24305),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    InMux I__3290 (
            .O(N__24302),
            .I(N__24299));
    LocalMux I__3289 (
            .O(N__24299),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    InMux I__3288 (
            .O(N__24296),
            .I(N__24293));
    LocalMux I__3287 (
            .O(N__24293),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    CascadeMux I__3286 (
            .O(N__24290),
            .I(N__24287));
    InMux I__3285 (
            .O(N__24287),
            .I(N__24284));
    LocalMux I__3284 (
            .O(N__24284),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ));
    InMux I__3283 (
            .O(N__24281),
            .I(N__24278));
    LocalMux I__3282 (
            .O(N__24278),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ));
    InMux I__3281 (
            .O(N__24275),
            .I(N__24272));
    LocalMux I__3280 (
            .O(N__24272),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    InMux I__3279 (
            .O(N__24269),
            .I(N__24266));
    LocalMux I__3278 (
            .O(N__24266),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ));
    CascadeMux I__3277 (
            .O(N__24263),
            .I(N__24260));
    InMux I__3276 (
            .O(N__24260),
            .I(N__24257));
    LocalMux I__3275 (
            .O(N__24257),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__3274 (
            .O(N__24254),
            .I(N__24251));
    InMux I__3273 (
            .O(N__24251),
            .I(N__24248));
    LocalMux I__3272 (
            .O(N__24248),
            .I(N__24245));
    Odrv4 I__3271 (
            .O(N__24245),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__3270 (
            .O(N__24242),
            .I(N__24239));
    LocalMux I__3269 (
            .O(N__24239),
            .I(N__24235));
    InMux I__3268 (
            .O(N__24238),
            .I(N__24232));
    Odrv12 I__3267 (
            .O(N__24235),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    LocalMux I__3266 (
            .O(N__24232),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__3265 (
            .O(N__24227),
            .I(N__24224));
    LocalMux I__3264 (
            .O(N__24224),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__3263 (
            .O(N__24221),
            .I(N__24218));
    LocalMux I__3262 (
            .O(N__24218),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    InMux I__3261 (
            .O(N__24215),
            .I(N__24212));
    LocalMux I__3260 (
            .O(N__24212),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    CascadeMux I__3259 (
            .O(N__24209),
            .I(N__24206));
    InMux I__3258 (
            .O(N__24206),
            .I(N__24203));
    LocalMux I__3257 (
            .O(N__24203),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    InMux I__3256 (
            .O(N__24200),
            .I(N__24197));
    LocalMux I__3255 (
            .O(N__24197),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    CascadeMux I__3254 (
            .O(N__24194),
            .I(N__24191));
    InMux I__3253 (
            .O(N__24191),
            .I(N__24188));
    LocalMux I__3252 (
            .O(N__24188),
            .I(N__24185));
    Odrv4 I__3251 (
            .O(N__24185),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ));
    CascadeMux I__3250 (
            .O(N__24182),
            .I(N__24179));
    InMux I__3249 (
            .O(N__24179),
            .I(N__24176));
    LocalMux I__3248 (
            .O(N__24176),
            .I(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ));
    InMux I__3247 (
            .O(N__24173),
            .I(N__24169));
    InMux I__3246 (
            .O(N__24172),
            .I(N__24166));
    LocalMux I__3245 (
            .O(N__24169),
            .I(N__24160));
    LocalMux I__3244 (
            .O(N__24166),
            .I(N__24160));
    InMux I__3243 (
            .O(N__24165),
            .I(N__24157));
    Span4Mux_h I__3242 (
            .O(N__24160),
            .I(N__24154));
    LocalMux I__3241 (
            .O(N__24157),
            .I(N__24151));
    Odrv4 I__3240 (
            .O(N__24154),
            .I(pwm_duty_input_3));
    Odrv4 I__3239 (
            .O(N__24151),
            .I(pwm_duty_input_3));
    CascadeMux I__3238 (
            .O(N__24146),
            .I(N__24143));
    InMux I__3237 (
            .O(N__24143),
            .I(N__24139));
    InMux I__3236 (
            .O(N__24142),
            .I(N__24136));
    LocalMux I__3235 (
            .O(N__24139),
            .I(N__24130));
    LocalMux I__3234 (
            .O(N__24136),
            .I(N__24130));
    InMux I__3233 (
            .O(N__24135),
            .I(N__24127));
    Span4Mux_h I__3232 (
            .O(N__24130),
            .I(N__24124));
    LocalMux I__3231 (
            .O(N__24127),
            .I(N__24121));
    Odrv4 I__3230 (
            .O(N__24124),
            .I(pwm_duty_input_4));
    Odrv4 I__3229 (
            .O(N__24121),
            .I(pwm_duty_input_4));
    CascadeMux I__3228 (
            .O(N__24116),
            .I(N__24113));
    InMux I__3227 (
            .O(N__24113),
            .I(N__24110));
    LocalMux I__3226 (
            .O(N__24110),
            .I(N__24105));
    InMux I__3225 (
            .O(N__24109),
            .I(N__24102));
    InMux I__3224 (
            .O(N__24108),
            .I(N__24099));
    Span4Mux_h I__3223 (
            .O(N__24105),
            .I(N__24096));
    LocalMux I__3222 (
            .O(N__24102),
            .I(N__24093));
    LocalMux I__3221 (
            .O(N__24099),
            .I(N__24090));
    Odrv4 I__3220 (
            .O(N__24096),
            .I(pwm_duty_input_5));
    Odrv4 I__3219 (
            .O(N__24093),
            .I(pwm_duty_input_5));
    Odrv4 I__3218 (
            .O(N__24090),
            .I(pwm_duty_input_5));
    InMux I__3217 (
            .O(N__24083),
            .I(N__24080));
    LocalMux I__3216 (
            .O(N__24080),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ));
    InMux I__3215 (
            .O(N__24077),
            .I(N__24066));
    InMux I__3214 (
            .O(N__24076),
            .I(N__24049));
    InMux I__3213 (
            .O(N__24075),
            .I(N__24049));
    InMux I__3212 (
            .O(N__24074),
            .I(N__24049));
    InMux I__3211 (
            .O(N__24073),
            .I(N__24049));
    InMux I__3210 (
            .O(N__24072),
            .I(N__24049));
    InMux I__3209 (
            .O(N__24071),
            .I(N__24049));
    InMux I__3208 (
            .O(N__24070),
            .I(N__24049));
    InMux I__3207 (
            .O(N__24069),
            .I(N__24049));
    LocalMux I__3206 (
            .O(N__24066),
            .I(\pwm_generator_inst.N_17 ));
    LocalMux I__3205 (
            .O(N__24049),
            .I(\pwm_generator_inst.N_17 ));
    CascadeMux I__3204 (
            .O(N__24044),
            .I(N__24035));
    CascadeMux I__3203 (
            .O(N__24043),
            .I(N__24030));
    CascadeMux I__3202 (
            .O(N__24042),
            .I(N__24027));
    CascadeMux I__3201 (
            .O(N__24041),
            .I(N__24023));
    InMux I__3200 (
            .O(N__24040),
            .I(N__24020));
    InMux I__3199 (
            .O(N__24039),
            .I(N__24017));
    InMux I__3198 (
            .O(N__24038),
            .I(N__24000));
    InMux I__3197 (
            .O(N__24035),
            .I(N__24000));
    InMux I__3196 (
            .O(N__24034),
            .I(N__24000));
    InMux I__3195 (
            .O(N__24033),
            .I(N__24000));
    InMux I__3194 (
            .O(N__24030),
            .I(N__24000));
    InMux I__3193 (
            .O(N__24027),
            .I(N__24000));
    InMux I__3192 (
            .O(N__24026),
            .I(N__24000));
    InMux I__3191 (
            .O(N__24023),
            .I(N__24000));
    LocalMux I__3190 (
            .O(N__24020),
            .I(\pwm_generator_inst.N_16 ));
    LocalMux I__3189 (
            .O(N__24017),
            .I(\pwm_generator_inst.N_16 ));
    LocalMux I__3188 (
            .O(N__24000),
            .I(\pwm_generator_inst.N_16 ));
    InMux I__3187 (
            .O(N__23993),
            .I(N__23990));
    LocalMux I__3186 (
            .O(N__23990),
            .I(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ));
    CascadeMux I__3185 (
            .O(N__23987),
            .I(\pwm_generator_inst.N_17_cascade_ ));
    InMux I__3184 (
            .O(N__23984),
            .I(N__23980));
    CascadeMux I__3183 (
            .O(N__23983),
            .I(N__23977));
    LocalMux I__3182 (
            .O(N__23980),
            .I(N__23973));
    InMux I__3181 (
            .O(N__23977),
            .I(N__23970));
    InMux I__3180 (
            .O(N__23976),
            .I(N__23967));
    Span4Mux_v I__3179 (
            .O(N__23973),
            .I(N__23964));
    LocalMux I__3178 (
            .O(N__23970),
            .I(N__23961));
    LocalMux I__3177 (
            .O(N__23967),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__3176 (
            .O(N__23964),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__3175 (
            .O(N__23961),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    InMux I__3174 (
            .O(N__23954),
            .I(N__23951));
    LocalMux I__3173 (
            .O(N__23951),
            .I(N__23948));
    Odrv12 I__3172 (
            .O(N__23948),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    CascadeMux I__3171 (
            .O(N__23945),
            .I(N__23942));
    InMux I__3170 (
            .O(N__23942),
            .I(N__23938));
    InMux I__3169 (
            .O(N__23941),
            .I(N__23935));
    LocalMux I__3168 (
            .O(N__23938),
            .I(N__23932));
    LocalMux I__3167 (
            .O(N__23935),
            .I(N__23929));
    Span4Mux_v I__3166 (
            .O(N__23932),
            .I(N__23926));
    Span4Mux_h I__3165 (
            .O(N__23929),
            .I(N__23923));
    Odrv4 I__3164 (
            .O(N__23926),
            .I(\pwm_generator_inst.O_10 ));
    Odrv4 I__3163 (
            .O(N__23923),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__3162 (
            .O(N__23918),
            .I(N__23915));
    LocalMux I__3161 (
            .O(N__23915),
            .I(N__23912));
    Span4Mux_h I__3160 (
            .O(N__23912),
            .I(N__23909));
    Odrv4 I__3159 (
            .O(N__23909),
            .I(\pwm_generator_inst.un19_threshold_axb_0 ));
    InMux I__3158 (
            .O(N__23906),
            .I(N__23903));
    LocalMux I__3157 (
            .O(N__23903),
            .I(N__23900));
    Glb2LocalMux I__3156 (
            .O(N__23900),
            .I(N__23897));
    GlobalMux I__3155 (
            .O(N__23897),
            .I(clk_12mhz));
    IoInMux I__3154 (
            .O(N__23894),
            .I(N__23891));
    LocalMux I__3153 (
            .O(N__23891),
            .I(N__23888));
    IoSpan4Mux I__3152 (
            .O(N__23888),
            .I(N__23885));
    Span4Mux_s0_v I__3151 (
            .O(N__23885),
            .I(N__23882));
    Odrv4 I__3150 (
            .O(N__23882),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__3149 (
            .O(N__23879),
            .I(N__23874));
    InMux I__3148 (
            .O(N__23878),
            .I(N__23860));
    InMux I__3147 (
            .O(N__23877),
            .I(N__23860));
    LocalMux I__3146 (
            .O(N__23874),
            .I(N__23857));
    InMux I__3145 (
            .O(N__23873),
            .I(N__23852));
    InMux I__3144 (
            .O(N__23872),
            .I(N__23852));
    InMux I__3143 (
            .O(N__23871),
            .I(N__23839));
    InMux I__3142 (
            .O(N__23870),
            .I(N__23833));
    InMux I__3141 (
            .O(N__23869),
            .I(N__23830));
    InMux I__3140 (
            .O(N__23868),
            .I(N__23827));
    InMux I__3139 (
            .O(N__23867),
            .I(N__23820));
    InMux I__3138 (
            .O(N__23866),
            .I(N__23820));
    InMux I__3137 (
            .O(N__23865),
            .I(N__23820));
    LocalMux I__3136 (
            .O(N__23860),
            .I(N__23813));
    Span4Mux_h I__3135 (
            .O(N__23857),
            .I(N__23813));
    LocalMux I__3134 (
            .O(N__23852),
            .I(N__23813));
    InMux I__3133 (
            .O(N__23851),
            .I(N__23810));
    InMux I__3132 (
            .O(N__23850),
            .I(N__23805));
    InMux I__3131 (
            .O(N__23849),
            .I(N__23805));
    InMux I__3130 (
            .O(N__23848),
            .I(N__23785));
    InMux I__3129 (
            .O(N__23847),
            .I(N__23785));
    InMux I__3128 (
            .O(N__23846),
            .I(N__23785));
    InMux I__3127 (
            .O(N__23845),
            .I(N__23785));
    InMux I__3126 (
            .O(N__23844),
            .I(N__23785));
    InMux I__3125 (
            .O(N__23843),
            .I(N__23785));
    InMux I__3124 (
            .O(N__23842),
            .I(N__23785));
    LocalMux I__3123 (
            .O(N__23839),
            .I(N__23782));
    InMux I__3122 (
            .O(N__23838),
            .I(N__23775));
    InMux I__3121 (
            .O(N__23837),
            .I(N__23775));
    InMux I__3120 (
            .O(N__23836),
            .I(N__23775));
    LocalMux I__3119 (
            .O(N__23833),
            .I(N__23766));
    LocalMux I__3118 (
            .O(N__23830),
            .I(N__23766));
    LocalMux I__3117 (
            .O(N__23827),
            .I(N__23766));
    LocalMux I__3116 (
            .O(N__23820),
            .I(N__23766));
    Span4Mux_h I__3115 (
            .O(N__23813),
            .I(N__23763));
    LocalMux I__3114 (
            .O(N__23810),
            .I(N__23758));
    LocalMux I__3113 (
            .O(N__23805),
            .I(N__23755));
    InMux I__3112 (
            .O(N__23804),
            .I(N__23752));
    InMux I__3111 (
            .O(N__23803),
            .I(N__23743));
    InMux I__3110 (
            .O(N__23802),
            .I(N__23743));
    InMux I__3109 (
            .O(N__23801),
            .I(N__23743));
    InMux I__3108 (
            .O(N__23800),
            .I(N__23743));
    LocalMux I__3107 (
            .O(N__23785),
            .I(N__23738));
    Span4Mux_h I__3106 (
            .O(N__23782),
            .I(N__23738));
    LocalMux I__3105 (
            .O(N__23775),
            .I(N__23731));
    Span4Mux_v I__3104 (
            .O(N__23766),
            .I(N__23731));
    Span4Mux_v I__3103 (
            .O(N__23763),
            .I(N__23731));
    InMux I__3102 (
            .O(N__23762),
            .I(N__23728));
    InMux I__3101 (
            .O(N__23761),
            .I(N__23725));
    Span4Mux_h I__3100 (
            .O(N__23758),
            .I(N__23718));
    Span4Mux_v I__3099 (
            .O(N__23755),
            .I(N__23718));
    LocalMux I__3098 (
            .O(N__23752),
            .I(N__23718));
    LocalMux I__3097 (
            .O(N__23743),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3096 (
            .O(N__23738),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3095 (
            .O(N__23731),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3094 (
            .O(N__23728),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3093 (
            .O(N__23725),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3092 (
            .O(N__23718),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__3091 (
            .O(N__23705),
            .I(N__23691));
    InMux I__3090 (
            .O(N__23704),
            .I(N__23691));
    InMux I__3089 (
            .O(N__23703),
            .I(N__23691));
    CascadeMux I__3088 (
            .O(N__23702),
            .I(N__23679));
    CascadeMux I__3087 (
            .O(N__23701),
            .I(N__23675));
    InMux I__3086 (
            .O(N__23700),
            .I(N__23668));
    InMux I__3085 (
            .O(N__23699),
            .I(N__23668));
    InMux I__3084 (
            .O(N__23698),
            .I(N__23668));
    LocalMux I__3083 (
            .O(N__23691),
            .I(N__23665));
    InMux I__3082 (
            .O(N__23690),
            .I(N__23662));
    CascadeMux I__3081 (
            .O(N__23689),
            .I(N__23648));
    CascadeMux I__3080 (
            .O(N__23688),
            .I(N__23643));
    InMux I__3079 (
            .O(N__23687),
            .I(N__23640));
    InMux I__3078 (
            .O(N__23686),
            .I(N__23637));
    InMux I__3077 (
            .O(N__23685),
            .I(N__23630));
    InMux I__3076 (
            .O(N__23684),
            .I(N__23630));
    InMux I__3075 (
            .O(N__23683),
            .I(N__23630));
    InMux I__3074 (
            .O(N__23682),
            .I(N__23625));
    InMux I__3073 (
            .O(N__23679),
            .I(N__23625));
    InMux I__3072 (
            .O(N__23678),
            .I(N__23620));
    InMux I__3071 (
            .O(N__23675),
            .I(N__23620));
    LocalMux I__3070 (
            .O(N__23668),
            .I(N__23617));
    Span4Mux_v I__3069 (
            .O(N__23665),
            .I(N__23614));
    LocalMux I__3068 (
            .O(N__23662),
            .I(N__23611));
    InMux I__3067 (
            .O(N__23661),
            .I(N__23608));
    InMux I__3066 (
            .O(N__23660),
            .I(N__23593));
    InMux I__3065 (
            .O(N__23659),
            .I(N__23593));
    InMux I__3064 (
            .O(N__23658),
            .I(N__23593));
    InMux I__3063 (
            .O(N__23657),
            .I(N__23593));
    InMux I__3062 (
            .O(N__23656),
            .I(N__23593));
    InMux I__3061 (
            .O(N__23655),
            .I(N__23593));
    InMux I__3060 (
            .O(N__23654),
            .I(N__23593));
    InMux I__3059 (
            .O(N__23653),
            .I(N__23584));
    InMux I__3058 (
            .O(N__23652),
            .I(N__23584));
    InMux I__3057 (
            .O(N__23651),
            .I(N__23584));
    InMux I__3056 (
            .O(N__23648),
            .I(N__23584));
    InMux I__3055 (
            .O(N__23647),
            .I(N__23577));
    InMux I__3054 (
            .O(N__23646),
            .I(N__23577));
    InMux I__3053 (
            .O(N__23643),
            .I(N__23577));
    LocalMux I__3052 (
            .O(N__23640),
            .I(N__23574));
    LocalMux I__3051 (
            .O(N__23637),
            .I(N__23571));
    LocalMux I__3050 (
            .O(N__23630),
            .I(N__23568));
    LocalMux I__3049 (
            .O(N__23625),
            .I(N__23563));
    LocalMux I__3048 (
            .O(N__23620),
            .I(N__23563));
    Span4Mux_v I__3047 (
            .O(N__23617),
            .I(N__23556));
    Span4Mux_s2_h I__3046 (
            .O(N__23614),
            .I(N__23556));
    Span4Mux_v I__3045 (
            .O(N__23611),
            .I(N__23556));
    LocalMux I__3044 (
            .O(N__23608),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    LocalMux I__3043 (
            .O(N__23593),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    LocalMux I__3042 (
            .O(N__23584),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    LocalMux I__3041 (
            .O(N__23577),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__3040 (
            .O(N__23574),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__3039 (
            .O(N__23571),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__3038 (
            .O(N__23568),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__3037 (
            .O(N__23563),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__3036 (
            .O(N__23556),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    CascadeMux I__3035 (
            .O(N__23537),
            .I(N__23534));
    InMux I__3034 (
            .O(N__23534),
            .I(N__23531));
    LocalMux I__3033 (
            .O(N__23531),
            .I(N__23528));
    Span4Mux_h I__3032 (
            .O(N__23528),
            .I(N__23525));
    Odrv4 I__3031 (
            .O(N__23525),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    CascadeMux I__3030 (
            .O(N__23522),
            .I(N__23496));
    CascadeMux I__3029 (
            .O(N__23521),
            .I(N__23493));
    CascadeMux I__3028 (
            .O(N__23520),
            .I(N__23490));
    CascadeMux I__3027 (
            .O(N__23519),
            .I(N__23487));
    InMux I__3026 (
            .O(N__23518),
            .I(N__23484));
    InMux I__3025 (
            .O(N__23517),
            .I(N__23477));
    InMux I__3024 (
            .O(N__23516),
            .I(N__23477));
    InMux I__3023 (
            .O(N__23515),
            .I(N__23477));
    CascadeMux I__3022 (
            .O(N__23514),
            .I(N__23473));
    CascadeMux I__3021 (
            .O(N__23513),
            .I(N__23470));
    InMux I__3020 (
            .O(N__23512),
            .I(N__23467));
    InMux I__3019 (
            .O(N__23511),
            .I(N__23464));
    InMux I__3018 (
            .O(N__23510),
            .I(N__23461));
    CascadeMux I__3017 (
            .O(N__23509),
            .I(N__23456));
    InMux I__3016 (
            .O(N__23508),
            .I(N__23447));
    InMux I__3015 (
            .O(N__23507),
            .I(N__23447));
    InMux I__3014 (
            .O(N__23506),
            .I(N__23440));
    InMux I__3013 (
            .O(N__23505),
            .I(N__23440));
    InMux I__3012 (
            .O(N__23504),
            .I(N__23440));
    InMux I__3011 (
            .O(N__23503),
            .I(N__23435));
    InMux I__3010 (
            .O(N__23502),
            .I(N__23435));
    InMux I__3009 (
            .O(N__23501),
            .I(N__23420));
    InMux I__3008 (
            .O(N__23500),
            .I(N__23420));
    InMux I__3007 (
            .O(N__23499),
            .I(N__23420));
    InMux I__3006 (
            .O(N__23496),
            .I(N__23420));
    InMux I__3005 (
            .O(N__23493),
            .I(N__23420));
    InMux I__3004 (
            .O(N__23490),
            .I(N__23420));
    InMux I__3003 (
            .O(N__23487),
            .I(N__23420));
    LocalMux I__3002 (
            .O(N__23484),
            .I(N__23415));
    LocalMux I__3001 (
            .O(N__23477),
            .I(N__23415));
    InMux I__3000 (
            .O(N__23476),
            .I(N__23408));
    InMux I__2999 (
            .O(N__23473),
            .I(N__23408));
    InMux I__2998 (
            .O(N__23470),
            .I(N__23408));
    LocalMux I__2997 (
            .O(N__23467),
            .I(N__23401));
    LocalMux I__2996 (
            .O(N__23464),
            .I(N__23401));
    LocalMux I__2995 (
            .O(N__23461),
            .I(N__23401));
    InMux I__2994 (
            .O(N__23460),
            .I(N__23394));
    InMux I__2993 (
            .O(N__23459),
            .I(N__23394));
    InMux I__2992 (
            .O(N__23456),
            .I(N__23394));
    InMux I__2991 (
            .O(N__23455),
            .I(N__23385));
    InMux I__2990 (
            .O(N__23454),
            .I(N__23385));
    InMux I__2989 (
            .O(N__23453),
            .I(N__23385));
    InMux I__2988 (
            .O(N__23452),
            .I(N__23385));
    LocalMux I__2987 (
            .O(N__23447),
            .I(N__23382));
    LocalMux I__2986 (
            .O(N__23440),
            .I(N__23379));
    LocalMux I__2985 (
            .O(N__23435),
            .I(N__23372));
    LocalMux I__2984 (
            .O(N__23420),
            .I(N__23372));
    Span4Mux_h I__2983 (
            .O(N__23415),
            .I(N__23372));
    LocalMux I__2982 (
            .O(N__23408),
            .I(N__23367));
    Span4Mux_v I__2981 (
            .O(N__23401),
            .I(N__23367));
    LocalMux I__2980 (
            .O(N__23394),
            .I(N__23364));
    LocalMux I__2979 (
            .O(N__23385),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2978 (
            .O(N__23382),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2977 (
            .O(N__23379),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2976 (
            .O(N__23372),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2975 (
            .O(N__23367),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv12 I__2974 (
            .O(N__23364),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    CascadeMux I__2973 (
            .O(N__23351),
            .I(N__23346));
    InMux I__2972 (
            .O(N__23350),
            .I(N__23342));
    InMux I__2971 (
            .O(N__23349),
            .I(N__23339));
    InMux I__2970 (
            .O(N__23346),
            .I(N__23336));
    InMux I__2969 (
            .O(N__23345),
            .I(N__23333));
    LocalMux I__2968 (
            .O(N__23342),
            .I(N__23330));
    LocalMux I__2967 (
            .O(N__23339),
            .I(N__23327));
    LocalMux I__2966 (
            .O(N__23336),
            .I(N__23324));
    LocalMux I__2965 (
            .O(N__23333),
            .I(N__23321));
    Span4Mux_v I__2964 (
            .O(N__23330),
            .I(N__23318));
    Span4Mux_v I__2963 (
            .O(N__23327),
            .I(N__23315));
    Span4Mux_v I__2962 (
            .O(N__23324),
            .I(N__23312));
    Span12Mux_v I__2961 (
            .O(N__23321),
            .I(N__23309));
    Odrv4 I__2960 (
            .O(N__23318),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__2959 (
            .O(N__23315),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__2958 (
            .O(N__23312),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv12 I__2957 (
            .O(N__23309),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    CascadeMux I__2956 (
            .O(N__23300),
            .I(N__23297));
    InMux I__2955 (
            .O(N__23297),
            .I(N__23294));
    LocalMux I__2954 (
            .O(N__23294),
            .I(N__23290));
    InMux I__2953 (
            .O(N__23293),
            .I(N__23285));
    Span4Mux_v I__2952 (
            .O(N__23290),
            .I(N__23282));
    InMux I__2951 (
            .O(N__23289),
            .I(N__23279));
    InMux I__2950 (
            .O(N__23288),
            .I(N__23276));
    LocalMux I__2949 (
            .O(N__23285),
            .I(N__23273));
    Odrv4 I__2948 (
            .O(N__23282),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__2947 (
            .O(N__23279),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__2946 (
            .O(N__23276),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__2945 (
            .O(N__23273),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__2944 (
            .O(N__23264),
            .I(N__23260));
    InMux I__2943 (
            .O(N__23263),
            .I(N__23257));
    LocalMux I__2942 (
            .O(N__23260),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    LocalMux I__2941 (
            .O(N__23257),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2940 (
            .O(N__23252),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2939 (
            .O(N__23249),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2938 (
            .O(N__23246),
            .I(N__23243));
    LocalMux I__2937 (
            .O(N__23243),
            .I(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ));
    CascadeMux I__2936 (
            .O(N__23240),
            .I(N__23237));
    InMux I__2935 (
            .O(N__23237),
            .I(N__23234));
    LocalMux I__2934 (
            .O(N__23234),
            .I(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ));
    InMux I__2933 (
            .O(N__23231),
            .I(N__23228));
    LocalMux I__2932 (
            .O(N__23228),
            .I(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ));
    CascadeMux I__2931 (
            .O(N__23225),
            .I(N__23222));
    InMux I__2930 (
            .O(N__23222),
            .I(N__23219));
    LocalMux I__2929 (
            .O(N__23219),
            .I(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ));
    InMux I__2928 (
            .O(N__23216),
            .I(N__23213));
    LocalMux I__2927 (
            .O(N__23213),
            .I(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ));
    CascadeMux I__2926 (
            .O(N__23210),
            .I(N__23207));
    InMux I__2925 (
            .O(N__23207),
            .I(N__23204));
    LocalMux I__2924 (
            .O(N__23204),
            .I(N__23201));
    Odrv4 I__2923 (
            .O(N__23201),
            .I(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ));
    InMux I__2922 (
            .O(N__23198),
            .I(N__23195));
    LocalMux I__2921 (
            .O(N__23195),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ));
    InMux I__2920 (
            .O(N__23192),
            .I(N__23189));
    LocalMux I__2919 (
            .O(N__23189),
            .I(N__23186));
    Odrv12 I__2918 (
            .O(N__23186),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    CascadeMux I__2917 (
            .O(N__23183),
            .I(N__23180));
    InMux I__2916 (
            .O(N__23180),
            .I(N__23176));
    CascadeMux I__2915 (
            .O(N__23179),
            .I(N__23172));
    LocalMux I__2914 (
            .O(N__23176),
            .I(N__23169));
    CascadeMux I__2913 (
            .O(N__23175),
            .I(N__23165));
    InMux I__2912 (
            .O(N__23172),
            .I(N__23162));
    Span4Mux_v I__2911 (
            .O(N__23169),
            .I(N__23159));
    InMux I__2910 (
            .O(N__23168),
            .I(N__23156));
    InMux I__2909 (
            .O(N__23165),
            .I(N__23153));
    LocalMux I__2908 (
            .O(N__23162),
            .I(N__23150));
    Odrv4 I__2907 (
            .O(N__23159),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__2906 (
            .O(N__23156),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__2905 (
            .O(N__23153),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__2904 (
            .O(N__23150),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    CascadeMux I__2903 (
            .O(N__23141),
            .I(N__23138));
    InMux I__2902 (
            .O(N__23138),
            .I(N__23134));
    InMux I__2901 (
            .O(N__23137),
            .I(N__23131));
    LocalMux I__2900 (
            .O(N__23134),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    LocalMux I__2899 (
            .O(N__23131),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2898 (
            .O(N__23126),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    CascadeMux I__2897 (
            .O(N__23123),
            .I(N__23120));
    InMux I__2896 (
            .O(N__23120),
            .I(N__23117));
    LocalMux I__2895 (
            .O(N__23117),
            .I(N__23113));
    InMux I__2894 (
            .O(N__23116),
            .I(N__23108));
    Span4Mux_v I__2893 (
            .O(N__23113),
            .I(N__23105));
    InMux I__2892 (
            .O(N__23112),
            .I(N__23102));
    InMux I__2891 (
            .O(N__23111),
            .I(N__23099));
    LocalMux I__2890 (
            .O(N__23108),
            .I(N__23096));
    Odrv4 I__2889 (
            .O(N__23105),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__2888 (
            .O(N__23102),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__2887 (
            .O(N__23099),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv12 I__2886 (
            .O(N__23096),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__2885 (
            .O(N__23087),
            .I(N__23083));
    InMux I__2884 (
            .O(N__23086),
            .I(N__23078));
    InMux I__2883 (
            .O(N__23083),
            .I(N__23078));
    LocalMux I__2882 (
            .O(N__23078),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2881 (
            .O(N__23075),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    CascadeMux I__2880 (
            .O(N__23072),
            .I(N__23069));
    InMux I__2879 (
            .O(N__23069),
            .I(N__23066));
    LocalMux I__2878 (
            .O(N__23066),
            .I(N__23061));
    InMux I__2877 (
            .O(N__23065),
            .I(N__23057));
    InMux I__2876 (
            .O(N__23064),
            .I(N__23054));
    Span4Mux_v I__2875 (
            .O(N__23061),
            .I(N__23051));
    InMux I__2874 (
            .O(N__23060),
            .I(N__23048));
    LocalMux I__2873 (
            .O(N__23057),
            .I(N__23043));
    LocalMux I__2872 (
            .O(N__23054),
            .I(N__23043));
    Odrv4 I__2871 (
            .O(N__23051),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__2870 (
            .O(N__23048),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv12 I__2869 (
            .O(N__23043),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__2868 (
            .O(N__23036),
            .I(N__23030));
    InMux I__2867 (
            .O(N__23035),
            .I(N__23030));
    LocalMux I__2866 (
            .O(N__23030),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2865 (
            .O(N__23027),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    CascadeMux I__2864 (
            .O(N__23024),
            .I(N__23021));
    InMux I__2863 (
            .O(N__23021),
            .I(N__23017));
    CascadeMux I__2862 (
            .O(N__23020),
            .I(N__23014));
    LocalMux I__2861 (
            .O(N__23017),
            .I(N__23011));
    InMux I__2860 (
            .O(N__23014),
            .I(N__23006));
    Span4Mux_v I__2859 (
            .O(N__23011),
            .I(N__23003));
    InMux I__2858 (
            .O(N__23010),
            .I(N__23000));
    InMux I__2857 (
            .O(N__23009),
            .I(N__22997));
    LocalMux I__2856 (
            .O(N__23006),
            .I(N__22994));
    Odrv4 I__2855 (
            .O(N__23003),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__2854 (
            .O(N__23000),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__2853 (
            .O(N__22997),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__2852 (
            .O(N__22994),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__2851 (
            .O(N__22985),
            .I(N__22979));
    InMux I__2850 (
            .O(N__22984),
            .I(N__22979));
    LocalMux I__2849 (
            .O(N__22979),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2848 (
            .O(N__22976),
            .I(bfn_4_20_0_));
    CascadeMux I__2847 (
            .O(N__22973),
            .I(N__22970));
    InMux I__2846 (
            .O(N__22970),
            .I(N__22966));
    InMux I__2845 (
            .O(N__22969),
            .I(N__22963));
    LocalMux I__2844 (
            .O(N__22966),
            .I(N__22959));
    LocalMux I__2843 (
            .O(N__22963),
            .I(N__22956));
    InMux I__2842 (
            .O(N__22962),
            .I(N__22952));
    Span4Mux_h I__2841 (
            .O(N__22959),
            .I(N__22947));
    Span4Mux_h I__2840 (
            .O(N__22956),
            .I(N__22947));
    InMux I__2839 (
            .O(N__22955),
            .I(N__22944));
    LocalMux I__2838 (
            .O(N__22952),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__2837 (
            .O(N__22947),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__2836 (
            .O(N__22944),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__2835 (
            .O(N__22937),
            .I(N__22931));
    InMux I__2834 (
            .O(N__22936),
            .I(N__22931));
    LocalMux I__2833 (
            .O(N__22931),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2832 (
            .O(N__22928),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    CascadeMux I__2831 (
            .O(N__22925),
            .I(N__22921));
    InMux I__2830 (
            .O(N__22924),
            .I(N__22918));
    InMux I__2829 (
            .O(N__22921),
            .I(N__22915));
    LocalMux I__2828 (
            .O(N__22918),
            .I(N__22912));
    LocalMux I__2827 (
            .O(N__22915),
            .I(N__22908));
    Span4Mux_h I__2826 (
            .O(N__22912),
            .I(N__22904));
    InMux I__2825 (
            .O(N__22911),
            .I(N__22901));
    Span4Mux_h I__2824 (
            .O(N__22908),
            .I(N__22898));
    InMux I__2823 (
            .O(N__22907),
            .I(N__22895));
    Odrv4 I__2822 (
            .O(N__22904),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__2821 (
            .O(N__22901),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__2820 (
            .O(N__22898),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__2819 (
            .O(N__22895),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__2818 (
            .O(N__22886),
            .I(N__22882));
    InMux I__2817 (
            .O(N__22885),
            .I(N__22879));
    LocalMux I__2816 (
            .O(N__22882),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    LocalMux I__2815 (
            .O(N__22879),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2814 (
            .O(N__22874),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2813 (
            .O(N__22871),
            .I(N__22868));
    LocalMux I__2812 (
            .O(N__22868),
            .I(N__22864));
    InMux I__2811 (
            .O(N__22867),
            .I(N__22859));
    Span4Mux_v I__2810 (
            .O(N__22864),
            .I(N__22856));
    InMux I__2809 (
            .O(N__22863),
            .I(N__22853));
    InMux I__2808 (
            .O(N__22862),
            .I(N__22850));
    LocalMux I__2807 (
            .O(N__22859),
            .I(N__22847));
    Odrv4 I__2806 (
            .O(N__22856),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__2805 (
            .O(N__22853),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__2804 (
            .O(N__22850),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__2803 (
            .O(N__22847),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__2802 (
            .O(N__22838),
            .I(N__22832));
    InMux I__2801 (
            .O(N__22837),
            .I(N__22832));
    LocalMux I__2800 (
            .O(N__22832),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2799 (
            .O(N__22829),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2798 (
            .O(N__22826),
            .I(N__22823));
    LocalMux I__2797 (
            .O(N__22823),
            .I(N__22820));
    Span4Mux_v I__2796 (
            .O(N__22820),
            .I(N__22814));
    InMux I__2795 (
            .O(N__22819),
            .I(N__22811));
    InMux I__2794 (
            .O(N__22818),
            .I(N__22808));
    InMux I__2793 (
            .O(N__22817),
            .I(N__22805));
    Odrv4 I__2792 (
            .O(N__22814),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__2791 (
            .O(N__22811),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__2790 (
            .O(N__22808),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__2789 (
            .O(N__22805),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    CascadeMux I__2788 (
            .O(N__22796),
            .I(N__22792));
    CascadeMux I__2787 (
            .O(N__22795),
            .I(N__22789));
    InMux I__2786 (
            .O(N__22792),
            .I(N__22786));
    InMux I__2785 (
            .O(N__22789),
            .I(N__22783));
    LocalMux I__2784 (
            .O(N__22786),
            .I(N__22780));
    LocalMux I__2783 (
            .O(N__22783),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    Odrv4 I__2782 (
            .O(N__22780),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2781 (
            .O(N__22775),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    CascadeMux I__2780 (
            .O(N__22772),
            .I(N__22769));
    InMux I__2779 (
            .O(N__22769),
            .I(N__22766));
    LocalMux I__2778 (
            .O(N__22766),
            .I(N__22761));
    InMux I__2777 (
            .O(N__22765),
            .I(N__22757));
    InMux I__2776 (
            .O(N__22764),
            .I(N__22754));
    Span4Mux_v I__2775 (
            .O(N__22761),
            .I(N__22751));
    InMux I__2774 (
            .O(N__22760),
            .I(N__22748));
    LocalMux I__2773 (
            .O(N__22757),
            .I(N__22743));
    LocalMux I__2772 (
            .O(N__22754),
            .I(N__22743));
    Odrv4 I__2771 (
            .O(N__22751),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__2770 (
            .O(N__22748),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__2769 (
            .O(N__22743),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    CascadeMux I__2768 (
            .O(N__22736),
            .I(N__22733));
    InMux I__2767 (
            .O(N__22733),
            .I(N__22730));
    LocalMux I__2766 (
            .O(N__22730),
            .I(N__22727));
    Span4Mux_v I__2765 (
            .O(N__22727),
            .I(N__22723));
    InMux I__2764 (
            .O(N__22726),
            .I(N__22720));
    Odrv4 I__2763 (
            .O(N__22723),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    LocalMux I__2762 (
            .O(N__22720),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2761 (
            .O(N__22715),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    CascadeMux I__2760 (
            .O(N__22712),
            .I(N__22709));
    InMux I__2759 (
            .O(N__22709),
            .I(N__22706));
    LocalMux I__2758 (
            .O(N__22706),
            .I(N__22701));
    InMux I__2757 (
            .O(N__22705),
            .I(N__22698));
    InMux I__2756 (
            .O(N__22704),
            .I(N__22695));
    Span4Mux_v I__2755 (
            .O(N__22701),
            .I(N__22691));
    LocalMux I__2754 (
            .O(N__22698),
            .I(N__22686));
    LocalMux I__2753 (
            .O(N__22695),
            .I(N__22686));
    InMux I__2752 (
            .O(N__22694),
            .I(N__22683));
    Odrv4 I__2751 (
            .O(N__22691),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__2750 (
            .O(N__22686),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__2749 (
            .O(N__22683),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__2748 (
            .O(N__22676),
            .I(N__22670));
    InMux I__2747 (
            .O(N__22675),
            .I(N__22670));
    LocalMux I__2746 (
            .O(N__22670),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2745 (
            .O(N__22667),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    CascadeMux I__2744 (
            .O(N__22664),
            .I(N__22661));
    InMux I__2743 (
            .O(N__22661),
            .I(N__22657));
    InMux I__2742 (
            .O(N__22660),
            .I(N__22652));
    LocalMux I__2741 (
            .O(N__22657),
            .I(N__22649));
    InMux I__2740 (
            .O(N__22656),
            .I(N__22646));
    InMux I__2739 (
            .O(N__22655),
            .I(N__22643));
    LocalMux I__2738 (
            .O(N__22652),
            .I(N__22640));
    Span4Mux_h I__2737 (
            .O(N__22649),
            .I(N__22631));
    LocalMux I__2736 (
            .O(N__22646),
            .I(N__22631));
    LocalMux I__2735 (
            .O(N__22643),
            .I(N__22631));
    Span4Mux_s3_h I__2734 (
            .O(N__22640),
            .I(N__22631));
    Odrv4 I__2733 (
            .O(N__22631),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__2732 (
            .O(N__22628),
            .I(N__22622));
    InMux I__2731 (
            .O(N__22627),
            .I(N__22622));
    LocalMux I__2730 (
            .O(N__22622),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2729 (
            .O(N__22619),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    CascadeMux I__2728 (
            .O(N__22616),
            .I(N__22613));
    InMux I__2727 (
            .O(N__22613),
            .I(N__22609));
    InMux I__2726 (
            .O(N__22612),
            .I(N__22605));
    LocalMux I__2725 (
            .O(N__22609),
            .I(N__22601));
    InMux I__2724 (
            .O(N__22608),
            .I(N__22598));
    LocalMux I__2723 (
            .O(N__22605),
            .I(N__22595));
    InMux I__2722 (
            .O(N__22604),
            .I(N__22592));
    Span4Mux_v I__2721 (
            .O(N__22601),
            .I(N__22587));
    LocalMux I__2720 (
            .O(N__22598),
            .I(N__22587));
    Span4Mux_h I__2719 (
            .O(N__22595),
            .I(N__22584));
    LocalMux I__2718 (
            .O(N__22592),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__2717 (
            .O(N__22587),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__2716 (
            .O(N__22584),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__2715 (
            .O(N__22577),
            .I(N__22573));
    InMux I__2714 (
            .O(N__22576),
            .I(N__22570));
    LocalMux I__2713 (
            .O(N__22573),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    LocalMux I__2712 (
            .O(N__22570),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2711 (
            .O(N__22565),
            .I(bfn_4_19_0_));
    InMux I__2710 (
            .O(N__22562),
            .I(N__22559));
    LocalMux I__2709 (
            .O(N__22559),
            .I(N__22556));
    Odrv4 I__2708 (
            .O(N__22556),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    CascadeMux I__2707 (
            .O(N__22553),
            .I(N__22550));
    InMux I__2706 (
            .O(N__22550),
            .I(N__22547));
    LocalMux I__2705 (
            .O(N__22547),
            .I(N__22543));
    InMux I__2704 (
            .O(N__22546),
            .I(N__22538));
    Span4Mux_v I__2703 (
            .O(N__22543),
            .I(N__22535));
    InMux I__2702 (
            .O(N__22542),
            .I(N__22532));
    InMux I__2701 (
            .O(N__22541),
            .I(N__22529));
    LocalMux I__2700 (
            .O(N__22538),
            .I(N__22526));
    Odrv4 I__2699 (
            .O(N__22535),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__2698 (
            .O(N__22532),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__2697 (
            .O(N__22529),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__2696 (
            .O(N__22526),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    CascadeMux I__2695 (
            .O(N__22517),
            .I(N__22514));
    InMux I__2694 (
            .O(N__22514),
            .I(N__22510));
    InMux I__2693 (
            .O(N__22513),
            .I(N__22507));
    LocalMux I__2692 (
            .O(N__22510),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    LocalMux I__2691 (
            .O(N__22507),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2690 (
            .O(N__22502),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2689 (
            .O(N__22499),
            .I(N__22496));
    LocalMux I__2688 (
            .O(N__22496),
            .I(N__22491));
    CascadeMux I__2687 (
            .O(N__22495),
            .I(N__22488));
    InMux I__2686 (
            .O(N__22494),
            .I(N__22484));
    Span4Mux_v I__2685 (
            .O(N__22491),
            .I(N__22481));
    InMux I__2684 (
            .O(N__22488),
            .I(N__22478));
    InMux I__2683 (
            .O(N__22487),
            .I(N__22475));
    LocalMux I__2682 (
            .O(N__22484),
            .I(N__22472));
    Odrv4 I__2681 (
            .O(N__22481),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__2680 (
            .O(N__22478),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__2679 (
            .O(N__22475),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__2678 (
            .O(N__22472),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__2677 (
            .O(N__22463),
            .I(N__22457));
    InMux I__2676 (
            .O(N__22462),
            .I(N__22457));
    LocalMux I__2675 (
            .O(N__22457),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2674 (
            .O(N__22454),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2673 (
            .O(N__22451),
            .I(N__22448));
    LocalMux I__2672 (
            .O(N__22448),
            .I(N__22445));
    Odrv12 I__2671 (
            .O(N__22445),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    CascadeMux I__2670 (
            .O(N__22442),
            .I(N__22439));
    InMux I__2669 (
            .O(N__22439),
            .I(N__22436));
    LocalMux I__2668 (
            .O(N__22436),
            .I(N__22432));
    CascadeMux I__2667 (
            .O(N__22435),
            .I(N__22427));
    Span4Mux_h I__2666 (
            .O(N__22432),
            .I(N__22424));
    InMux I__2665 (
            .O(N__22431),
            .I(N__22421));
    InMux I__2664 (
            .O(N__22430),
            .I(N__22418));
    InMux I__2663 (
            .O(N__22427),
            .I(N__22415));
    Sp12to4 I__2662 (
            .O(N__22424),
            .I(N__22408));
    LocalMux I__2661 (
            .O(N__22421),
            .I(N__22408));
    LocalMux I__2660 (
            .O(N__22418),
            .I(N__22408));
    LocalMux I__2659 (
            .O(N__22415),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv12 I__2658 (
            .O(N__22408),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__2657 (
            .O(N__22403),
            .I(N__22399));
    InMux I__2656 (
            .O(N__22402),
            .I(N__22394));
    InMux I__2655 (
            .O(N__22399),
            .I(N__22394));
    LocalMux I__2654 (
            .O(N__22394),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2653 (
            .O(N__22391),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    CascadeMux I__2652 (
            .O(N__22388),
            .I(N__22385));
    InMux I__2651 (
            .O(N__22385),
            .I(N__22381));
    CascadeMux I__2650 (
            .O(N__22384),
            .I(N__22378));
    LocalMux I__2649 (
            .O(N__22381),
            .I(N__22375));
    InMux I__2648 (
            .O(N__22378),
            .I(N__22372));
    Span4Mux_h I__2647 (
            .O(N__22375),
            .I(N__22368));
    LocalMux I__2646 (
            .O(N__22372),
            .I(N__22364));
    InMux I__2645 (
            .O(N__22371),
            .I(N__22361));
    Span4Mux_v I__2644 (
            .O(N__22368),
            .I(N__22358));
    InMux I__2643 (
            .O(N__22367),
            .I(N__22355));
    Span4Mux_v I__2642 (
            .O(N__22364),
            .I(N__22350));
    LocalMux I__2641 (
            .O(N__22361),
            .I(N__22350));
    Odrv4 I__2640 (
            .O(N__22358),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__2639 (
            .O(N__22355),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__2638 (
            .O(N__22350),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__2637 (
            .O(N__22343),
            .I(N__22340));
    LocalMux I__2636 (
            .O(N__22340),
            .I(N__22336));
    InMux I__2635 (
            .O(N__22339),
            .I(N__22333));
    Odrv4 I__2634 (
            .O(N__22336),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    LocalMux I__2633 (
            .O(N__22333),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2632 (
            .O(N__22328),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2631 (
            .O(N__22325),
            .I(N__22322));
    LocalMux I__2630 (
            .O(N__22322),
            .I(N__22319));
    Odrv12 I__2629 (
            .O(N__22319),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__2628 (
            .O(N__22316),
            .I(N__22313));
    InMux I__2627 (
            .O(N__22313),
            .I(N__22310));
    LocalMux I__2626 (
            .O(N__22310),
            .I(N__22305));
    InMux I__2625 (
            .O(N__22309),
            .I(N__22302));
    InMux I__2624 (
            .O(N__22308),
            .I(N__22299));
    Span4Mux_v I__2623 (
            .O(N__22305),
            .I(N__22294));
    LocalMux I__2622 (
            .O(N__22302),
            .I(N__22294));
    LocalMux I__2621 (
            .O(N__22299),
            .I(N__22291));
    Span4Mux_h I__2620 (
            .O(N__22294),
            .I(N__22288));
    Span4Mux_v I__2619 (
            .O(N__22291),
            .I(N__22285));
    Odrv4 I__2618 (
            .O(N__22288),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__2617 (
            .O(N__22285),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2616 (
            .O(N__22280),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__2615 (
            .O(N__22277),
            .I(N__22273));
    InMux I__2614 (
            .O(N__22276),
            .I(N__22270));
    LocalMux I__2613 (
            .O(N__22273),
            .I(N__22266));
    LocalMux I__2612 (
            .O(N__22270),
            .I(N__22263));
    InMux I__2611 (
            .O(N__22269),
            .I(N__22260));
    Span4Mux_v I__2610 (
            .O(N__22266),
            .I(N__22257));
    Span4Mux_v I__2609 (
            .O(N__22263),
            .I(N__22251));
    LocalMux I__2608 (
            .O(N__22260),
            .I(N__22251));
    Span4Mux_h I__2607 (
            .O(N__22257),
            .I(N__22248));
    InMux I__2606 (
            .O(N__22256),
            .I(N__22245));
    Odrv4 I__2605 (
            .O(N__22251),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__2604 (
            .O(N__22248),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__2603 (
            .O(N__22245),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    CascadeMux I__2602 (
            .O(N__22238),
            .I(N__22235));
    InMux I__2601 (
            .O(N__22235),
            .I(N__22230));
    InMux I__2600 (
            .O(N__22234),
            .I(N__22227));
    InMux I__2599 (
            .O(N__22233),
            .I(N__22224));
    LocalMux I__2598 (
            .O(N__22230),
            .I(N__22221));
    LocalMux I__2597 (
            .O(N__22227),
            .I(N__22218));
    LocalMux I__2596 (
            .O(N__22224),
            .I(N__22215));
    Span12Mux_v I__2595 (
            .O(N__22221),
            .I(N__22212));
    Span4Mux_h I__2594 (
            .O(N__22218),
            .I(N__22209));
    Span4Mux_v I__2593 (
            .O(N__22215),
            .I(N__22206));
    Odrv12 I__2592 (
            .O(N__22212),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2591 (
            .O(N__22209),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2590 (
            .O(N__22206),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2589 (
            .O(N__22199),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    InMux I__2588 (
            .O(N__22196),
            .I(N__22191));
    CascadeMux I__2587 (
            .O(N__22195),
            .I(N__22187));
    InMux I__2586 (
            .O(N__22194),
            .I(N__22184));
    LocalMux I__2585 (
            .O(N__22191),
            .I(N__22181));
    CascadeMux I__2584 (
            .O(N__22190),
            .I(N__22178));
    InMux I__2583 (
            .O(N__22187),
            .I(N__22175));
    LocalMux I__2582 (
            .O(N__22184),
            .I(N__22172));
    Span4Mux_v I__2581 (
            .O(N__22181),
            .I(N__22169));
    InMux I__2580 (
            .O(N__22178),
            .I(N__22166));
    LocalMux I__2579 (
            .O(N__22175),
            .I(N__22161));
    Span4Mux_h I__2578 (
            .O(N__22172),
            .I(N__22161));
    Odrv4 I__2577 (
            .O(N__22169),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__2576 (
            .O(N__22166),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__2575 (
            .O(N__22161),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__2574 (
            .O(N__22154),
            .I(N__22150));
    InMux I__2573 (
            .O(N__22153),
            .I(N__22146));
    LocalMux I__2572 (
            .O(N__22150),
            .I(N__22143));
    InMux I__2571 (
            .O(N__22149),
            .I(N__22140));
    LocalMux I__2570 (
            .O(N__22146),
            .I(N__22137));
    Span4Mux_s3_h I__2569 (
            .O(N__22143),
            .I(N__22132));
    LocalMux I__2568 (
            .O(N__22140),
            .I(N__22132));
    Span4Mux_h I__2567 (
            .O(N__22137),
            .I(N__22129));
    Span4Mux_v I__2566 (
            .O(N__22132),
            .I(N__22126));
    Odrv4 I__2565 (
            .O(N__22129),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv4 I__2564 (
            .O(N__22126),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2563 (
            .O(N__22121),
            .I(bfn_4_18_0_));
    InMux I__2562 (
            .O(N__22118),
            .I(N__22115));
    LocalMux I__2561 (
            .O(N__22115),
            .I(N__22112));
    Odrv12 I__2560 (
            .O(N__22112),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    CascadeMux I__2559 (
            .O(N__22109),
            .I(N__22106));
    InMux I__2558 (
            .O(N__22106),
            .I(N__22101));
    CascadeMux I__2557 (
            .O(N__22105),
            .I(N__22098));
    CascadeMux I__2556 (
            .O(N__22104),
            .I(N__22095));
    LocalMux I__2555 (
            .O(N__22101),
            .I(N__22092));
    InMux I__2554 (
            .O(N__22098),
            .I(N__22089));
    InMux I__2553 (
            .O(N__22095),
            .I(N__22086));
    Span4Mux_h I__2552 (
            .O(N__22092),
            .I(N__22081));
    LocalMux I__2551 (
            .O(N__22089),
            .I(N__22081));
    LocalMux I__2550 (
            .O(N__22086),
            .I(N__22078));
    Span4Mux_v I__2549 (
            .O(N__22081),
            .I(N__22074));
    Span12Mux_v I__2548 (
            .O(N__22078),
            .I(N__22071));
    InMux I__2547 (
            .O(N__22077),
            .I(N__22068));
    Odrv4 I__2546 (
            .O(N__22074),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv12 I__2545 (
            .O(N__22071),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__2544 (
            .O(N__22068),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__2543 (
            .O(N__22061),
            .I(N__22055));
    InMux I__2542 (
            .O(N__22060),
            .I(N__22055));
    LocalMux I__2541 (
            .O(N__22055),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2540 (
            .O(N__22052),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2539 (
            .O(N__22049),
            .I(N__22046));
    LocalMux I__2538 (
            .O(N__22046),
            .I(N__22043));
    Odrv12 I__2537 (
            .O(N__22043),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__2536 (
            .O(N__22040),
            .I(N__22036));
    CascadeMux I__2535 (
            .O(N__22039),
            .I(N__22033));
    InMux I__2534 (
            .O(N__22036),
            .I(N__22029));
    InMux I__2533 (
            .O(N__22033),
            .I(N__22026));
    InMux I__2532 (
            .O(N__22032),
            .I(N__22023));
    LocalMux I__2531 (
            .O(N__22029),
            .I(N__22019));
    LocalMux I__2530 (
            .O(N__22026),
            .I(N__22016));
    LocalMux I__2529 (
            .O(N__22023),
            .I(N__22013));
    InMux I__2528 (
            .O(N__22022),
            .I(N__22010));
    Span4Mux_v I__2527 (
            .O(N__22019),
            .I(N__22007));
    Span4Mux_v I__2526 (
            .O(N__22016),
            .I(N__22002));
    Span4Mux_s3_h I__2525 (
            .O(N__22013),
            .I(N__22002));
    LocalMux I__2524 (
            .O(N__22010),
            .I(N__21999));
    Odrv4 I__2523 (
            .O(N__22007),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__2522 (
            .O(N__22002),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv12 I__2521 (
            .O(N__21999),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__2520 (
            .O(N__21992),
            .I(N__21986));
    InMux I__2519 (
            .O(N__21991),
            .I(N__21986));
    LocalMux I__2518 (
            .O(N__21986),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2517 (
            .O(N__21983),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2516 (
            .O(N__21980),
            .I(N__21974));
    InMux I__2515 (
            .O(N__21979),
            .I(N__21971));
    InMux I__2514 (
            .O(N__21978),
            .I(N__21968));
    InMux I__2513 (
            .O(N__21977),
            .I(N__21965));
    LocalMux I__2512 (
            .O(N__21974),
            .I(N__21962));
    LocalMux I__2511 (
            .O(N__21971),
            .I(N__21959));
    LocalMux I__2510 (
            .O(N__21968),
            .I(N__21952));
    LocalMux I__2509 (
            .O(N__21965),
            .I(N__21952));
    Span4Mux_s3_h I__2508 (
            .O(N__21962),
            .I(N__21952));
    Odrv4 I__2507 (
            .O(N__21959),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__2506 (
            .O(N__21952),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__2505 (
            .O(N__21947),
            .I(N__21943));
    InMux I__2504 (
            .O(N__21946),
            .I(N__21940));
    LocalMux I__2503 (
            .O(N__21943),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    LocalMux I__2502 (
            .O(N__21940),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2501 (
            .O(N__21935),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2500 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__2499 (
            .O(N__21929),
            .I(N__21926));
    Odrv4 I__2498 (
            .O(N__21926),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__2497 (
            .O(N__21923),
            .I(N__21920));
    InMux I__2496 (
            .O(N__21920),
            .I(N__21915));
    InMux I__2495 (
            .O(N__21919),
            .I(N__21912));
    InMux I__2494 (
            .O(N__21918),
            .I(N__21908));
    LocalMux I__2493 (
            .O(N__21915),
            .I(N__21905));
    LocalMux I__2492 (
            .O(N__21912),
            .I(N__21902));
    InMux I__2491 (
            .O(N__21911),
            .I(N__21899));
    LocalMux I__2490 (
            .O(N__21908),
            .I(N__21896));
    Span4Mux_v I__2489 (
            .O(N__21905),
            .I(N__21893));
    Sp12to4 I__2488 (
            .O(N__21902),
            .I(N__21888));
    LocalMux I__2487 (
            .O(N__21899),
            .I(N__21888));
    Span4Mux_s3_h I__2486 (
            .O(N__21896),
            .I(N__21885));
    Odrv4 I__2485 (
            .O(N__21893),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv12 I__2484 (
            .O(N__21888),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__2483 (
            .O(N__21885),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__2482 (
            .O(N__21878),
            .I(N__21875));
    LocalMux I__2481 (
            .O(N__21875),
            .I(N__21871));
    InMux I__2480 (
            .O(N__21874),
            .I(N__21868));
    Odrv4 I__2479 (
            .O(N__21871),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    LocalMux I__2478 (
            .O(N__21868),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2477 (
            .O(N__21863),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    CascadeMux I__2476 (
            .O(N__21860),
            .I(N__21857));
    InMux I__2475 (
            .O(N__21857),
            .I(N__21852));
    InMux I__2474 (
            .O(N__21856),
            .I(N__21849));
    InMux I__2473 (
            .O(N__21855),
            .I(N__21844));
    LocalMux I__2472 (
            .O(N__21852),
            .I(N__21841));
    LocalMux I__2471 (
            .O(N__21849),
            .I(N__21838));
    InMux I__2470 (
            .O(N__21848),
            .I(N__21835));
    InMux I__2469 (
            .O(N__21847),
            .I(N__21832));
    LocalMux I__2468 (
            .O(N__21844),
            .I(N__21829));
    Span4Mux_v I__2467 (
            .O(N__21841),
            .I(N__21826));
    Span4Mux_v I__2466 (
            .O(N__21838),
            .I(N__21823));
    LocalMux I__2465 (
            .O(N__21835),
            .I(N__21820));
    LocalMux I__2464 (
            .O(N__21832),
            .I(N__21811));
    Span4Mux_v I__2463 (
            .O(N__21829),
            .I(N__21811));
    Span4Mux_h I__2462 (
            .O(N__21826),
            .I(N__21811));
    Span4Mux_s1_h I__2461 (
            .O(N__21823),
            .I(N__21811));
    Odrv12 I__2460 (
            .O(N__21820),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__2459 (
            .O(N__21811),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__2458 (
            .O(N__21806),
            .I(N__21803));
    LocalMux I__2457 (
            .O(N__21803),
            .I(N__21800));
    Odrv4 I__2456 (
            .O(N__21800),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__2455 (
            .O(N__21797),
            .I(N__21794));
    InMux I__2454 (
            .O(N__21794),
            .I(N__21790));
    InMux I__2453 (
            .O(N__21793),
            .I(N__21786));
    LocalMux I__2452 (
            .O(N__21790),
            .I(N__21783));
    InMux I__2451 (
            .O(N__21789),
            .I(N__21780));
    LocalMux I__2450 (
            .O(N__21786),
            .I(N__21777));
    Span4Mux_v I__2449 (
            .O(N__21783),
            .I(N__21774));
    LocalMux I__2448 (
            .O(N__21780),
            .I(N__21771));
    Odrv12 I__2447 (
            .O(N__21777),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__2446 (
            .O(N__21774),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv12 I__2445 (
            .O(N__21771),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__2444 (
            .O(N__21764),
            .I(N__21761));
    LocalMux I__2443 (
            .O(N__21761),
            .I(N__21758));
    Span4Mux_h I__2442 (
            .O(N__21758),
            .I(N__21755));
    Span4Mux_v I__2441 (
            .O(N__21755),
            .I(N__21752));
    Odrv4 I__2440 (
            .O(N__21752),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2439 (
            .O(N__21749),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2438 (
            .O(N__21746),
            .I(N__21743));
    LocalMux I__2437 (
            .O(N__21743),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__2436 (
            .O(N__21740),
            .I(N__21736));
    InMux I__2435 (
            .O(N__21739),
            .I(N__21732));
    InMux I__2434 (
            .O(N__21736),
            .I(N__21729));
    InMux I__2433 (
            .O(N__21735),
            .I(N__21726));
    LocalMux I__2432 (
            .O(N__21732),
            .I(N__21721));
    LocalMux I__2431 (
            .O(N__21729),
            .I(N__21721));
    LocalMux I__2430 (
            .O(N__21726),
            .I(N__21717));
    Span4Mux_h I__2429 (
            .O(N__21721),
            .I(N__21714));
    CascadeMux I__2428 (
            .O(N__21720),
            .I(N__21711));
    Span4Mux_v I__2427 (
            .O(N__21717),
            .I(N__21708));
    Span4Mux_v I__2426 (
            .O(N__21714),
            .I(N__21705));
    InMux I__2425 (
            .O(N__21711),
            .I(N__21702));
    Odrv4 I__2424 (
            .O(N__21708),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__2423 (
            .O(N__21705),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__2422 (
            .O(N__21702),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__2421 (
            .O(N__21695),
            .I(N__21692));
    LocalMux I__2420 (
            .O(N__21692),
            .I(N__21687));
    InMux I__2419 (
            .O(N__21691),
            .I(N__21684));
    InMux I__2418 (
            .O(N__21690),
            .I(N__21681));
    Span4Mux_v I__2417 (
            .O(N__21687),
            .I(N__21674));
    LocalMux I__2416 (
            .O(N__21684),
            .I(N__21674));
    LocalMux I__2415 (
            .O(N__21681),
            .I(N__21674));
    Span4Mux_v I__2414 (
            .O(N__21674),
            .I(N__21671));
    Odrv4 I__2413 (
            .O(N__21671),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2412 (
            .O(N__21668),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__2411 (
            .O(N__21665),
            .I(N__21662));
    LocalMux I__2410 (
            .O(N__21662),
            .I(N__21659));
    Odrv4 I__2409 (
            .O(N__21659),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__2408 (
            .O(N__21656),
            .I(N__21651));
    CascadeMux I__2407 (
            .O(N__21655),
            .I(N__21648));
    InMux I__2406 (
            .O(N__21654),
            .I(N__21645));
    InMux I__2405 (
            .O(N__21651),
            .I(N__21642));
    InMux I__2404 (
            .O(N__21648),
            .I(N__21639));
    LocalMux I__2403 (
            .O(N__21645),
            .I(N__21633));
    LocalMux I__2402 (
            .O(N__21642),
            .I(N__21633));
    LocalMux I__2401 (
            .O(N__21639),
            .I(N__21630));
    InMux I__2400 (
            .O(N__21638),
            .I(N__21627));
    Span4Mux_v I__2399 (
            .O(N__21633),
            .I(N__21624));
    Span4Mux_v I__2398 (
            .O(N__21630),
            .I(N__21621));
    LocalMux I__2397 (
            .O(N__21627),
            .I(N__21618));
    Odrv4 I__2396 (
            .O(N__21624),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__2395 (
            .O(N__21621),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv12 I__2394 (
            .O(N__21618),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__2393 (
            .O(N__21611),
            .I(N__21608));
    LocalMux I__2392 (
            .O(N__21608),
            .I(N__21602));
    InMux I__2391 (
            .O(N__21607),
            .I(N__21599));
    InMux I__2390 (
            .O(N__21606),
            .I(N__21594));
    InMux I__2389 (
            .O(N__21605),
            .I(N__21594));
    Span4Mux_v I__2388 (
            .O(N__21602),
            .I(N__21587));
    LocalMux I__2387 (
            .O(N__21599),
            .I(N__21587));
    LocalMux I__2386 (
            .O(N__21594),
            .I(N__21587));
    Span4Mux_v I__2385 (
            .O(N__21587),
            .I(N__21584));
    Odrv4 I__2384 (
            .O(N__21584),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2383 (
            .O(N__21581),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__2382 (
            .O(N__21578),
            .I(N__21573));
    InMux I__2381 (
            .O(N__21577),
            .I(N__21569));
    InMux I__2380 (
            .O(N__21576),
            .I(N__21566));
    LocalMux I__2379 (
            .O(N__21573),
            .I(N__21563));
    InMux I__2378 (
            .O(N__21572),
            .I(N__21560));
    LocalMux I__2377 (
            .O(N__21569),
            .I(N__21557));
    LocalMux I__2376 (
            .O(N__21566),
            .I(N__21554));
    Span4Mux_v I__2375 (
            .O(N__21563),
            .I(N__21551));
    LocalMux I__2374 (
            .O(N__21560),
            .I(N__21544));
    Span4Mux_h I__2373 (
            .O(N__21557),
            .I(N__21544));
    Span4Mux_s3_h I__2372 (
            .O(N__21554),
            .I(N__21544));
    Odrv4 I__2371 (
            .O(N__21551),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__2370 (
            .O(N__21544),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    CascadeMux I__2369 (
            .O(N__21539),
            .I(N__21536));
    InMux I__2368 (
            .O(N__21536),
            .I(N__21533));
    LocalMux I__2367 (
            .O(N__21533),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__2366 (
            .O(N__21530),
            .I(N__21527));
    InMux I__2365 (
            .O(N__21527),
            .I(N__21524));
    LocalMux I__2364 (
            .O(N__21524),
            .I(N__21519));
    InMux I__2363 (
            .O(N__21523),
            .I(N__21516));
    InMux I__2362 (
            .O(N__21522),
            .I(N__21513));
    Span4Mux_v I__2361 (
            .O(N__21519),
            .I(N__21506));
    LocalMux I__2360 (
            .O(N__21516),
            .I(N__21506));
    LocalMux I__2359 (
            .O(N__21513),
            .I(N__21506));
    Span4Mux_v I__2358 (
            .O(N__21506),
            .I(N__21503));
    Odrv4 I__2357 (
            .O(N__21503),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2356 (
            .O(N__21500),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__2355 (
            .O(N__21497),
            .I(N__21494));
    LocalMux I__2354 (
            .O(N__21494),
            .I(N__21491));
    Odrv4 I__2353 (
            .O(N__21491),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__2352 (
            .O(N__21488),
            .I(N__21483));
    InMux I__2351 (
            .O(N__21487),
            .I(N__21480));
    InMux I__2350 (
            .O(N__21486),
            .I(N__21476));
    InMux I__2349 (
            .O(N__21483),
            .I(N__21473));
    LocalMux I__2348 (
            .O(N__21480),
            .I(N__21470));
    InMux I__2347 (
            .O(N__21479),
            .I(N__21467));
    LocalMux I__2346 (
            .O(N__21476),
            .I(N__21464));
    LocalMux I__2345 (
            .O(N__21473),
            .I(N__21461));
    Span4Mux_h I__2344 (
            .O(N__21470),
            .I(N__21454));
    LocalMux I__2343 (
            .O(N__21467),
            .I(N__21454));
    Span4Mux_h I__2342 (
            .O(N__21464),
            .I(N__21454));
    Odrv4 I__2341 (
            .O(N__21461),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__2340 (
            .O(N__21454),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__2339 (
            .O(N__21449),
            .I(N__21446));
    InMux I__2338 (
            .O(N__21446),
            .I(N__21443));
    LocalMux I__2337 (
            .O(N__21443),
            .I(N__21438));
    InMux I__2336 (
            .O(N__21442),
            .I(N__21435));
    InMux I__2335 (
            .O(N__21441),
            .I(N__21432));
    Span4Mux_v I__2334 (
            .O(N__21438),
            .I(N__21425));
    LocalMux I__2333 (
            .O(N__21435),
            .I(N__21425));
    LocalMux I__2332 (
            .O(N__21432),
            .I(N__21425));
    Span4Mux_v I__2331 (
            .O(N__21425),
            .I(N__21422));
    Odrv4 I__2330 (
            .O(N__21422),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2329 (
            .O(N__21419),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    CascadeMux I__2328 (
            .O(N__21416),
            .I(N__21413));
    InMux I__2327 (
            .O(N__21413),
            .I(N__21410));
    LocalMux I__2326 (
            .O(N__21410),
            .I(N__21407));
    Span4Mux_h I__2325 (
            .O(N__21407),
            .I(N__21404));
    Odrv4 I__2324 (
            .O(N__21404),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    CascadeMux I__2323 (
            .O(N__21401),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_ ));
    InMux I__2322 (
            .O(N__21398),
            .I(N__21394));
    InMux I__2321 (
            .O(N__21397),
            .I(N__21390));
    LocalMux I__2320 (
            .O(N__21394),
            .I(N__21387));
    InMux I__2319 (
            .O(N__21393),
            .I(N__21384));
    LocalMux I__2318 (
            .O(N__21390),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    Odrv4 I__2317 (
            .O(N__21387),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    LocalMux I__2316 (
            .O(N__21384),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    CascadeMux I__2315 (
            .O(N__21377),
            .I(N__21374));
    InMux I__2314 (
            .O(N__21374),
            .I(N__21371));
    LocalMux I__2313 (
            .O(N__21371),
            .I(N__21368));
    Span4Mux_h I__2312 (
            .O(N__21368),
            .I(N__21365));
    Odrv4 I__2311 (
            .O(N__21365),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    InMux I__2310 (
            .O(N__21362),
            .I(N__21359));
    LocalMux I__2309 (
            .O(N__21359),
            .I(\pwm_generator_inst.un19_threshold_axb_3 ));
    InMux I__2308 (
            .O(N__21356),
            .I(N__21353));
    LocalMux I__2307 (
            .O(N__21353),
            .I(N__21350));
    Odrv4 I__2306 (
            .O(N__21350),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__2305 (
            .O(N__21347),
            .I(N__21344));
    LocalMux I__2304 (
            .O(N__21344),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ));
    InMux I__2303 (
            .O(N__21341),
            .I(N__21338));
    LocalMux I__2302 (
            .O(N__21338),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    InMux I__2301 (
            .O(N__21335),
            .I(N__21329));
    InMux I__2300 (
            .O(N__21334),
            .I(N__21329));
    LocalMux I__2299 (
            .O(N__21329),
            .I(N__21325));
    InMux I__2298 (
            .O(N__21328),
            .I(N__21322));
    Span4Mux_v I__2297 (
            .O(N__21325),
            .I(N__21319));
    LocalMux I__2296 (
            .O(N__21322),
            .I(N__21316));
    Odrv4 I__2295 (
            .O(N__21319),
            .I(pwm_duty_input_9));
    Odrv4 I__2294 (
            .O(N__21316),
            .I(pwm_duty_input_9));
    CascadeMux I__2293 (
            .O(N__21311),
            .I(N__21307));
    InMux I__2292 (
            .O(N__21310),
            .I(N__21301));
    InMux I__2291 (
            .O(N__21307),
            .I(N__21301));
    InMux I__2290 (
            .O(N__21306),
            .I(N__21298));
    LocalMux I__2289 (
            .O(N__21301),
            .I(N__21295));
    LocalMux I__2288 (
            .O(N__21298),
            .I(N__21292));
    Span4Mux_h I__2287 (
            .O(N__21295),
            .I(N__21289));
    Span4Mux_s1_h I__2286 (
            .O(N__21292),
            .I(N__21286));
    Odrv4 I__2285 (
            .O(N__21289),
            .I(pwm_duty_input_8));
    Odrv4 I__2284 (
            .O(N__21286),
            .I(pwm_duty_input_8));
    CascadeMux I__2283 (
            .O(N__21281),
            .I(N__21278));
    InMux I__2282 (
            .O(N__21278),
            .I(N__21271));
    InMux I__2281 (
            .O(N__21277),
            .I(N__21271));
    InMux I__2280 (
            .O(N__21276),
            .I(N__21268));
    LocalMux I__2279 (
            .O(N__21271),
            .I(N__21265));
    LocalMux I__2278 (
            .O(N__21268),
            .I(N__21262));
    Span4Mux_h I__2277 (
            .O(N__21265),
            .I(N__21259));
    Span4Mux_v I__2276 (
            .O(N__21262),
            .I(N__21256));
    Odrv4 I__2275 (
            .O(N__21259),
            .I(pwm_duty_input_6));
    Odrv4 I__2274 (
            .O(N__21256),
            .I(pwm_duty_input_6));
    InMux I__2273 (
            .O(N__21251),
            .I(N__21247));
    InMux I__2272 (
            .O(N__21250),
            .I(N__21244));
    LocalMux I__2271 (
            .O(N__21247),
            .I(N__21241));
    LocalMux I__2270 (
            .O(N__21244),
            .I(N__21237));
    Span4Mux_v I__2269 (
            .O(N__21241),
            .I(N__21234));
    InMux I__2268 (
            .O(N__21240),
            .I(N__21231));
    Span4Mux_s1_h I__2267 (
            .O(N__21237),
            .I(N__21228));
    Odrv4 I__2266 (
            .O(N__21234),
            .I(pwm_duty_input_7));
    LocalMux I__2265 (
            .O(N__21231),
            .I(pwm_duty_input_7));
    Odrv4 I__2264 (
            .O(N__21228),
            .I(pwm_duty_input_7));
    InMux I__2263 (
            .O(N__21221),
            .I(N__21218));
    LocalMux I__2262 (
            .O(N__21218),
            .I(N__21215));
    Odrv4 I__2261 (
            .O(N__21215),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    InMux I__2260 (
            .O(N__21212),
            .I(N__21207));
    InMux I__2259 (
            .O(N__21211),
            .I(N__21204));
    InMux I__2258 (
            .O(N__21210),
            .I(N__21201));
    LocalMux I__2257 (
            .O(N__21207),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    LocalMux I__2256 (
            .O(N__21204),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    LocalMux I__2255 (
            .O(N__21201),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    InMux I__2254 (
            .O(N__21194),
            .I(N__21191));
    LocalMux I__2253 (
            .O(N__21191),
            .I(N__21188));
    Odrv4 I__2252 (
            .O(N__21188),
            .I(\pwm_generator_inst.un19_threshold_axb_2 ));
    CascadeMux I__2251 (
            .O(N__21185),
            .I(N__21182));
    InMux I__2250 (
            .O(N__21182),
            .I(N__21179));
    LocalMux I__2249 (
            .O(N__21179),
            .I(N__21176));
    Odrv4 I__2248 (
            .O(N__21176),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    CascadeMux I__2247 (
            .O(N__21173),
            .I(N__21170));
    InMux I__2246 (
            .O(N__21170),
            .I(N__21167));
    LocalMux I__2245 (
            .O(N__21167),
            .I(N__21164));
    Span4Mux_v I__2244 (
            .O(N__21164),
            .I(N__21161));
    Odrv4 I__2243 (
            .O(N__21161),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__2242 (
            .O(N__21158),
            .I(\pwm_generator_inst.un19_threshold_cry_1 ));
    InMux I__2241 (
            .O(N__21155),
            .I(\pwm_generator_inst.un19_threshold_cry_2 ));
    InMux I__2240 (
            .O(N__21152),
            .I(N__21149));
    LocalMux I__2239 (
            .O(N__21149),
            .I(\pwm_generator_inst.un19_threshold_axb_4 ));
    InMux I__2238 (
            .O(N__21146),
            .I(\pwm_generator_inst.un19_threshold_cry_3 ));
    InMux I__2237 (
            .O(N__21143),
            .I(N__21140));
    LocalMux I__2236 (
            .O(N__21140),
            .I(\pwm_generator_inst.un19_threshold_axb_5 ));
    InMux I__2235 (
            .O(N__21137),
            .I(\pwm_generator_inst.un19_threshold_cry_4 ));
    InMux I__2234 (
            .O(N__21134),
            .I(N__21131));
    LocalMux I__2233 (
            .O(N__21131),
            .I(\pwm_generator_inst.un19_threshold_axb_6 ));
    InMux I__2232 (
            .O(N__21128),
            .I(\pwm_generator_inst.un19_threshold_cry_5 ));
    InMux I__2231 (
            .O(N__21125),
            .I(N__21122));
    LocalMux I__2230 (
            .O(N__21122),
            .I(\pwm_generator_inst.un19_threshold_axb_7 ));
    InMux I__2229 (
            .O(N__21119),
            .I(\pwm_generator_inst.un19_threshold_cry_6 ));
    InMux I__2228 (
            .O(N__21116),
            .I(N__21113));
    LocalMux I__2227 (
            .O(N__21113),
            .I(\pwm_generator_inst.un19_threshold_axb_8 ));
    InMux I__2226 (
            .O(N__21110),
            .I(bfn_3_24_0_));
    InMux I__2225 (
            .O(N__21107),
            .I(N__21104));
    LocalMux I__2224 (
            .O(N__21104),
            .I(N__21101));
    Span4Mux_v I__2223 (
            .O(N__21101),
            .I(N__21098));
    Odrv4 I__2222 (
            .O(N__21098),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    InMux I__2221 (
            .O(N__21095),
            .I(\pwm_generator_inst.un19_threshold_cry_8 ));
    CascadeMux I__2220 (
            .O(N__21092),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ));
    InMux I__2219 (
            .O(N__21089),
            .I(N__21086));
    LocalMux I__2218 (
            .O(N__21086),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__2217 (
            .O(N__21083),
            .I(N__21080));
    LocalMux I__2216 (
            .O(N__21080),
            .I(N__21077));
    Odrv4 I__2215 (
            .O(N__21077),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ));
    CascadeMux I__2214 (
            .O(N__21074),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ));
    InMux I__2213 (
            .O(N__21071),
            .I(N__21068));
    LocalMux I__2212 (
            .O(N__21068),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__2211 (
            .O(N__21065),
            .I(N__21056));
    InMux I__2210 (
            .O(N__21064),
            .I(N__21051));
    InMux I__2209 (
            .O(N__21063),
            .I(N__21051));
    InMux I__2208 (
            .O(N__21062),
            .I(N__21044));
    InMux I__2207 (
            .O(N__21061),
            .I(N__21044));
    InMux I__2206 (
            .O(N__21060),
            .I(N__21044));
    InMux I__2205 (
            .O(N__21059),
            .I(N__21041));
    LocalMux I__2204 (
            .O(N__21056),
            .I(N__21036));
    LocalMux I__2203 (
            .O(N__21051),
            .I(N__21036));
    LocalMux I__2202 (
            .O(N__21044),
            .I(N__21033));
    LocalMux I__2201 (
            .O(N__21041),
            .I(N__21030));
    Span4Mux_v I__2200 (
            .O(N__21036),
            .I(N__21027));
    Span4Mux_s3_h I__2199 (
            .O(N__21033),
            .I(N__21024));
    Span4Mux_s3_h I__2198 (
            .O(N__21030),
            .I(N__21021));
    Odrv4 I__2197 (
            .O(N__21027),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    Odrv4 I__2196 (
            .O(N__21024),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    Odrv4 I__2195 (
            .O(N__21021),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    InMux I__2194 (
            .O(N__21014),
            .I(N__21011));
    LocalMux I__2193 (
            .O(N__21011),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    CascadeMux I__2192 (
            .O(N__21008),
            .I(N__21005));
    InMux I__2191 (
            .O(N__21005),
            .I(N__21002));
    LocalMux I__2190 (
            .O(N__21002),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__2189 (
            .O(N__20999),
            .I(N__20996));
    LocalMux I__2188 (
            .O(N__20996),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    InMux I__2187 (
            .O(N__20993),
            .I(N__20990));
    LocalMux I__2186 (
            .O(N__20990),
            .I(N__20987));
    Span4Mux_v I__2185 (
            .O(N__20987),
            .I(N__20984));
    Odrv4 I__2184 (
            .O(N__20984),
            .I(\pwm_generator_inst.un19_threshold_axb_1 ));
    InMux I__2183 (
            .O(N__20981),
            .I(\pwm_generator_inst.un19_threshold_cry_0 ));
    CascadeMux I__2182 (
            .O(N__20978),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ));
    InMux I__2181 (
            .O(N__20975),
            .I(N__20972));
    LocalMux I__2180 (
            .O(N__20972),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ));
    InMux I__2179 (
            .O(N__20969),
            .I(N__20966));
    LocalMux I__2178 (
            .O(N__20966),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ));
    CascadeMux I__2177 (
            .O(N__20963),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ));
    InMux I__2176 (
            .O(N__20960),
            .I(N__20957));
    LocalMux I__2175 (
            .O(N__20957),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    InMux I__2174 (
            .O(N__20954),
            .I(N__20951));
    LocalMux I__2173 (
            .O(N__20951),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__2172 (
            .O(N__20948),
            .I(N__20945));
    LocalMux I__2171 (
            .O(N__20945),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__2170 (
            .O(N__20942),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ));
    InMux I__2169 (
            .O(N__20939),
            .I(N__20936));
    LocalMux I__2168 (
            .O(N__20936),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ));
    CascadeMux I__2167 (
            .O(N__20933),
            .I(N__20930));
    InMux I__2166 (
            .O(N__20930),
            .I(N__20927));
    LocalMux I__2165 (
            .O(N__20927),
            .I(N__20924));
    Odrv4 I__2164 (
            .O(N__20924),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    CascadeMux I__2163 (
            .O(N__20921),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    CascadeMux I__2162 (
            .O(N__20918),
            .I(\current_shift_inst.PI_CTRL.N_44_cascade_ ));
    InMux I__2161 (
            .O(N__20915),
            .I(N__20912));
    LocalMux I__2160 (
            .O(N__20912),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ));
    CascadeMux I__2159 (
            .O(N__20909),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_ ));
    InMux I__2158 (
            .O(N__20906),
            .I(N__20903));
    LocalMux I__2157 (
            .O(N__20903),
            .I(N__20900));
    Odrv4 I__2156 (
            .O(N__20900),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    InMux I__2155 (
            .O(N__20897),
            .I(N__20894));
    LocalMux I__2154 (
            .O(N__20894),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    InMux I__2153 (
            .O(N__20891),
            .I(N__20888));
    LocalMux I__2152 (
            .O(N__20888),
            .I(\current_shift_inst.PI_CTRL.N_77 ));
    InMux I__2151 (
            .O(N__20885),
            .I(N__20881));
    InMux I__2150 (
            .O(N__20884),
            .I(N__20877));
    LocalMux I__2149 (
            .O(N__20881),
            .I(N__20874));
    InMux I__2148 (
            .O(N__20880),
            .I(N__20871));
    LocalMux I__2147 (
            .O(N__20877),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv12 I__2146 (
            .O(N__20874),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    LocalMux I__2145 (
            .O(N__20871),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__2144 (
            .O(N__20864),
            .I(N__20861));
    LocalMux I__2143 (
            .O(N__20861),
            .I(N__20858));
    Span4Mux_s1_v I__2142 (
            .O(N__20858),
            .I(N__20855));
    Odrv4 I__2141 (
            .O(N__20855),
            .I(rgb_drv_RNOZ0));
    CascadeMux I__2140 (
            .O(N__20852),
            .I(N__20849));
    InMux I__2139 (
            .O(N__20849),
            .I(N__20846));
    LocalMux I__2138 (
            .O(N__20846),
            .I(N__20843));
    Span4Mux_h I__2137 (
            .O(N__20843),
            .I(N__20840));
    Odrv4 I__2136 (
            .O(N__20840),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__2135 (
            .O(N__20837),
            .I(N__20834));
    LocalMux I__2134 (
            .O(N__20834),
            .I(N__20831));
    Odrv4 I__2133 (
            .O(N__20831),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    CascadeMux I__2132 (
            .O(N__20828),
            .I(N__20825));
    InMux I__2131 (
            .O(N__20825),
            .I(N__20822));
    LocalMux I__2130 (
            .O(N__20822),
            .I(N__20819));
    Span4Mux_h I__2129 (
            .O(N__20819),
            .I(N__20816));
    Odrv4 I__2128 (
            .O(N__20816),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    CascadeMux I__2127 (
            .O(N__20813),
            .I(N__20810));
    InMux I__2126 (
            .O(N__20810),
            .I(N__20807));
    LocalMux I__2125 (
            .O(N__20807),
            .I(N__20804));
    Span4Mux_v I__2124 (
            .O(N__20804),
            .I(N__20801));
    Odrv4 I__2123 (
            .O(N__20801),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__2122 (
            .O(N__20798),
            .I(N__20794));
    CascadeMux I__2121 (
            .O(N__20797),
            .I(N__20791));
    LocalMux I__2120 (
            .O(N__20794),
            .I(N__20788));
    InMux I__2119 (
            .O(N__20791),
            .I(N__20785));
    Span4Mux_h I__2118 (
            .O(N__20788),
            .I(N__20780));
    LocalMux I__2117 (
            .O(N__20785),
            .I(N__20780));
    Span4Mux_v I__2116 (
            .O(N__20780),
            .I(N__20777));
    Odrv4 I__2115 (
            .O(N__20777),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    CascadeMux I__2114 (
            .O(N__20774),
            .I(N__20771));
    InMux I__2113 (
            .O(N__20771),
            .I(N__20768));
    LocalMux I__2112 (
            .O(N__20768),
            .I(N__20765));
    Span4Mux_h I__2111 (
            .O(N__20765),
            .I(N__20762));
    Odrv4 I__2110 (
            .O(N__20762),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__2109 (
            .O(N__20759),
            .I(N__20756));
    LocalMux I__2108 (
            .O(N__20756),
            .I(N__20753));
    Span4Mux_v I__2107 (
            .O(N__20753),
            .I(N__20750));
    Odrv4 I__2106 (
            .O(N__20750),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__2105 (
            .O(N__20747),
            .I(N__20744));
    LocalMux I__2104 (
            .O(N__20744),
            .I(N__20741));
    Odrv4 I__2103 (
            .O(N__20741),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    InMux I__2102 (
            .O(N__20738),
            .I(N__20735));
    LocalMux I__2101 (
            .O(N__20735),
            .I(N__20732));
    Odrv4 I__2100 (
            .O(N__20732),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__2099 (
            .O(N__20729),
            .I(N__20726));
    LocalMux I__2098 (
            .O(N__20726),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__2097 (
            .O(N__20723),
            .I(N__20718));
    InMux I__2096 (
            .O(N__20722),
            .I(N__20715));
    InMux I__2095 (
            .O(N__20721),
            .I(N__20712));
    LocalMux I__2094 (
            .O(N__20718),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__2093 (
            .O(N__20715),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__2092 (
            .O(N__20712),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    CascadeMux I__2091 (
            .O(N__20705),
            .I(N__20702));
    InMux I__2090 (
            .O(N__20702),
            .I(N__20698));
    InMux I__2089 (
            .O(N__20701),
            .I(N__20694));
    LocalMux I__2088 (
            .O(N__20698),
            .I(N__20691));
    InMux I__2087 (
            .O(N__20697),
            .I(N__20688));
    LocalMux I__2086 (
            .O(N__20694),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    Odrv4 I__2085 (
            .O(N__20691),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__2084 (
            .O(N__20688),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    InMux I__2083 (
            .O(N__20681),
            .I(N__20677));
    InMux I__2082 (
            .O(N__20680),
            .I(N__20673));
    LocalMux I__2081 (
            .O(N__20677),
            .I(N__20670));
    InMux I__2080 (
            .O(N__20676),
            .I(N__20667));
    LocalMux I__2079 (
            .O(N__20673),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    Odrv4 I__2078 (
            .O(N__20670),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    LocalMux I__2077 (
            .O(N__20667),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__2076 (
            .O(N__20660),
            .I(N__20657));
    LocalMux I__2075 (
            .O(N__20657),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    CascadeMux I__2074 (
            .O(N__20654),
            .I(N__20647));
    InMux I__2073 (
            .O(N__20653),
            .I(N__20640));
    InMux I__2072 (
            .O(N__20652),
            .I(N__20640));
    InMux I__2071 (
            .O(N__20651),
            .I(N__20640));
    InMux I__2070 (
            .O(N__20650),
            .I(N__20632));
    InMux I__2069 (
            .O(N__20647),
            .I(N__20632));
    LocalMux I__2068 (
            .O(N__20640),
            .I(N__20629));
    InMux I__2067 (
            .O(N__20639),
            .I(N__20622));
    InMux I__2066 (
            .O(N__20638),
            .I(N__20622));
    InMux I__2065 (
            .O(N__20637),
            .I(N__20622));
    LocalMux I__2064 (
            .O(N__20632),
            .I(N__20615));
    Span4Mux_v I__2063 (
            .O(N__20629),
            .I(N__20615));
    LocalMux I__2062 (
            .O(N__20622),
            .I(N__20615));
    Odrv4 I__2061 (
            .O(N__20615),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    CascadeMux I__2060 (
            .O(N__20612),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    CascadeMux I__2059 (
            .O(N__20609),
            .I(N__20605));
    CascadeMux I__2058 (
            .O(N__20608),
            .I(N__20602));
    InMux I__2057 (
            .O(N__20605),
            .I(N__20598));
    InMux I__2056 (
            .O(N__20602),
            .I(N__20593));
    InMux I__2055 (
            .O(N__20601),
            .I(N__20593));
    LocalMux I__2054 (
            .O(N__20598),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__2053 (
            .O(N__20593),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__2052 (
            .O(N__20588),
            .I(N__20584));
    InMux I__2051 (
            .O(N__20587),
            .I(N__20581));
    LocalMux I__2050 (
            .O(N__20584),
            .I(N__20578));
    LocalMux I__2049 (
            .O(N__20581),
            .I(pwm_duty_input_0));
    Odrv4 I__2048 (
            .O(N__20578),
            .I(pwm_duty_input_0));
    InMux I__2047 (
            .O(N__20573),
            .I(N__20570));
    LocalMux I__2046 (
            .O(N__20570),
            .I(N__20566));
    InMux I__2045 (
            .O(N__20569),
            .I(N__20563));
    Span4Mux_v I__2044 (
            .O(N__20566),
            .I(N__20560));
    LocalMux I__2043 (
            .O(N__20563),
            .I(pwm_duty_input_1));
    Odrv4 I__2042 (
            .O(N__20560),
            .I(pwm_duty_input_1));
    InMux I__2041 (
            .O(N__20555),
            .I(N__20551));
    InMux I__2040 (
            .O(N__20554),
            .I(N__20548));
    LocalMux I__2039 (
            .O(N__20551),
            .I(N__20545));
    LocalMux I__2038 (
            .O(N__20548),
            .I(N__20540));
    Span4Mux_v I__2037 (
            .O(N__20545),
            .I(N__20540));
    Odrv4 I__2036 (
            .O(N__20540),
            .I(pwm_duty_input_2));
    InMux I__2035 (
            .O(N__20537),
            .I(N__20534));
    LocalMux I__2034 (
            .O(N__20534),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    CascadeMux I__2033 (
            .O(N__20531),
            .I(N__20527));
    InMux I__2032 (
            .O(N__20530),
            .I(N__20524));
    InMux I__2031 (
            .O(N__20527),
            .I(N__20521));
    LocalMux I__2030 (
            .O(N__20524),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    LocalMux I__2029 (
            .O(N__20521),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    InMux I__2028 (
            .O(N__20516),
            .I(N__20513));
    LocalMux I__2027 (
            .O(N__20513),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    CascadeMux I__2026 (
            .O(N__20510),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15_cascade_ ));
    CascadeMux I__2025 (
            .O(N__20507),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ));
    CascadeMux I__2024 (
            .O(N__20504),
            .I(\current_shift_inst.PI_CTRL.N_43_cascade_ ));
    InMux I__2023 (
            .O(N__20501),
            .I(N__20498));
    LocalMux I__2022 (
            .O(N__20498),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__2021 (
            .O(N__20495),
            .I(N__20492));
    LocalMux I__2020 (
            .O(N__20492),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    CascadeMux I__2019 (
            .O(N__20489),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ));
    InMux I__2018 (
            .O(N__20486),
            .I(N__20483));
    LocalMux I__2017 (
            .O(N__20483),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    CascadeMux I__2016 (
            .O(N__20480),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ));
    InMux I__2015 (
            .O(N__20477),
            .I(N__20474));
    LocalMux I__2014 (
            .O(N__20474),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    InMux I__2013 (
            .O(N__20471),
            .I(N__20468));
    LocalMux I__2012 (
            .O(N__20468),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__2011 (
            .O(N__20465),
            .I(N__20462));
    LocalMux I__2010 (
            .O(N__20462),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    CascadeMux I__2009 (
            .O(N__20459),
            .I(N__20456));
    InMux I__2008 (
            .O(N__20456),
            .I(N__20453));
    LocalMux I__2007 (
            .O(N__20453),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__2006 (
            .O(N__20450),
            .I(N__20447));
    LocalMux I__2005 (
            .O(N__20447),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    CascadeMux I__2004 (
            .O(N__20444),
            .I(N__20441));
    InMux I__2003 (
            .O(N__20441),
            .I(N__20438));
    LocalMux I__2002 (
            .O(N__20438),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    CascadeMux I__2001 (
            .O(N__20435),
            .I(N__20432));
    InMux I__2000 (
            .O(N__20432),
            .I(N__20429));
    LocalMux I__1999 (
            .O(N__20429),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    CascadeMux I__1998 (
            .O(N__20426),
            .I(N__20423));
    InMux I__1997 (
            .O(N__20423),
            .I(N__20420));
    LocalMux I__1996 (
            .O(N__20420),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__1995 (
            .O(N__20417),
            .I(N__20414));
    LocalMux I__1994 (
            .O(N__20414),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__1993 (
            .O(N__20411),
            .I(N__20408));
    InMux I__1992 (
            .O(N__20408),
            .I(N__20405));
    LocalMux I__1991 (
            .O(N__20405),
            .I(N__20402));
    Odrv4 I__1990 (
            .O(N__20402),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__1989 (
            .O(N__20399),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__1988 (
            .O(N__20396),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__1987 (
            .O(N__20393),
            .I(N__20390));
    LocalMux I__1986 (
            .O(N__20390),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__1985 (
            .O(N__20387),
            .I(N__20384));
    LocalMux I__1984 (
            .O(N__20384),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    CascadeMux I__1983 (
            .O(N__20381),
            .I(N__20378));
    InMux I__1982 (
            .O(N__20378),
            .I(N__20375));
    LocalMux I__1981 (
            .O(N__20375),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    CascadeMux I__1980 (
            .O(N__20372),
            .I(N__20369));
    InMux I__1979 (
            .O(N__20369),
            .I(N__20366));
    LocalMux I__1978 (
            .O(N__20366),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__1977 (
            .O(N__20363),
            .I(N__20360));
    LocalMux I__1976 (
            .O(N__20360),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__1975 (
            .O(N__20357),
            .I(N__20354));
    LocalMux I__1974 (
            .O(N__20354),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    CascadeMux I__1973 (
            .O(N__20351),
            .I(N__20348));
    InMux I__1972 (
            .O(N__20348),
            .I(N__20345));
    LocalMux I__1971 (
            .O(N__20345),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__1970 (
            .O(N__20342),
            .I(N__20339));
    LocalMux I__1969 (
            .O(N__20339),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1968 (
            .O(N__20336),
            .I(N__20333));
    LocalMux I__1967 (
            .O(N__20333),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    InMux I__1966 (
            .O(N__20330),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    InMux I__1965 (
            .O(N__20327),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    InMux I__1964 (
            .O(N__20324),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__1963 (
            .O(N__20321),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    InMux I__1962 (
            .O(N__20318),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    InMux I__1961 (
            .O(N__20315),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    InMux I__1960 (
            .O(N__20312),
            .I(bfn_1_26_0_));
    InMux I__1959 (
            .O(N__20309),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__1958 (
            .O(N__20306),
            .I(N__20303));
    LocalMux I__1957 (
            .O(N__20303),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1956 (
            .O(N__20300),
            .I(N__20297));
    LocalMux I__1955 (
            .O(N__20297),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__1954 (
            .O(N__20294),
            .I(N__20291));
    LocalMux I__1953 (
            .O(N__20291),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1952 (
            .O(N__20288),
            .I(N__20285));
    LocalMux I__1951 (
            .O(N__20285),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__1950 (
            .O(N__20282),
            .I(N__20279));
    LocalMux I__1949 (
            .O(N__20279),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1948 (
            .O(N__20276),
            .I(N__20273));
    LocalMux I__1947 (
            .O(N__20273),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    InMux I__1946 (
            .O(N__20270),
            .I(N__20267));
    LocalMux I__1945 (
            .O(N__20267),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1944 (
            .O(N__20264),
            .I(N__20261));
    LocalMux I__1943 (
            .O(N__20261),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    InMux I__1942 (
            .O(N__20258),
            .I(N__20255));
    LocalMux I__1941 (
            .O(N__20255),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1940 (
            .O(N__20252),
            .I(N__20249));
    LocalMux I__1939 (
            .O(N__20249),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__1938 (
            .O(N__20246),
            .I(N__20243));
    LocalMux I__1937 (
            .O(N__20243),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1936 (
            .O(N__20240),
            .I(N__20237));
    LocalMux I__1935 (
            .O(N__20237),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    InMux I__1934 (
            .O(N__20234),
            .I(N__20231));
    LocalMux I__1933 (
            .O(N__20231),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__1932 (
            .O(N__20228),
            .I(N__20225));
    LocalMux I__1931 (
            .O(N__20225),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__1930 (
            .O(N__20222),
            .I(N__20219));
    LocalMux I__1929 (
            .O(N__20219),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1928 (
            .O(N__20216),
            .I(N__20213));
    LocalMux I__1927 (
            .O(N__20213),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__1926 (
            .O(N__20210),
            .I(N__20207));
    LocalMux I__1925 (
            .O(N__20207),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    InMux I__1924 (
            .O(N__20204),
            .I(N__20200));
    InMux I__1923 (
            .O(N__20203),
            .I(N__20197));
    LocalMux I__1922 (
            .O(N__20200),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    LocalMux I__1921 (
            .O(N__20197),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    CascadeMux I__1920 (
            .O(N__20192),
            .I(N__20189));
    InMux I__1919 (
            .O(N__20189),
            .I(N__20186));
    LocalMux I__1918 (
            .O(N__20186),
            .I(N__20182));
    InMux I__1917 (
            .O(N__20185),
            .I(N__20179));
    Odrv4 I__1916 (
            .O(N__20182),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__1915 (
            .O(N__20179),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__1914 (
            .O(N__20174),
            .I(N__20171));
    LocalMux I__1913 (
            .O(N__20171),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    InMux I__1912 (
            .O(N__20168),
            .I(N__20159));
    InMux I__1911 (
            .O(N__20167),
            .I(N__20159));
    InMux I__1910 (
            .O(N__20166),
            .I(N__20159));
    LocalMux I__1909 (
            .O(N__20159),
            .I(\current_shift_inst.PI_CTRL.N_161 ));
    InMux I__1908 (
            .O(N__20156),
            .I(N__20153));
    LocalMux I__1907 (
            .O(N__20153),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1906 (
            .O(N__20150),
            .I(N__20147));
    LocalMux I__1905 (
            .O(N__20147),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    CascadeMux I__1904 (
            .O(N__20144),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ));
    CascadeMux I__1903 (
            .O(N__20141),
            .I(\current_shift_inst.PI_CTRL.N_98_cascade_ ));
    CascadeMux I__1902 (
            .O(N__20138),
            .I(\current_shift_inst.PI_CTRL.N_96_cascade_ ));
    InMux I__1901 (
            .O(N__20135),
            .I(N__20132));
    LocalMux I__1900 (
            .O(N__20132),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    InMux I__1899 (
            .O(N__20129),
            .I(N__20126));
    LocalMux I__1898 (
            .O(N__20126),
            .I(N__20123));
    Odrv12 I__1897 (
            .O(N__20123),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    CascadeMux I__1896 (
            .O(N__20120),
            .I(N__20117));
    InMux I__1895 (
            .O(N__20117),
            .I(N__20114));
    LocalMux I__1894 (
            .O(N__20114),
            .I(N__20111));
    Span4Mux_v I__1893 (
            .O(N__20111),
            .I(N__20108));
    Odrv4 I__1892 (
            .O(N__20108),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__1891 (
            .O(N__20105),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    CascadeMux I__1890 (
            .O(N__20102),
            .I(N__20099));
    InMux I__1889 (
            .O(N__20099),
            .I(N__20096));
    LocalMux I__1888 (
            .O(N__20096),
            .I(N__20093));
    Odrv12 I__1887 (
            .O(N__20093),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__1886 (
            .O(N__20090),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    CascadeMux I__1885 (
            .O(N__20087),
            .I(N__20084));
    InMux I__1884 (
            .O(N__20084),
            .I(N__20081));
    LocalMux I__1883 (
            .O(N__20081),
            .I(N__20078));
    Span4Mux_v I__1882 (
            .O(N__20078),
            .I(N__20075));
    Odrv4 I__1881 (
            .O(N__20075),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__1880 (
            .O(N__20072),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__1879 (
            .O(N__20069),
            .I(N__20066));
    LocalMux I__1878 (
            .O(N__20066),
            .I(N__20063));
    Span4Mux_v I__1877 (
            .O(N__20063),
            .I(N__20060));
    Odrv4 I__1876 (
            .O(N__20060),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    CascadeMux I__1875 (
            .O(N__20057),
            .I(N__20054));
    InMux I__1874 (
            .O(N__20054),
            .I(N__20051));
    LocalMux I__1873 (
            .O(N__20051),
            .I(N__20048));
    Odrv12 I__1872 (
            .O(N__20048),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ));
    InMux I__1871 (
            .O(N__20045),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__1870 (
            .O(N__20042),
            .I(N__20039));
    LocalMux I__1869 (
            .O(N__20039),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    CascadeMux I__1868 (
            .O(N__20036),
            .I(N__20033));
    InMux I__1867 (
            .O(N__20033),
            .I(N__20030));
    LocalMux I__1866 (
            .O(N__20030),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__1865 (
            .O(N__20027),
            .I(N__20024));
    LocalMux I__1864 (
            .O(N__20024),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__1863 (
            .O(N__20021),
            .I(N__20018));
    LocalMux I__1862 (
            .O(N__20018),
            .I(N__20015));
    Span4Mux_v I__1861 (
            .O(N__20015),
            .I(N__20012));
    Odrv4 I__1860 (
            .O(N__20012),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__1859 (
            .O(N__20009),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    InMux I__1858 (
            .O(N__20006),
            .I(N__20003));
    LocalMux I__1857 (
            .O(N__20003),
            .I(N__20000));
    Odrv12 I__1856 (
            .O(N__20000),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__1855 (
            .O(N__19997),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__1854 (
            .O(N__19994),
            .I(N__19991));
    InMux I__1853 (
            .O(N__19991),
            .I(N__19988));
    LocalMux I__1852 (
            .O(N__19988),
            .I(N__19985));
    Span4Mux_v I__1851 (
            .O(N__19985),
            .I(N__19982));
    Odrv4 I__1850 (
            .O(N__19982),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__1849 (
            .O(N__19979),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    CascadeMux I__1848 (
            .O(N__19976),
            .I(N__19973));
    InMux I__1847 (
            .O(N__19973),
            .I(N__19970));
    LocalMux I__1846 (
            .O(N__19970),
            .I(N__19967));
    Span4Mux_v I__1845 (
            .O(N__19967),
            .I(N__19964));
    Odrv4 I__1844 (
            .O(N__19964),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__1843 (
            .O(N__19961),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    CascadeMux I__1842 (
            .O(N__19958),
            .I(N__19955));
    InMux I__1841 (
            .O(N__19955),
            .I(N__19952));
    LocalMux I__1840 (
            .O(N__19952),
            .I(N__19949));
    Span4Mux_v I__1839 (
            .O(N__19949),
            .I(N__19946));
    Odrv4 I__1838 (
            .O(N__19946),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__1837 (
            .O(N__19943),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__1836 (
            .O(N__19940),
            .I(N__19937));
    InMux I__1835 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__1834 (
            .O(N__19934),
            .I(N__19931));
    Span4Mux_v I__1833 (
            .O(N__19931),
            .I(N__19928));
    Odrv4 I__1832 (
            .O(N__19928),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__1831 (
            .O(N__19925),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    CascadeMux I__1830 (
            .O(N__19922),
            .I(N__19919));
    InMux I__1829 (
            .O(N__19919),
            .I(N__19916));
    LocalMux I__1828 (
            .O(N__19916),
            .I(N__19913));
    Span4Mux_v I__1827 (
            .O(N__19913),
            .I(N__19910));
    Odrv4 I__1826 (
            .O(N__19910),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__1825 (
            .O(N__19907),
            .I(bfn_1_16_0_));
    CascadeMux I__1824 (
            .O(N__19904),
            .I(N__19901));
    InMux I__1823 (
            .O(N__19901),
            .I(N__19898));
    LocalMux I__1822 (
            .O(N__19898),
            .I(N__19895));
    Span4Mux_v I__1821 (
            .O(N__19895),
            .I(N__19892));
    Odrv4 I__1820 (
            .O(N__19892),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__1819 (
            .O(N__19889),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    CascadeMux I__1818 (
            .O(N__19886),
            .I(N__19883));
    InMux I__1817 (
            .O(N__19883),
            .I(N__19880));
    LocalMux I__1816 (
            .O(N__19880),
            .I(N__19877));
    Span4Mux_v I__1815 (
            .O(N__19877),
            .I(N__19874));
    Odrv4 I__1814 (
            .O(N__19874),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    InMux I__1813 (
            .O(N__19871),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    CascadeMux I__1812 (
            .O(N__19868),
            .I(N__19865));
    InMux I__1811 (
            .O(N__19865),
            .I(N__19862));
    LocalMux I__1810 (
            .O(N__19862),
            .I(N__19859));
    Odrv4 I__1809 (
            .O(N__19859),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    InMux I__1808 (
            .O(N__19856),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    CascadeMux I__1807 (
            .O(N__19853),
            .I(N__19850));
    InMux I__1806 (
            .O(N__19850),
            .I(N__19847));
    LocalMux I__1805 (
            .O(N__19847),
            .I(N__19844));
    Odrv4 I__1804 (
            .O(N__19844),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    InMux I__1803 (
            .O(N__19841),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__1802 (
            .O(N__19838),
            .I(N__19835));
    InMux I__1801 (
            .O(N__19835),
            .I(N__19832));
    LocalMux I__1800 (
            .O(N__19832),
            .I(N__19829));
    Span4Mux_v I__1799 (
            .O(N__19829),
            .I(N__19826));
    Odrv4 I__1798 (
            .O(N__19826),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__1797 (
            .O(N__19823),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    CascadeMux I__1796 (
            .O(N__19820),
            .I(N__19817));
    InMux I__1795 (
            .O(N__19817),
            .I(N__19814));
    LocalMux I__1794 (
            .O(N__19814),
            .I(N__19811));
    Odrv4 I__1793 (
            .O(N__19811),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__1792 (
            .O(N__19808),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__1791 (
            .O(N__19805),
            .I(N__19802));
    InMux I__1790 (
            .O(N__19802),
            .I(N__19799));
    LocalMux I__1789 (
            .O(N__19799),
            .I(N__19796));
    Span4Mux_h I__1788 (
            .O(N__19796),
            .I(N__19793));
    Odrv4 I__1787 (
            .O(N__19793),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    InMux I__1786 (
            .O(N__19790),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__1785 (
            .O(N__19787),
            .I(N__19784));
    InMux I__1784 (
            .O(N__19784),
            .I(N__19781));
    LocalMux I__1783 (
            .O(N__19781),
            .I(N__19778));
    Odrv12 I__1782 (
            .O(N__19778),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    InMux I__1781 (
            .O(N__19775),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    CascadeMux I__1780 (
            .O(N__19772),
            .I(N__19769));
    InMux I__1779 (
            .O(N__19769),
            .I(N__19766));
    LocalMux I__1778 (
            .O(N__19766),
            .I(N__19763));
    Span4Mux_v I__1777 (
            .O(N__19763),
            .I(N__19760));
    Odrv4 I__1776 (
            .O(N__19760),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    InMux I__1775 (
            .O(N__19757),
            .I(bfn_1_15_0_));
    CascadeMux I__1774 (
            .O(N__19754),
            .I(N__19751));
    InMux I__1773 (
            .O(N__19751),
            .I(N__19748));
    LocalMux I__1772 (
            .O(N__19748),
            .I(N__19745));
    Span4Mux_v I__1771 (
            .O(N__19745),
            .I(N__19742));
    Odrv4 I__1770 (
            .O(N__19742),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__1769 (
            .O(N__19739),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__1768 (
            .O(N__19736),
            .I(N__19733));
    InMux I__1767 (
            .O(N__19733),
            .I(N__19730));
    LocalMux I__1766 (
            .O(N__19730),
            .I(N__19727));
    Span4Mux_v I__1765 (
            .O(N__19727),
            .I(N__19724));
    Odrv4 I__1764 (
            .O(N__19724),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__1763 (
            .O(N__19721),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    InMux I__1762 (
            .O(N__19718),
            .I(N__19715));
    LocalMux I__1761 (
            .O(N__19715),
            .I(N__19712));
    Odrv4 I__1760 (
            .O(N__19712),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__1759 (
            .O(N__19709),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CascadeMux I__1758 (
            .O(N__19706),
            .I(N__19703));
    InMux I__1757 (
            .O(N__19703),
            .I(N__19700));
    LocalMux I__1756 (
            .O(N__19700),
            .I(N__19697));
    Odrv4 I__1755 (
            .O(N__19697),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    InMux I__1754 (
            .O(N__19694),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    CascadeMux I__1753 (
            .O(N__19691),
            .I(N__19688));
    InMux I__1752 (
            .O(N__19688),
            .I(N__19685));
    LocalMux I__1751 (
            .O(N__19685),
            .I(N__19682));
    Span4Mux_h I__1750 (
            .O(N__19682),
            .I(N__19679));
    Odrv4 I__1749 (
            .O(N__19679),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    InMux I__1748 (
            .O(N__19676),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__1747 (
            .O(N__19673),
            .I(N__19670));
    InMux I__1746 (
            .O(N__19670),
            .I(N__19667));
    LocalMux I__1745 (
            .O(N__19667),
            .I(N__19664));
    Odrv4 I__1744 (
            .O(N__19664),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__1743 (
            .O(N__19661),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__1742 (
            .O(N__19658),
            .I(N__19655));
    InMux I__1741 (
            .O(N__19655),
            .I(N__19652));
    LocalMux I__1740 (
            .O(N__19652),
            .I(N__19649));
    Span4Mux_v I__1739 (
            .O(N__19649),
            .I(N__19646));
    Odrv4 I__1738 (
            .O(N__19646),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__1737 (
            .O(N__19643),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__1736 (
            .O(N__19640),
            .I(N__19637));
    InMux I__1735 (
            .O(N__19637),
            .I(N__19634));
    LocalMux I__1734 (
            .O(N__19634),
            .I(N__19631));
    Span4Mux_v I__1733 (
            .O(N__19631),
            .I(N__19628));
    Odrv4 I__1732 (
            .O(N__19628),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__1731 (
            .O(N__19625),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    CascadeMux I__1730 (
            .O(N__19622),
            .I(N__19619));
    InMux I__1729 (
            .O(N__19619),
            .I(N__19616));
    LocalMux I__1728 (
            .O(N__19616),
            .I(N__19613));
    Span4Mux_v I__1727 (
            .O(N__19613),
            .I(N__19610));
    Odrv4 I__1726 (
            .O(N__19610),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    InMux I__1725 (
            .O(N__19607),
            .I(bfn_1_14_0_));
    CascadeMux I__1724 (
            .O(N__19604),
            .I(N__19601));
    InMux I__1723 (
            .O(N__19601),
            .I(N__19598));
    LocalMux I__1722 (
            .O(N__19598),
            .I(N__19595));
    Span4Mux_v I__1721 (
            .O(N__19595),
            .I(N__19592));
    Odrv4 I__1720 (
            .O(N__19592),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__1719 (
            .O(N__19589),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    InMux I__1718 (
            .O(N__19586),
            .I(N__19583));
    LocalMux I__1717 (
            .O(N__19583),
            .I(N__19580));
    Span4Mux_v I__1716 (
            .O(N__19580),
            .I(N__19577));
    Odrv4 I__1715 (
            .O(N__19577),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    InMux I__1714 (
            .O(N__19574),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    InMux I__1713 (
            .O(N__19571),
            .I(N__19568));
    LocalMux I__1712 (
            .O(N__19568),
            .I(N__19565));
    Span4Mux_v I__1711 (
            .O(N__19565),
            .I(N__19562));
    Odrv4 I__1710 (
            .O(N__19562),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    InMux I__1709 (
            .O(N__19559),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__1708 (
            .O(N__19556),
            .I(N__19553));
    LocalMux I__1707 (
            .O(N__19553),
            .I(N__19550));
    Span4Mux_v I__1706 (
            .O(N__19550),
            .I(N__19547));
    Odrv4 I__1705 (
            .O(N__19547),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    InMux I__1704 (
            .O(N__19544),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    InMux I__1703 (
            .O(N__19541),
            .I(N__19538));
    LocalMux I__1702 (
            .O(N__19538),
            .I(N__19535));
    Span4Mux_h I__1701 (
            .O(N__19535),
            .I(N__19532));
    Span4Mux_v I__1700 (
            .O(N__19532),
            .I(N__19529));
    Odrv4 I__1699 (
            .O(N__19529),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    InMux I__1698 (
            .O(N__19526),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__1697 (
            .O(N__19523),
            .I(N__19520));
    LocalMux I__1696 (
            .O(N__19520),
            .I(N__19517));
    Span4Mux_v I__1695 (
            .O(N__19517),
            .I(N__19514));
    Span4Mux_s1_h I__1694 (
            .O(N__19514),
            .I(N__19511));
    Odrv4 I__1693 (
            .O(N__19511),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    InMux I__1692 (
            .O(N__19508),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    InMux I__1691 (
            .O(N__19505),
            .I(N__19502));
    LocalMux I__1690 (
            .O(N__19502),
            .I(N__19499));
    Span4Mux_v I__1689 (
            .O(N__19499),
            .I(N__19496));
    Odrv4 I__1688 (
            .O(N__19496),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    InMux I__1687 (
            .O(N__19493),
            .I(N__19479));
    CascadeMux I__1686 (
            .O(N__19492),
            .I(N__19476));
    CascadeMux I__1685 (
            .O(N__19491),
            .I(N__19473));
    CascadeMux I__1684 (
            .O(N__19490),
            .I(N__19470));
    CascadeMux I__1683 (
            .O(N__19489),
            .I(N__19467));
    CascadeMux I__1682 (
            .O(N__19488),
            .I(N__19464));
    CascadeMux I__1681 (
            .O(N__19487),
            .I(N__19461));
    CascadeMux I__1680 (
            .O(N__19486),
            .I(N__19458));
    CascadeMux I__1679 (
            .O(N__19485),
            .I(N__19455));
    CascadeMux I__1678 (
            .O(N__19484),
            .I(N__19452));
    CascadeMux I__1677 (
            .O(N__19483),
            .I(N__19449));
    CascadeMux I__1676 (
            .O(N__19482),
            .I(N__19446));
    LocalMux I__1675 (
            .O(N__19479),
            .I(N__19443));
    InMux I__1674 (
            .O(N__19476),
            .I(N__19436));
    InMux I__1673 (
            .O(N__19473),
            .I(N__19436));
    InMux I__1672 (
            .O(N__19470),
            .I(N__19436));
    InMux I__1671 (
            .O(N__19467),
            .I(N__19427));
    InMux I__1670 (
            .O(N__19464),
            .I(N__19427));
    InMux I__1669 (
            .O(N__19461),
            .I(N__19427));
    InMux I__1668 (
            .O(N__19458),
            .I(N__19427));
    InMux I__1667 (
            .O(N__19455),
            .I(N__19422));
    InMux I__1666 (
            .O(N__19452),
            .I(N__19422));
    InMux I__1665 (
            .O(N__19449),
            .I(N__19417));
    InMux I__1664 (
            .O(N__19446),
            .I(N__19417));
    Odrv4 I__1663 (
            .O(N__19443),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1662 (
            .O(N__19436),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1661 (
            .O(N__19427),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1660 (
            .O(N__19422),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1659 (
            .O(N__19417),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    InMux I__1658 (
            .O(N__19406),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__1657 (
            .O(N__19403),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    InMux I__1656 (
            .O(N__19400),
            .I(N__19397));
    LocalMux I__1655 (
            .O(N__19397),
            .I(N__19394));
    Span4Mux_v I__1654 (
            .O(N__19394),
            .I(N__19391));
    Odrv4 I__1653 (
            .O(N__19391),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    CascadeMux I__1652 (
            .O(N__19388),
            .I(N__19385));
    InMux I__1651 (
            .O(N__19385),
            .I(N__19382));
    LocalMux I__1650 (
            .O(N__19382),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    InMux I__1649 (
            .O(N__19379),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__1648 (
            .O(N__19376),
            .I(N__19373));
    LocalMux I__1647 (
            .O(N__19373),
            .I(N__19370));
    Span4Mux_v I__1646 (
            .O(N__19370),
            .I(N__19367));
    Odrv4 I__1645 (
            .O(N__19367),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    CascadeMux I__1644 (
            .O(N__19364),
            .I(N__19361));
    InMux I__1643 (
            .O(N__19361),
            .I(N__19358));
    LocalMux I__1642 (
            .O(N__19358),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    InMux I__1641 (
            .O(N__19355),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    InMux I__1640 (
            .O(N__19352),
            .I(N__19349));
    LocalMux I__1639 (
            .O(N__19349),
            .I(N__19346));
    Span4Mux_v I__1638 (
            .O(N__19346),
            .I(N__19343));
    Odrv4 I__1637 (
            .O(N__19343),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__1636 (
            .O(N__19340),
            .I(N__19337));
    InMux I__1635 (
            .O(N__19337),
            .I(N__19334));
    LocalMux I__1634 (
            .O(N__19334),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    InMux I__1633 (
            .O(N__19331),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    InMux I__1632 (
            .O(N__19328),
            .I(N__19325));
    LocalMux I__1631 (
            .O(N__19325),
            .I(N__19322));
    Span4Mux_v I__1630 (
            .O(N__19322),
            .I(N__19319));
    Odrv4 I__1629 (
            .O(N__19319),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    InMux I__1628 (
            .O(N__19316),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    InMux I__1627 (
            .O(N__19313),
            .I(N__19310));
    LocalMux I__1626 (
            .O(N__19310),
            .I(N__19307));
    Span4Mux_v I__1625 (
            .O(N__19307),
            .I(N__19304));
    Odrv4 I__1624 (
            .O(N__19304),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    InMux I__1623 (
            .O(N__19301),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    InMux I__1622 (
            .O(N__19298),
            .I(N__19295));
    LocalMux I__1621 (
            .O(N__19295),
            .I(N__19292));
    Span4Mux_v I__1620 (
            .O(N__19292),
            .I(N__19289));
    Odrv4 I__1619 (
            .O(N__19289),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    InMux I__1618 (
            .O(N__19286),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    InMux I__1617 (
            .O(N__19283),
            .I(N__19280));
    LocalMux I__1616 (
            .O(N__19280),
            .I(N__19277));
    Span4Mux_v I__1615 (
            .O(N__19277),
            .I(N__19274));
    Odrv4 I__1614 (
            .O(N__19274),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    InMux I__1613 (
            .O(N__19271),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    InMux I__1612 (
            .O(N__19268),
            .I(N__19265));
    LocalMux I__1611 (
            .O(N__19265),
            .I(N__19262));
    Span4Mux_v I__1610 (
            .O(N__19262),
            .I(N__19259));
    Odrv4 I__1609 (
            .O(N__19259),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    InMux I__1608 (
            .O(N__19256),
            .I(bfn_1_12_0_));
    InMux I__1607 (
            .O(N__19253),
            .I(N__19250));
    LocalMux I__1606 (
            .O(N__19250),
            .I(N__19247));
    Span4Mux_v I__1605 (
            .O(N__19247),
            .I(N__19244));
    Odrv4 I__1604 (
            .O(N__19244),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    InMux I__1603 (
            .O(N__19241),
            .I(N__19238));
    LocalMux I__1602 (
            .O(N__19238),
            .I(N__19235));
    Span4Mux_v I__1601 (
            .O(N__19235),
            .I(N__19232));
    Odrv4 I__1600 (
            .O(N__19232),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__1599 (
            .O(N__19229),
            .I(N__19226));
    InMux I__1598 (
            .O(N__19226),
            .I(N__19223));
    LocalMux I__1597 (
            .O(N__19223),
            .I(N__19220));
    Odrv4 I__1596 (
            .O(N__19220),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    IoInMux I__1595 (
            .O(N__19217),
            .I(N__19214));
    LocalMux I__1594 (
            .O(N__19214),
            .I(N__19211));
    Span4Mux_s3_v I__1593 (
            .O(N__19211),
            .I(N__19208));
    Span4Mux_h I__1592 (
            .O(N__19208),
            .I(N__19205));
    Sp12to4 I__1591 (
            .O(N__19205),
            .I(N__19202));
    Span12Mux_v I__1590 (
            .O(N__19202),
            .I(N__19199));
    Span12Mux_v I__1589 (
            .O(N__19199),
            .I(N__19196));
    Odrv12 I__1588 (
            .O(N__19196),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1587 (
            .O(N__19193),
            .I(N__19190));
    LocalMux I__1586 (
            .O(N__19190),
            .I(N__19187));
    IoSpan4Mux I__1585 (
            .O(N__19187),
            .I(N__19184));
    IoSpan4Mux I__1584 (
            .O(N__19184),
            .I(N__19181));
    Odrv4 I__1583 (
            .O(N__19181),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_9_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_26_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_9_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_28_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_9_28_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_17_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_22_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_17_22_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_4_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_17_0_));
    defparam IN_MUX_bfv_4_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_4_18_0_));
    defparam IN_MUX_bfv_4_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_4_19_0_));
    defparam IN_MUX_bfv_4_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_4_20_0_));
    defparam IN_MUX_bfv_10_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_26_0_));
    defparam IN_MUX_bfv_10_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_27_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_10_27_0_));
    defparam IN_MUX_bfv_10_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_28_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_10_28_0_));
    defparam IN_MUX_bfv_3_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_23_0_));
    defparam IN_MUX_bfv_3_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_24_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_cry_7 ),
            .carryinitout(bfn_3_24_0_));
    defparam IN_MUX_bfv_1_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_24_0_));
    defparam IN_MUX_bfv_1_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_25_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_1_25_0_));
    defparam IN_MUX_bfv_1_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_26_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_1_26_0_));
    defparam IN_MUX_bfv_5_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_23_0_));
    defparam IN_MUX_bfv_5_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_24_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_5_24_0_));
    defparam IN_MUX_bfv_5_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_26_0_));
    defparam IN_MUX_bfv_5_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_27_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_5_27_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_16_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_5_0_));
    defparam IN_MUX_bfv_16_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_6_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_16_6_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_16_7_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_15 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_23 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .carryinitout(bfn_9_18_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19217),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19193),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__35558),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_162_i_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__31541),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un1_start_g ));
    ICE_GB \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0  (
            .USERSIGNALTOGLOBALBUFFER(N__36230),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_hc.un1_start_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__48437),
            .CLKHFEN(N__48439),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__48438),
            .RGB2PWM(N__24452),
            .RGB1(rgb_g),
            .CURREN(N__48404),
            .RGB2(rgb_b),
            .RGB1PWM(N__20864),
            .RGB0PWM(N__49574),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__19253),
            .in2(_gnd_net_),
            .in3(N__19493),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__19241),
            .in2(N__19229),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__19400),
            .in2(N__19388),
            .in3(N__19379),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__19376),
            .in2(N__19364),
            .in3(N__19355),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__19352),
            .in2(N__19340),
            .in3(N__19331),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__19328),
            .in2(N__19482),
            .in3(N__19316),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__19313),
            .in2(N__19484),
            .in3(N__19301),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__19298),
            .in2(N__19483),
            .in3(N__19286),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__19283),
            .in2(N__19485),
            .in3(N__19271),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__19268),
            .in2(N__19486),
            .in3(N__19256),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__19586),
            .in2(N__19490),
            .in3(N__19574),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__19571),
            .in2(N__19487),
            .in3(N__19559),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__19556),
            .in2(N__19491),
            .in3(N__19544),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__19541),
            .in2(N__19488),
            .in3(N__19526),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__19523),
            .in2(N__19492),
            .in3(N__19508),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__19505),
            .in2(N__19489),
            .in3(N__19406),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19403),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__21856),
            .in2(N__20797),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__21789),
            .in2(N__19736),
            .in3(N__19721),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__19718),
            .in2(N__21720),
            .in3(N__19709),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__21638),
            .in2(N__19706),
            .in3(N__19694),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__21576),
            .in2(N__19691),
            .in3(N__19676),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__21486),
            .in2(N__19673),
            .in3(N__19661),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__23345),
            .in2(N__19658),
            .in3(N__19643),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__22256),
            .in2(N__19640),
            .in3(N__19625),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__22194),
            .in2(N__19622),
            .in3(N__19607),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__22077),
            .in2(N__19604),
            .in3(N__19589),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__22032),
            .in2(N__19868),
            .in3(N__19856),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__21980),
            .in2(N__19853),
            .in3(N__19841),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__21918),
            .in2(N__19838),
            .in3(N__19823),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__22760),
            .in2(N__19820),
            .in3(N__19808),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__22694),
            .in2(N__19805),
            .in3(N__19790),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__22660),
            .in2(N__19787),
            .in3(N__19775),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__22608),
            .in2(N__19772),
            .in3(N__19757),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__22542),
            .in2(N__19754),
            .in3(N__19739),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__20021),
            .in2(N__22495),
            .in3(N__20009),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__20006),
            .in2(N__22435),
            .in3(N__19997),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__22367),
            .in2(N__19994),
            .in3(N__19979),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__23168),
            .in2(N__19976),
            .in3(N__19961),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__23111),
            .in2(N__19958),
            .in3(N__19943),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__23060),
            .in2(N__19940),
            .in3(N__19925),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__23010),
            .in2(N__19922),
            .in3(N__19907),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__22962),
            .in2(N__19904),
            .in3(N__19889),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__22911),
            .in2(N__19886),
            .in3(N__19871),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(N__22863),
            .in2(N__20120),
            .in3(N__20105),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(N__22819),
            .in2(N__20102),
            .in3(N__20090),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(N__23289),
            .in2(N__20087),
            .in3(N__20072),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_16_6  (
            .in0(N__20069),
            .in1(N__23762),
            .in2(N__20057),
            .in3(N__20045),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_1_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_1_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_1_17_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__24242),
            .in2(_gnd_net_),
            .in3(N__21855),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50267),
            .ce(),
            .sr(N__49536));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_17_3 .LUT_INIT=16'b1111111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_1_17_3  (
            .in0(N__23836),
            .in1(N__23704),
            .in2(N__23513),
            .in3(N__20042),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50267),
            .ce(),
            .sr(N__49536));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_1_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_1_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_1_17_6 .LUT_INIT=16'b1111010111100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_1_17_6  (
            .in0(N__23703),
            .in1(N__23476),
            .in2(N__20036),
            .in3(N__23838),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50267),
            .ce(),
            .sr(N__49536));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_1_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_1_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_1_17_7 .LUT_INIT=16'b1111111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_1_17_7  (
            .in0(N__23837),
            .in1(N__23705),
            .in2(N__23514),
            .in3(N__20027),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50267),
            .ce(),
            .sr(N__49536));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_1_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_1_20_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_1_20_4  (
            .in0(_gnd_net_),
            .in1(N__21442),
            .in2(_gnd_net_),
            .in3(N__22153),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_1_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_1_20_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_1_20_5  (
            .in0(N__21523),
            .in1(N__22234),
            .in2(N__20144),
            .in3(N__22309),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_21_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_21_2  (
            .in0(_gnd_net_),
            .in1(N__21605),
            .in2(_gnd_net_),
            .in3(N__21690),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_21_3 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_21_3  (
            .in0(N__20185),
            .in1(N__28452),
            .in2(N__20141),
            .in3(N__21059),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(\current_shift_inst.PI_CTRL.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_1_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_1_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_1_21_4 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_1_21_4  (
            .in0(N__21691),
            .in1(N__20135),
            .in2(N__20138),
            .in3(N__20203),
            .lcout(\current_shift_inst.PI_CTRL.N_161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_1_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_1_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_1_21_5 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_1_21_5  (
            .in0(N__20638),
            .in1(N__21607),
            .in2(N__20609),
            .in3(N__28451),
            .lcout(\current_shift_inst.PI_CTRL.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_21_6 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_21_6  (
            .in0(N__28453),
            .in1(N__21606),
            .in2(N__20608),
            .in3(N__20639),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_21_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_21_7  (
            .in0(N__20637),
            .in1(N__28450),
            .in2(_gnd_net_),
            .in3(N__20601),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_0  (
            .in0(N__20167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20129),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50212),
            .ce(),
            .sr(N__49548));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_1  (
            .in0(_gnd_net_),
            .in1(N__21764),
            .in2(_gnd_net_),
            .in3(N__20168),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50212),
            .ce(),
            .sr(N__49548));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_22_2 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_22_2  (
            .in0(N__21061),
            .in1(N__28465),
            .in2(N__20654),
            .in3(N__22154),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50212),
            .ce(),
            .sr(N__49548));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_4 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_4  (
            .in0(N__21695),
            .in1(N__20210),
            .in2(_gnd_net_),
            .in3(N__20204),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50212),
            .ce(),
            .sr(N__49548));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_5 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_5  (
            .in0(N__28464),
            .in1(N__21060),
            .in2(N__21530),
            .in3(N__20650),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50212),
            .ce(),
            .sr(N__49548));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_6 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_6  (
            .in0(N__21062),
            .in1(N__21611),
            .in2(N__20192),
            .in3(N__20174),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50212),
            .ce(),
            .sr(N__49548));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(N__24428),
            .in2(_gnd_net_),
            .in3(N__20166),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50212),
            .ce(),
            .sr(N__49548));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_23_0 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_23_0  (
            .in0(N__20651),
            .in1(N__28469),
            .in2(N__22238),
            .in3(N__21065),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50202),
            .ce(),
            .sr(N__49551));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_3 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_3  (
            .in0(N__28467),
            .in1(N__21063),
            .in2(N__21449),
            .in3(N__20652),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50202),
            .ce(),
            .sr(N__49551));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_23_5 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_23_5  (
            .in0(N__28468),
            .in1(N__21064),
            .in2(N__22316),
            .in3(N__20653),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50202),
            .ce(),
            .sr(N__49551));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_1_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_1_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_1_24_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_1_24_0  (
            .in0(N__20156),
            .in1(N__20150),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_1_24_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_1_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_1_24_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_1_24_1  (
            .in0(N__20306),
            .in1(N__20300),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_1_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_1_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_1_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_1_24_2  (
            .in0(_gnd_net_),
            .in1(N__20288),
            .in2(_gnd_net_),
            .in3(N__20294),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_1_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_1_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_1_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_1_24_3  (
            .in0(_gnd_net_),
            .in1(N__20276),
            .in2(_gnd_net_),
            .in3(N__20282),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_1_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_1_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_1_24_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_1_24_4  (
            .in0(_gnd_net_),
            .in1(N__20264),
            .in2(_gnd_net_),
            .in3(N__20270),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_1_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_1_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_1_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_1_24_5  (
            .in0(_gnd_net_),
            .in1(N__20252),
            .in2(_gnd_net_),
            .in3(N__20258),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_1_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_1_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_1_24_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_1_24_6  (
            .in0(_gnd_net_),
            .in1(N__20240),
            .in2(_gnd_net_),
            .in3(N__20246),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_1_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_1_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_1_24_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_1_24_7  (
            .in0(_gnd_net_),
            .in1(N__20228),
            .in2(_gnd_net_),
            .in3(N__20234),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_1_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_1_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_1_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_1_25_0  (
            .in0(_gnd_net_),
            .in1(N__20216),
            .in2(_gnd_net_),
            .in3(N__20222),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_1_25_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_1_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_1_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_1_25_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_1_25_1  (
            .in0(N__20342),
            .in1(N__20336),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_1_25_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_1_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_1_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_1_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23983),
            .in3(N__20330),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_1_25_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_1_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_1_25_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_1_25_3  (
            .in0(N__30519),
            .in1(N__28393),
            .in2(_gnd_net_),
            .in3(N__20327),
            .lcout(\pwm_generator_inst.un19_threshold_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_1_25_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_1_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_1_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_1_25_4  (
            .in0(_gnd_net_),
            .in1(N__21210),
            .in2(_gnd_net_),
            .in3(N__20324),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_1_25_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_1_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_1_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_1_25_5  (
            .in0(_gnd_net_),
            .in1(N__21393),
            .in2(_gnd_net_),
            .in3(N__20321),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_1_25_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_1_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_1_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_1_25_6  (
            .in0(_gnd_net_),
            .in1(N__20880),
            .in2(_gnd_net_),
            .in3(N__20318),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_1_25_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_1_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_1_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_1_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20531),
            .in3(N__20315),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_1_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_1_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_1_26_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_1_26_0  (
            .in0(_gnd_net_),
            .in1(N__20697),
            .in2(_gnd_net_),
            .in3(N__20312),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_26_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_1_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_1_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_1_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_1_26_1  (
            .in0(_gnd_net_),
            .in1(N__20676),
            .in2(_gnd_net_),
            .in3(N__20309),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_1_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_1_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_1_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_1_26_2  (
            .in0(_gnd_net_),
            .in1(N__20722),
            .in2(_gnd_net_),
            .in3(N__20399),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_1_26_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_1_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_1_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_1_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20396),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_13_0 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_2_13_0  (
            .in0(N__23699),
            .in1(N__20393),
            .in2(_gnd_net_),
            .in3(N__23460),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50305),
            .ce(),
            .sr(N__49517));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_2_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_2_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_2_13_3 .LUT_INIT=16'b1100110001000101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_2_13_3  (
            .in0(N__23877),
            .in1(N__20387),
            .in2(N__23509),
            .in3(N__23700),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50305),
            .ce(),
            .sr(N__49517));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_2_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_2_13_6 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_2_13_6  (
            .in0(N__23698),
            .in1(N__23878),
            .in2(N__20381),
            .in3(N__23459),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50305),
            .ce(),
            .sr(N__49517));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_2_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_2_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_2_14_2 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_2_14_2  (
            .in0(N__23849),
            .in1(N__23678),
            .in2(N__20372),
            .in3(N__23503),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50294),
            .ce(),
            .sr(N__49522));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_2_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_2_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_2_14_5 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_2_14_5  (
            .in0(N__23502),
            .in1(N__23850),
            .in2(N__23701),
            .in3(N__20363),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50294),
            .ce(),
            .sr(N__49522));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_0 .LUT_INIT=16'b1111111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_0  (
            .in0(N__23843),
            .in1(N__23658),
            .in2(N__23520),
            .in3(N__20357),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(N__49526));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_2_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_2_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_2_15_1 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_2_15_1  (
            .in0(N__23656),
            .in1(N__23848),
            .in2(N__20351),
            .in3(N__23501),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(N__49526));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_15_2 .LUT_INIT=16'b1111111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_2_15_2  (
            .in0(N__23842),
            .in1(N__23657),
            .in2(N__23519),
            .in3(N__20471),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(N__49526));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_2_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_2_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_2_15_4 .LUT_INIT=16'b1111111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_2_15_4  (
            .in0(N__23844),
            .in1(N__23659),
            .in2(N__23521),
            .in3(N__20465),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(N__49526));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_5 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_5  (
            .in0(N__23654),
            .in1(N__23846),
            .in2(N__20459),
            .in3(N__23499),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(N__49526));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_2_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_2_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_2_15_6 .LUT_INIT=16'b1111111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_2_15_6  (
            .in0(N__23845),
            .in1(N__23660),
            .in2(N__23522),
            .in3(N__20450),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(N__49526));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_2_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_2_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_2_15_7 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_2_15_7  (
            .in0(N__23655),
            .in1(N__23847),
            .in2(N__20444),
            .in3(N__23500),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(N__49526));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_2_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_2_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_2_16_0 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_2_16_0  (
            .in0(N__23454),
            .in1(N__23803),
            .in2(N__20435),
            .in3(N__23653),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(N__49530));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_16_4 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_2_16_4  (
            .in0(N__23452),
            .in1(N__23801),
            .in2(N__20426),
            .in3(N__23651),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(N__49530));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_2_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_2_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_2_16_5 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_2_16_5  (
            .in0(N__23800),
            .in1(N__23455),
            .in2(N__23689),
            .in3(N__20417),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(N__49530));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_16_6 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_2_16_6  (
            .in0(N__23453),
            .in1(N__23802),
            .in2(N__20411),
            .in3(N__23652),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(N__49530));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_1  (
            .in0(N__23350),
            .in1(N__22276),
            .in2(_gnd_net_),
            .in3(N__21572),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_2  (
            .in0(N__20891),
            .in1(N__22196),
            .in2(N__20507),
            .in3(N__21487),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_2_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_2_17_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_2_17_3  (
            .in0(N__20501),
            .in1(N__20495),
            .in2(N__20504),
            .in3(N__20660),
            .lcout(\current_shift_inst.PI_CTRL.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_17_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_17_5  (
            .in0(N__22765),
            .in1(N__22656),
            .in2(N__22039),
            .in3(N__21977),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_2_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_2_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_2_17_6  (
            .in0(N__22817),
            .in1(N__21919),
            .in2(N__22109),
            .in3(N__22705),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_2_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_2_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_2_18_0  (
            .in0(N__22612),
            .in1(N__22494),
            .in2(N__23179),
            .in3(N__22546),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_2_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_2_18_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_2_18_2  (
            .in0(N__22867),
            .in1(N__22907),
            .in2(N__23020),
            .in3(N__23293),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_2_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_2_18_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_2_18_5  (
            .in0(N__22371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22955),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_2_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_2_18_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_2_18_6  (
            .in0(N__22430),
            .in1(N__23064),
            .in2(N__20489),
            .in3(N__20486),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_2_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_2_18_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_2_18_7  (
            .in0(N__23116),
            .in1(N__23761),
            .in2(N__20480),
            .in3(N__20477),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_2_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_2_19_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_2_19_1  (
            .in0(N__22431),
            .in1(N__23065),
            .in2(N__22384),
            .in3(N__23804),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_19_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_19_4  (
            .in0(N__20948),
            .in1(N__20954),
            .in2(N__21008),
            .in3(N__21089),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_21_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_21_0  (
            .in0(_gnd_net_),
            .in1(N__22149),
            .in2(_gnd_net_),
            .in3(N__21522),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_21_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_21_1  (
            .in0(N__22233),
            .in1(N__22308),
            .in2(N__20612),
            .in3(N__21441),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_22_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_22_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_22_7  (
            .in0(N__20587),
            .in1(N__20569),
            .in2(_gnd_net_),
            .in3(N__20554),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_23_3  (
            .in0(_gnd_net_),
            .in1(N__23976),
            .in2(_gnd_net_),
            .in3(N__23941),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_2_24_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_2_24_0 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_2_24_0  (
            .in0(N__20537),
            .in1(N__28280),
            .in2(N__30520),
            .in3(N__20885),
            .lcout(\pwm_generator_inst.un19_threshold_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_24_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_24_1  (
            .in0(N__20530),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28255),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_2_24_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_2_24_2 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_2_24_2  (
            .in0(N__20516),
            .in1(N__28256),
            .in2(N__20510),
            .in3(N__30503),
            .lcout(\pwm_generator_inst.un19_threshold_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_2_24_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_2_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_2_24_4 .LUT_INIT=16'b1011011110000100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_2_24_4  (
            .in0(N__20747),
            .in1(N__30502),
            .in2(N__20705),
            .in3(N__28232),
            .lcout(\pwm_generator_inst.un19_threshold_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_24_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_24_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_24_5  (
            .in0(_gnd_net_),
            .in1(N__21240),
            .in2(_gnd_net_),
            .in3(N__24109),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_2_24_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_2_24_6 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_2_24_6  (
            .in0(N__20738),
            .in1(N__28559),
            .in2(N__30521),
            .in3(N__20681),
            .lcout(\pwm_generator_inst.un19_threshold_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_2_25_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_2_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_2_25_1 .LUT_INIT=16'b1011100001110100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_2_25_1  (
            .in0(N__20721),
            .in1(N__30500),
            .in2(N__28535),
            .in3(N__20729),
            .lcout(\pwm_generator_inst.un19_threshold_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_26_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_26_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_26_0  (
            .in0(N__28525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20723),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_26_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_26_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_26_1  (
            .in0(_gnd_net_),
            .in1(N__20701),
            .in2(_gnd_net_),
            .in3(N__28225),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_26_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_26_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_26_3  (
            .in0(N__20680),
            .in1(N__28552),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_26_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_26_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_26_4  (
            .in0(_gnd_net_),
            .in1(N__28318),
            .in2(_gnd_net_),
            .in3(N__21397),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_26_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_26_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_26_6  (
            .in0(_gnd_net_),
            .in1(N__28357),
            .in2(_gnd_net_),
            .in3(N__21212),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_2_26_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_2_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_2_26_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_2_26_7  (
            .in0(N__28273),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20884),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_LC_2_29_7.C_ON=1'b0;
    defparam rgb_drv_RNO_LC_2_29_7.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_LC_2_29_7.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_drv_RNO_LC_2_29_7 (
            .in0(N__49573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33560),
            .lcout(rgb_drv_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_13_2 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_3_13_2  (
            .in0(N__23873),
            .in1(N__23684),
            .in2(N__20852),
            .in3(N__23516),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50295),
            .ce(),
            .sr(N__49515));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_13_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_3_13_4  (
            .in0(N__20837),
            .in1(N__23685),
            .in2(_gnd_net_),
            .in3(N__23517),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50295),
            .ce(),
            .sr(N__49515));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_3_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_3_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_3_13_6 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_3_13_6  (
            .in0(N__23872),
            .in1(N__23683),
            .in2(N__20828),
            .in3(N__23515),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50295),
            .ce(),
            .sr(N__49515));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_3_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_3_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_3_14_2 .LUT_INIT=16'b1101000011010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_3_14_2  (
            .in0(N__23868),
            .in1(N__23682),
            .in2(N__20813),
            .in3(N__23508),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50282),
            .ce(),
            .sr(N__49518));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_3_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_3_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_3_14_5 .LUT_INIT=16'b0011001011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_3_14_5  (
            .in0(N__23507),
            .in1(N__21847),
            .in2(N__23702),
            .in3(N__20798),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50282),
            .ce(),
            .sr(N__49518));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_3_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_3_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_3_15_2 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_3_15_2  (
            .in0(N__23865),
            .in1(N__23646),
            .in2(N__20774),
            .in3(N__23506),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50270),
            .ce(),
            .sr(N__49523));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_15_3 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_3_15_3  (
            .in0(N__23504),
            .in1(N__23867),
            .in2(N__23688),
            .in3(N__20759),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50270),
            .ce(),
            .sr(N__49523));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_3_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_3_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_3_15_4 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_3_15_4  (
            .in0(N__23866),
            .in1(N__23505),
            .in2(N__20933),
            .in3(N__23647),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50270),
            .ce(),
            .sr(N__49523));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_3_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_3_15_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_3_15_7  (
            .in0(N__22487),
            .in1(N__22541),
            .in2(N__23175),
            .in3(N__22604),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_16_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_16_0  (
            .in0(N__22269),
            .in1(N__23349),
            .in2(N__22190),
            .in3(N__21479),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_16_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_16_1  (
            .in0(N__21654),
            .in1(N__21578),
            .in2(N__20921),
            .in3(N__21735),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_3_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_3_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_3_16_2  (
            .in0(N__22818),
            .in1(N__23112),
            .in2(N__20918),
            .in3(N__20915),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_3  (
            .in0(N__20975),
            .in1(N__20897),
            .in2(N__20909),
            .in3(N__20906),
            .lcout(\current_shift_inst.PI_CTRL.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_5  (
            .in0(N__22862),
            .in1(N__23009),
            .in2(N__22925),
            .in3(N__22969),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_3_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_3_17_0 .LUT_INIT=16'b0000001100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_3_17_0  (
            .in0(N__21848),
            .in1(N__21739),
            .in2(N__21656),
            .in3(N__21793),
            .lcout(\current_shift_inst.PI_CTRL.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_3_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_3_17_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_3_17_3  (
            .in0(N__22704),
            .in1(N__21911),
            .in2(N__22105),
            .in3(N__22655),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_17_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_17_4  (
            .in0(N__21978),
            .in1(N__20969),
            .in2(N__20978),
            .in3(N__23288),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_3_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_3_17_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__22764),
            .in2(_gnd_net_),
            .in3(N__22022),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_3_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_3_18_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_3_18_1  (
            .in0(N__22627),
            .in1(N__22675),
            .in2(N__22796),
            .in3(N__22060),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_3_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_3_18_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_3_18_5  (
            .in0(N__22628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22676),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_3_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_3_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_3_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__21946),
            .in2(_gnd_net_),
            .in3(N__22061),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_3_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_3_19_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__22513),
            .in2(_gnd_net_),
            .in3(N__22576),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_3_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_3_19_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_3_19_1  (
            .in0(N__21991),
            .in1(N__21947),
            .in2(N__20963),
            .in3(N__20960),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_3_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_3_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_3_19_2  (
            .in0(N__23036),
            .in1(N__22726),
            .in2(N__23087),
            .in3(N__21874),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_3_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_3_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_3_19_3  (
            .in0(N__22343),
            .in1(N__23086),
            .in2(N__22795),
            .in3(N__23035),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_3_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_3_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_3_19_4  (
            .in0(N__22838),
            .in1(N__21992),
            .in2(N__20942),
            .in3(N__20939),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_3_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_3_19_6 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_3_19_6  (
            .in0(N__22339),
            .in1(N__23137),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_3_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_3_19_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_3_19_7  (
            .in0(N__22885),
            .in1(N__22837),
            .in2(N__21092),
            .in3(N__23263),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_3_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_3_20_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_3_20_0  (
            .in0(N__22985),
            .in1(N__21083),
            .in2(N__23141),
            .in3(N__22937),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_20_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_20_1  (
            .in0(N__20999),
            .in1(N__21014),
            .in2(N__21074),
            .in3(N__21071),
            .lcout(\current_shift_inst.PI_CTRL.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_3_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_3_20_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_3_20_4  (
            .in0(N__22463),
            .in1(N__21878),
            .in2(N__22736),
            .in3(N__22402),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_3_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_3_20_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_3_20_5  (
            .in0(N__22936),
            .in1(N__22984),
            .in2(N__22403),
            .in3(N__22462),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_3_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_3_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_3_20_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_3_20_7  (
            .in0(N__23264),
            .in1(N__22577),
            .in2(N__22517),
            .in3(N__22886),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_23_0  (
            .in0(_gnd_net_),
            .in1(N__23918),
            .in2(N__30529),
            .in3(N__30525),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ),
            .ltout(),
            .carryin(bfn_3_23_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_23_1  (
            .in0(_gnd_net_),
            .in1(N__20993),
            .in2(_gnd_net_),
            .in3(N__20981),
            .lcout(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_23_2  (
            .in0(_gnd_net_),
            .in1(N__21194),
            .in2(_gnd_net_),
            .in3(N__21158),
            .lcout(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_23_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_23_3  (
            .in0(_gnd_net_),
            .in1(N__21362),
            .in2(_gnd_net_),
            .in3(N__21155),
            .lcout(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_23_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_23_4  (
            .in0(_gnd_net_),
            .in1(N__21152),
            .in2(_gnd_net_),
            .in3(N__21146),
            .lcout(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_23_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_23_5  (
            .in0(_gnd_net_),
            .in1(N__21143),
            .in2(_gnd_net_),
            .in3(N__21137),
            .lcout(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_23_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_23_6  (
            .in0(_gnd_net_),
            .in1(N__21134),
            .in2(_gnd_net_),
            .in3(N__21128),
            .lcout(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_23_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_23_7  (
            .in0(_gnd_net_),
            .in1(N__21125),
            .in2(_gnd_net_),
            .in3(N__21119),
            .lcout(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_24_0  (
            .in0(_gnd_net_),
            .in1(N__21116),
            .in2(_gnd_net_),
            .in3(N__21110),
            .lcout(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ),
            .ltout(),
            .carryin(bfn_3_24_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_24_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_24_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_24_1  (
            .in0(N__21107),
            .in1(N__28508),
            .in2(N__30530),
            .in3(N__21095),
            .lcout(),
            .ltout(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_3_24_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_3_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_3_24_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_3_24_2  (
            .in0(N__32424),
            .in1(N__24077),
            .in2(N__21401),
            .in3(N__24040),
            .lcout(\pwm_generator_inst.threshold_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_3_24_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_3_24_3 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_3_24_3  (
            .in0(N__28319),
            .in1(N__21398),
            .in2(N__21377),
            .in3(N__30501),
            .lcout(\pwm_generator_inst.un19_threshold_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_24_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_24_5 .LUT_INIT=16'b1010111110101011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_3_24_5  (
            .in0(N__21341),
            .in1(N__24172),
            .in2(N__24146),
            .in3(N__21356),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_24_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_24_6 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_24_6  (
            .in0(N__21347),
            .in1(N__21334),
            .in2(N__21311),
            .in3(N__21277),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_24_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_24_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_24_7  (
            .in0(N__21335),
            .in1(N__21310),
            .in2(N__21281),
            .in3(N__21251),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_3_25_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_3_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_3_25_4 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_3_25_4  (
            .in0(N__21221),
            .in1(N__21211),
            .in2(N__28364),
            .in3(N__30499),
            .lcout(\pwm_generator_inst.un19_threshold_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_4_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_4_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_4_13_4 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_4_13_4  (
            .in0(N__23879),
            .in1(N__23687),
            .in2(N__21185),
            .in3(N__23518),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50283),
            .ce(),
            .sr(N__49510));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_14_4 .LUT_INIT=16'b1101000011010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_4_14_4  (
            .in0(N__23870),
            .in1(N__23686),
            .in2(N__21173),
            .in3(N__23511),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50271),
            .ce(),
            .sr(N__49516));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27673),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(N__49519));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_4_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_4_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_4_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27295),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(N__49519));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_4_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_4_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_4_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27700),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(N__49519));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_4_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_4_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_4_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27352),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(N__49519));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_4_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_4_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_4_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27592),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(N__49519));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27497),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(N__49519));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_4_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_4_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_4_15_7 .LUT_INIT=16'b1111000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_4_15_7  (
            .in0(N__23869),
            .in1(N__23510),
            .in2(N__21416),
            .in3(N__23661),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(N__49519));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_4_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_4_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_4_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27328),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50247),
            .ce(),
            .sr(N__49524));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27275),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50247),
            .ce(),
            .sr(N__49524));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_4_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_4_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_4_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27733),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50247),
            .ce(),
            .sr(N__49524));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_4_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_4_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_4_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27799),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50247),
            .ce(),
            .sr(N__49524));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27550),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50247),
            .ce(),
            .sr(N__49524));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_4_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_4_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_4_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_4_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27863),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50247),
            .ce(),
            .sr(N__49524));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_4_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_4_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_4_17_0  (
            .in0(_gnd_net_),
            .in1(N__24238),
            .in2(N__21860),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_17_1  (
            .in0(_gnd_net_),
            .in1(N__21806),
            .in2(N__21797),
            .in3(N__21749),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__50235),
            .ce(),
            .sr(N__49527));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_17_2  (
            .in0(_gnd_net_),
            .in1(N__21746),
            .in2(N__21740),
            .in3(N__21668),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__50235),
            .ce(),
            .sr(N__49527));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_17_3  (
            .in0(_gnd_net_),
            .in1(N__21665),
            .in2(N__21655),
            .in3(N__21581),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__50235),
            .ce(),
            .sr(N__49527));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(N__21577),
            .in2(N__21539),
            .in3(N__21500),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__50235),
            .ce(),
            .sr(N__49527));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_17_5  (
            .in0(_gnd_net_),
            .in1(N__21497),
            .in2(N__21488),
            .in3(N__21419),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__50235),
            .ce(),
            .sr(N__49527));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_17_6  (
            .in0(_gnd_net_),
            .in1(N__22325),
            .in2(N__23351),
            .in3(N__22280),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__50235),
            .ce(),
            .sr(N__49527));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_17_7  (
            .in0(_gnd_net_),
            .in1(N__22277),
            .in2(N__24263),
            .in3(N__22199),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__50235),
            .ce(),
            .sr(N__49527));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__24227),
            .in2(N__22195),
            .in3(N__22121),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_4_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__50224),
            .ce(),
            .sr(N__49531));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_18_1  (
            .in0(_gnd_net_),
            .in1(N__22118),
            .in2(N__22104),
            .in3(N__22052),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__50224),
            .ce(),
            .sr(N__49531));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_18_2  (
            .in0(_gnd_net_),
            .in1(N__22049),
            .in2(N__22040),
            .in3(N__21983),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__50224),
            .ce(),
            .sr(N__49531));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(N__21979),
            .in2(N__24254),
            .in3(N__21935),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__50224),
            .ce(),
            .sr(N__49531));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(N__21932),
            .in2(N__21923),
            .in3(N__21863),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__50224),
            .ce(),
            .sr(N__49531));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_18_5  (
            .in0(_gnd_net_),
            .in1(N__24221),
            .in2(N__22772),
            .in3(N__22715),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__50224),
            .ce(),
            .sr(N__49531));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_18_6  (
            .in0(_gnd_net_),
            .in1(N__24326),
            .in2(N__22712),
            .in3(N__22667),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__50224),
            .ce(),
            .sr(N__49531));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_18_7  (
            .in0(_gnd_net_),
            .in1(N__24215),
            .in2(N__22664),
            .in3(N__22619),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__50224),
            .ce(),
            .sr(N__49531));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_19_0  (
            .in0(_gnd_net_),
            .in1(N__24296),
            .in2(N__22616),
            .in3(N__22565),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_4_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__50213),
            .ce(),
            .sr(N__49534));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_19_1  (
            .in0(_gnd_net_),
            .in1(N__22562),
            .in2(N__22553),
            .in3(N__22502),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__50213),
            .ce(),
            .sr(N__49534));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_19_2  (
            .in0(_gnd_net_),
            .in1(N__22499),
            .in2(N__24209),
            .in3(N__22454),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__50213),
            .ce(),
            .sr(N__49534));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_19_3  (
            .in0(_gnd_net_),
            .in1(N__22451),
            .in2(N__22442),
            .in3(N__22391),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__50213),
            .ce(),
            .sr(N__49534));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(N__24200),
            .in2(N__22388),
            .in3(N__22328),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__50213),
            .ce(),
            .sr(N__49534));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_19_5  (
            .in0(_gnd_net_),
            .in1(N__23192),
            .in2(N__23183),
            .in3(N__23126),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__50213),
            .ce(),
            .sr(N__49534));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(N__24308),
            .in2(N__23123),
            .in3(N__23075),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__50213),
            .ce(),
            .sr(N__49534));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_19_7  (
            .in0(_gnd_net_),
            .in1(N__24302),
            .in2(N__23072),
            .in3(N__23027),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__50213),
            .ce(),
            .sr(N__49534));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_20_0  (
            .in0(_gnd_net_),
            .in1(N__24275),
            .in2(N__23024),
            .in3(N__22976),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_4_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__50203),
            .ce(),
            .sr(N__49537));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(N__24281),
            .in2(N__22973),
            .in3(N__22928),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__50203),
            .ce(),
            .sr(N__49537));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_20_2  (
            .in0(_gnd_net_),
            .in1(N__22924),
            .in2(N__24194),
            .in3(N__22874),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__50203),
            .ce(),
            .sr(N__49537));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_20_3  (
            .in0(_gnd_net_),
            .in1(N__22871),
            .in2(N__24320),
            .in3(N__22829),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__50203),
            .ce(),
            .sr(N__49537));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(N__22826),
            .in2(N__24290),
            .in3(N__22775),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__50203),
            .ce(),
            .sr(N__49537));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_20_5  (
            .in0(_gnd_net_),
            .in1(N__24269),
            .in2(N__23300),
            .in3(N__23252),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__50203),
            .ce(),
            .sr(N__49537));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_20_6  (
            .in0(N__23851),
            .in1(N__28478),
            .in2(_gnd_net_),
            .in3(N__23249),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50203),
            .ce(),
            .sr(N__49537));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_4_23_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_4_23_0 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_4_23_0  (
            .in0(N__24071),
            .in1(N__32391),
            .in2(N__24042),
            .in3(N__23246),
            .lcout(\pwm_generator_inst.threshold_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_4_23_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_4_23_1 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_4_23_1  (
            .in0(N__32393),
            .in1(N__24073),
            .in2(N__23240),
            .in3(N__24033),
            .lcout(\pwm_generator_inst.threshold_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_4_23_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_4_23_2 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_4_23_2  (
            .in0(N__24072),
            .in1(N__32392),
            .in2(N__24043),
            .in3(N__23231),
            .lcout(\pwm_generator_inst.threshold_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_4_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_4_23_3 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_4_23_3  (
            .in0(N__32394),
            .in1(N__24074),
            .in2(N__23225),
            .in3(N__24034),
            .lcout(\pwm_generator_inst.threshold_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_4_23_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_4_23_4 .LUT_INIT=16'b1111111101000111;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_4_23_4  (
            .in0(N__24075),
            .in1(N__32395),
            .in2(N__24044),
            .in3(N__23216),
            .lcout(\pwm_generator_inst.un14_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_4_23_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_4_23_5 .LUT_INIT=16'b1111001011110111;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_4_23_5  (
            .in0(N__32390),
            .in1(N__24070),
            .in2(N__23210),
            .in3(N__24026),
            .lcout(\pwm_generator_inst.un14_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_4_23_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_4_23_6 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_4_23_6  (
            .in0(N__24069),
            .in1(N__32389),
            .in2(N__24041),
            .in3(N__23198),
            .lcout(\pwm_generator_inst.threshold_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_4_23_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_4_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_4_23_7 .LUT_INIT=16'b1111001011110111;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_4_23_7  (
            .in0(N__32396),
            .in1(N__24076),
            .in2(N__24182),
            .in3(N__24038),
            .lcout(\pwm_generator_inst.un14_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_24_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_24_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_24_6  (
            .in0(N__24173),
            .in1(N__24142),
            .in2(N__24116),
            .in3(N__24083),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(\pwm_generator_inst.N_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_4_24_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_4_24_7 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_4_24_7  (
            .in0(N__24039),
            .in1(N__23993),
            .in2(N__23987),
            .in3(N__32423),
            .lcout(\pwm_generator_inst.un14_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_7 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_7  (
            .in0(N__23984),
            .in1(N__23954),
            .in2(N__23945),
            .in3(N__30498),
            .lcout(\pwm_generator_inst.un19_threshold_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_4_30_3.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_4_30_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_4_30_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_4_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23906),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_5_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_5_10_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_5_10_1  (
            .in0(N__29074),
            .in1(N__29106),
            .in2(_gnd_net_),
            .in3(N__34816),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_5_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_5_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_5_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_28_LC_5_11_4  (
            .in0(N__29111),
            .in1(N__29070),
            .in2(_gnd_net_),
            .in3(N__34817),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50296),
            .ce(N__29767),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_5_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_5_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_5_14_0 .LUT_INIT=16'b1101000011010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_5_14_0  (
            .in0(N__23871),
            .in1(N__23690),
            .in2(N__23537),
            .in3(N__23512),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50260),
            .ce(),
            .sr(N__49511));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_16_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_5_16_5  (
            .in0(N__27649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50236),
            .ce(),
            .sr(N__49520));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_16_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(N__27520),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50236),
            .ce(),
            .sr(N__49520));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27386),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50225),
            .ce(),
            .sr(N__49525));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_5_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27622),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50225),
            .ce(),
            .sr(N__49525));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27466),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50225),
            .ce(),
            .sr(N__49525));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_17_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_5_17_7  (
            .in0(_gnd_net_),
            .in1(N__27922),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50225),
            .ce(),
            .sr(N__49525));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27826),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50214),
            .ce(),
            .sr(N__49528));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_5_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_5_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_5_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27764),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50214),
            .ce(),
            .sr(N__49528));
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_5_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_5_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_5_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_27_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28075),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50214),
            .ce(),
            .sr(N__49528));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27955),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50214),
            .ce(),
            .sr(N__49528));
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_5_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_5_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_5_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_28_LC_5_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28048),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50214),
            .ce(),
            .sr(N__49528));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_5_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28201),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50214),
            .ce(),
            .sr(N__49528));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28171),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50204),
            .ce(),
            .sr(N__49532));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27892),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50204),
            .ce(),
            .sr(N__49532));
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_5_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_5_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_5_19_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_29_LC_5_19_4  (
            .in0(N__28025),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50204),
            .ce(),
            .sr(N__49532));
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_5_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_5_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_5_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_26_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28111),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50204),
            .ce(),
            .sr(N__49532));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_5_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28142),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50195),
            .ce(),
            .sr(N__49535));
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_5_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_5_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_5_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_30_LC_5_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27991),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50195),
            .ce(),
            .sr(N__49535));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_5_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_5_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_5_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_5_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29725),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50189),
            .ce(),
            .sr(N__49538));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24434),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50185),
            .ce(),
            .sr(N__49540));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_23_0  (
            .in0(_gnd_net_),
            .in1(N__24410),
            .in2(N__24419),
            .in3(N__24710),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_5_23_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_23_1  (
            .in0(_gnd_net_),
            .in1(N__24395),
            .in2(N__24404),
            .in3(N__24686),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_23_2  (
            .in0(_gnd_net_),
            .in1(N__24380),
            .in2(N__24389),
            .in3(N__24662),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_23_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_23_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_23_3  (
            .in0(N__24638),
            .in1(N__24362),
            .in2(N__24371),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_23_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_23_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_23_4  (
            .in0(_gnd_net_),
            .in1(N__24356),
            .in2(N__24350),
            .in3(N__24614),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_23_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_23_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_23_5  (
            .in0(N__24590),
            .in1(N__24332),
            .in2(N__24341),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_23_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_23_6  (
            .in0(_gnd_net_),
            .in1(N__24533),
            .in2(N__24542),
            .in3(N__24566),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_23_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_23_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_23_7  (
            .in0(_gnd_net_),
            .in1(N__24527),
            .in2(N__24521),
            .in3(N__24854),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_24_0  (
            .in0(_gnd_net_),
            .in1(N__24503),
            .in2(N__24512),
            .in3(N__24830),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_5_24_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_24_1  (
            .in0(_gnd_net_),
            .in1(N__24485),
            .in2(N__24497),
            .in3(N__24758),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_5_24_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_5_24_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_5_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_5_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24479),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50180),
            .ce(),
            .sr(N__49544));
    defparam rgb_drv_RNO_0_LC_5_25_0.C_ON=1'b0;
    defparam rgb_drv_RNO_0_LC_5_25_0.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_0_LC_5_25_0.LUT_INIT=16'b1010101001010101;
    LogicCell40 rgb_drv_RNO_0_LC_5_25_0 (
            .in0(N__49572),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33553),
            .lcout(N_38_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_5_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_5_25_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_5_25_2  (
            .in0(N__24757),
            .in1(N__24829),
            .in2(_gnd_net_),
            .in3(N__24852),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto9_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_5_25_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_5_25_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_5_25_3  (
            .in0(N__24565),
            .in1(N__24589),
            .in2(N__24437),
            .in3(N__24716),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_5_25_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_5_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_5_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_5_25_5  (
            .in0(_gnd_net_),
            .in1(N__24705),
            .in2(_gnd_net_),
            .in3(N__24657),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_5_25_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_5_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_5_25_6 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_5_25_6  (
            .in0(N__24612),
            .in1(N__24684),
            .in2(N__24719),
            .in3(N__24636),
            .lcout(\pwm_generator_inst.un1_counterlt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_5_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_5_26_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_5_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_5_26_0  (
            .in0(N__24800),
            .in1(N__24709),
            .in2(_gnd_net_),
            .in3(N__24689),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_26_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__50176),
            .ce(),
            .sr(N__49549));
    defparam \pwm_generator_inst.counter_1_LC_5_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_5_26_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_5_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_5_26_1  (
            .in0(N__24794),
            .in1(N__24685),
            .in2(_gnd_net_),
            .in3(N__24665),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__50176),
            .ce(),
            .sr(N__49549));
    defparam \pwm_generator_inst.counter_2_LC_5_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_5_26_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_5_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_5_26_2  (
            .in0(N__24801),
            .in1(N__24661),
            .in2(_gnd_net_),
            .in3(N__24641),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__50176),
            .ce(),
            .sr(N__49549));
    defparam \pwm_generator_inst.counter_3_LC_5_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_5_26_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_5_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_5_26_3  (
            .in0(N__24795),
            .in1(N__24637),
            .in2(_gnd_net_),
            .in3(N__24617),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__50176),
            .ce(),
            .sr(N__49549));
    defparam \pwm_generator_inst.counter_4_LC_5_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_5_26_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_5_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_5_26_4  (
            .in0(N__24802),
            .in1(N__24613),
            .in2(_gnd_net_),
            .in3(N__24593),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__50176),
            .ce(),
            .sr(N__49549));
    defparam \pwm_generator_inst.counter_5_LC_5_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_5_26_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_5_26_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_5_26_5  (
            .in0(N__24796),
            .in1(N__24588),
            .in2(_gnd_net_),
            .in3(N__24569),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__50176),
            .ce(),
            .sr(N__49549));
    defparam \pwm_generator_inst.counter_6_LC_5_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_5_26_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_5_26_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_5_26_6  (
            .in0(N__24803),
            .in1(N__24564),
            .in2(_gnd_net_),
            .in3(N__24545),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__50176),
            .ce(),
            .sr(N__49549));
    defparam \pwm_generator_inst.counter_7_LC_5_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_5_26_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_5_26_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_5_26_7  (
            .in0(N__24797),
            .in1(N__24853),
            .in2(_gnd_net_),
            .in3(N__24833),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__50176),
            .ce(),
            .sr(N__49549));
    defparam \pwm_generator_inst.counter_8_LC_5_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_5_27_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_5_27_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_5_27_0  (
            .in0(N__24799),
            .in1(N__24828),
            .in2(_gnd_net_),
            .in3(N__24806),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_27_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__50173),
            .ce(),
            .sr(N__49552));
    defparam \pwm_generator_inst.counter_9_LC_5_27_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_5_27_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_5_27_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_5_27_1  (
            .in0(N__24756),
            .in1(N__24798),
            .in2(_gnd_net_),
            .in3(N__24761),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50173),
            .ce(),
            .sr(N__49552));
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_7_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_7_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_7_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_29_LC_7_6_5  (
            .in0(N__34758),
            .in1(N__28907),
            .in2(_gnd_net_),
            .in3(N__28886),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50319),
            .ce(N__29760),
            .sr(N__49460));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_7_0  (
            .in0(N__25075),
            .in1(N__25485),
            .in2(_gnd_net_),
            .in3(N__24734),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__50314),
            .ce(N__25160),
            .sr(N__49468));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_7_1  (
            .in0(N__25067),
            .in1(N__25464),
            .in2(_gnd_net_),
            .in3(N__24731),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__50314),
            .ce(N__25160),
            .sr(N__49468));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_7_2  (
            .in0(N__25076),
            .in1(N__25441),
            .in2(_gnd_net_),
            .in3(N__24728),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__50314),
            .ce(N__25160),
            .sr(N__49468));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_7_3  (
            .in0(N__25068),
            .in1(N__25417),
            .in2(_gnd_net_),
            .in3(N__24725),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__50314),
            .ce(N__25160),
            .sr(N__49468));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_7_4  (
            .in0(N__25077),
            .in1(N__25393),
            .in2(_gnd_net_),
            .in3(N__24722),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__50314),
            .ce(N__25160),
            .sr(N__49468));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_7_5  (
            .in0(N__25069),
            .in1(N__25369),
            .in2(_gnd_net_),
            .in3(N__24881),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__50314),
            .ce(N__25160),
            .sr(N__49468));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_7_6  (
            .in0(N__25078),
            .in1(N__25345),
            .in2(_gnd_net_),
            .in3(N__24878),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__50314),
            .ce(N__25160),
            .sr(N__49468));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_7_7  (
            .in0(N__25070),
            .in1(N__25321),
            .in2(_gnd_net_),
            .in3(N__24875),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__50314),
            .ce(N__25160),
            .sr(N__49468));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_8_0  (
            .in0(N__25066),
            .in1(N__25297),
            .in2(_gnd_net_),
            .in3(N__24872),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__50306),
            .ce(N__25149),
            .sr(N__49475));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_8_1  (
            .in0(N__25102),
            .in1(N__25678),
            .in2(_gnd_net_),
            .in3(N__24869),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__50306),
            .ce(N__25149),
            .sr(N__49475));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_8_2  (
            .in0(N__25063),
            .in1(N__25654),
            .in2(_gnd_net_),
            .in3(N__24866),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__50306),
            .ce(N__25149),
            .sr(N__49475));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_8_3  (
            .in0(N__25099),
            .in1(N__25630),
            .in2(_gnd_net_),
            .in3(N__24863),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__50306),
            .ce(N__25149),
            .sr(N__49475));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_8_4  (
            .in0(N__25064),
            .in1(N__25606),
            .in2(_gnd_net_),
            .in3(N__24860),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__50306),
            .ce(N__25149),
            .sr(N__49475));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_8_5  (
            .in0(N__25100),
            .in1(N__25582),
            .in2(_gnd_net_),
            .in3(N__24857),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__50306),
            .ce(N__25149),
            .sr(N__49475));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_8_6  (
            .in0(N__25065),
            .in1(N__25558),
            .in2(_gnd_net_),
            .in3(N__24908),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__50306),
            .ce(N__25149),
            .sr(N__49475));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_8_7  (
            .in0(N__25101),
            .in1(N__25534),
            .in2(_gnd_net_),
            .in3(N__24905),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__50306),
            .ce(N__25149),
            .sr(N__49475));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_9_0  (
            .in0(N__25079),
            .in1(N__25510),
            .in2(_gnd_net_),
            .in3(N__24902),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__50297),
            .ce(N__25156),
            .sr(N__49482));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_9_1  (
            .in0(N__25095),
            .in1(N__25891),
            .in2(_gnd_net_),
            .in3(N__24899),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__50297),
            .ce(N__25156),
            .sr(N__49482));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_9_2  (
            .in0(N__25080),
            .in1(N__25867),
            .in2(_gnd_net_),
            .in3(N__24896),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__50297),
            .ce(N__25156),
            .sr(N__49482));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_9_3  (
            .in0(N__25096),
            .in1(N__25843),
            .in2(_gnd_net_),
            .in3(N__24893),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__50297),
            .ce(N__25156),
            .sr(N__49482));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_9_4  (
            .in0(N__25081),
            .in1(N__25819),
            .in2(_gnd_net_),
            .in3(N__24890),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__50297),
            .ce(N__25156),
            .sr(N__49482));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_9_5  (
            .in0(N__25097),
            .in1(N__25795),
            .in2(_gnd_net_),
            .in3(N__24887),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__50297),
            .ce(N__25156),
            .sr(N__49482));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_9_6  (
            .in0(N__25082),
            .in1(N__25771),
            .in2(_gnd_net_),
            .in3(N__24884),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__50297),
            .ce(N__25156),
            .sr(N__49482));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_9_7  (
            .in0(N__25098),
            .in1(N__25747),
            .in2(_gnd_net_),
            .in3(N__24929),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__50297),
            .ce(N__25156),
            .sr(N__49482));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_10_0  (
            .in0(N__25071),
            .in1(N__25723),
            .in2(_gnd_net_),
            .in3(N__24926),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__50284),
            .ce(N__25148),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_10_1  (
            .in0(N__25108),
            .in1(N__25699),
            .in2(_gnd_net_),
            .in3(N__24923),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__50284),
            .ce(N__25148),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_10_2  (
            .in0(N__25072),
            .in1(N__25984),
            .in2(_gnd_net_),
            .in3(N__24920),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__50284),
            .ce(N__25148),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_10_3  (
            .in0(N__25109),
            .in1(N__25948),
            .in2(_gnd_net_),
            .in3(N__24917),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__50284),
            .ce(N__25148),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_10_4  (
            .in0(N__25073),
            .in1(N__26000),
            .in2(_gnd_net_),
            .in3(N__24914),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__50284),
            .ce(N__25148),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_10_5  (
            .in0(N__25964),
            .in1(N__25074),
            .in2(_gnd_net_),
            .in3(N__24911),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50284),
            .ce(N__25148),
            .sr(N__49488));
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_7_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_7_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNIG7JF_2_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__24950),
            .in2(_gnd_net_),
            .in3(N__24976),
            .lcout(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_11_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_11_2  (
            .in0(N__31255),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31294),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_7_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_7_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__31389),
            .in2(_gnd_net_),
            .in3(N__31350),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_7_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_7_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_7_11_5  (
            .in0(N__33870),
            .in1(N__33900),
            .in2(_gnd_net_),
            .in3(N__34742),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_7_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_7_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_7_11_7  (
            .in0(N__31390),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31351),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_12_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_12_0  (
            .in0(N__24945),
            .in1(N__26218),
            .in2(N__24977),
            .in3(N__25275),
            .lcout(\phase_controller_inst2.start_timer_tr_RNO_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26408),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_7_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_7_12_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__31595),
            .in2(_gnd_net_),
            .in3(N__27413),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_7_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_7_13_0 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_7_13_0  (
            .in0(N__24974),
            .in1(N__35074),
            .in2(N__31259),
            .in3(N__37661),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50248),
            .ce(),
            .sr(N__49500));
    defparam \phase_controller_inst2.start_timer_tr_LC_7_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_7_13_1 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_7_13_1  (
            .in0(N__46926),
            .in1(N__24983),
            .in2(N__31573),
            .in3(N__25121),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50248),
            .ce(),
            .sr(N__49500));
    defparam \phase_controller_inst2.state_2_LC_7_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_7_13_5 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst2.state_2_LC_7_13_5  (
            .in0(N__25185),
            .in1(N__24949),
            .in2(N__26268),
            .in3(N__24975),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50248),
            .ce(),
            .sr(N__49500));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_7_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_7_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31565),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50248),
            .ce(),
            .sr(N__49500));
    defparam \phase_controller_inst2.state_3_LC_7_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_7_13_7 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \phase_controller_inst2.state_3_LC_7_13_7  (
            .in0(N__25186),
            .in1(N__25120),
            .in2(N__26269),
            .in3(N__33581),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50248),
            .ce(),
            .sr(N__49500));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_7_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_7_14_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_7_14_0  (
            .in0(N__26137),
            .in1(N__26157),
            .in2(N__25241),
            .in3(N__29162),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_7_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_7_14_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_7_14_1  (
            .in0(N__29161),
            .in1(N__26136),
            .in2(N__26159),
            .in3(N__25237),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_7_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_7_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_7_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_27_LC_7_14_3  (
            .in0(N__31178),
            .in1(N__31199),
            .in2(_gnd_net_),
            .in3(N__34815),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50237),
            .ce(N__29768),
            .sr(N__49504));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_7_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_7_14_5 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_7_14_5  (
            .in0(N__25207),
            .in1(N__26100),
            .in2(N__25229),
            .in3(N__26118),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_7_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_7_14_6 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_7_14_6  (
            .in0(N__26119),
            .in1(N__25228),
            .in2(N__26102),
            .in3(N__25208),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__25193),
            .in2(_gnd_net_),
            .in3(N__26264),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_7_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_7_15_2 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__26406),
            .in2(N__26306),
            .in3(N__26330),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_201_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_7_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_7_15_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_7_15_5  (
            .in0(N__31604),
            .in1(N__26446),
            .in2(_gnd_net_),
            .in3(N__31569),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_7_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_7_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(N__26073),
            .in2(_gnd_net_),
            .in3(N__25252),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_1_LC_7_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_7_16_0 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst2.state_1_LC_7_16_0  (
            .in0(N__26207),
            .in1(N__25277),
            .in2(_gnd_net_),
            .in3(N__26425),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50215),
            .ce(),
            .sr(N__49512));
    defparam \phase_controller_inst2.state_0_LC_7_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_7_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_7_16_5 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \phase_controller_inst2.state_0_LC_7_16_5  (
            .in0(N__26075),
            .in1(N__25276),
            .in2(N__26217),
            .in3(N__25253),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50215),
            .ce(),
            .sr(N__49512));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_7_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_7_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_7_16_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_7_16_7  (
            .in0(N__26407),
            .in1(N__26302),
            .in2(_gnd_net_),
            .in3(N__26327),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50215),
            .ce(),
            .sr(N__49512));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_8_5_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_8_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_8_5_3  (
            .in0(N__28966),
            .in1(N__28938),
            .in2(_gnd_net_),
            .in3(N__34709),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_6_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_6_0  (
            .in0(N__29189),
            .in1(N__34019),
            .in2(N__30807),
            .in3(N__32168),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_8_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_8_6_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_8_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25489),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50315),
            .ce(N__26381),
            .sr(N__49454));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_8_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_8_6_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_8_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25468),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50315),
            .ce(N__26381),
            .sr(N__49454));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_8_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_8_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_8_6_6  (
            .in0(N__29190),
            .in1(N__29217),
            .in2(_gnd_net_),
            .in3(N__34581),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_6_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__30800),
            .in2(N__34711),
            .in3(N__30831),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_7_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__25440),
            .in2(N__25490),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__50307),
            .ce(N__26380),
            .sr(N__49461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__25416),
            .in2(N__25469),
            .in3(N__25448),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__50307),
            .ce(N__26380),
            .sr(N__49461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__25392),
            .in2(N__25445),
            .in3(N__25424),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__50307),
            .ce(N__26380),
            .sr(N__49461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__25368),
            .in2(N__25421),
            .in3(N__25400),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__50307),
            .ce(N__26380),
            .sr(N__49461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__25344),
            .in2(N__25397),
            .in3(N__25376),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__50307),
            .ce(N__26380),
            .sr(N__49461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__25320),
            .in2(N__25373),
            .in3(N__25352),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__50307),
            .ce(N__26380),
            .sr(N__49461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__25296),
            .in2(N__25349),
            .in3(N__25328),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__50307),
            .ce(N__26380),
            .sr(N__49461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__25677),
            .in2(N__25325),
            .in3(N__25304),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__50307),
            .ce(N__26380),
            .sr(N__49461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__25653),
            .in2(N__25301),
            .in3(N__25280),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__50298),
            .ce(N__26371),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__25629),
            .in2(N__25682),
            .in3(N__25661),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__50298),
            .ce(N__26371),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__25605),
            .in2(N__25658),
            .in3(N__25637),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__50298),
            .ce(N__26371),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__25581),
            .in2(N__25634),
            .in3(N__25613),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__50298),
            .ce(N__26371),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__25557),
            .in2(N__25610),
            .in3(N__25589),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__50298),
            .ce(N__26371),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__25533),
            .in2(N__25586),
            .in3(N__25565),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__50298),
            .ce(N__26371),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__25509),
            .in2(N__25562),
            .in3(N__25541),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__50298),
            .ce(N__26371),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__25890),
            .in2(N__25538),
            .in3(N__25517),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__50298),
            .ce(N__26371),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__25866),
            .in2(N__25514),
            .in3(N__25493),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__50285),
            .ce(N__26379),
            .sr(N__49476));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__25842),
            .in2(N__25895),
            .in3(N__25874),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__50285),
            .ce(N__26379),
            .sr(N__49476));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__25818),
            .in2(N__25871),
            .in3(N__25850),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__50285),
            .ce(N__26379),
            .sr(N__49476));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__25794),
            .in2(N__25847),
            .in3(N__25826),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__50285),
            .ce(N__26379),
            .sr(N__49476));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__25770),
            .in2(N__25823),
            .in3(N__25802),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__50285),
            .ce(N__26379),
            .sr(N__49476));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__25746),
            .in2(N__25799),
            .in3(N__25778),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__50285),
            .ce(N__26379),
            .sr(N__49476));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__25722),
            .in2(N__25775),
            .in3(N__25754),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__50285),
            .ce(N__26379),
            .sr(N__49476));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__25698),
            .in2(N__25751),
            .in3(N__25730),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__50285),
            .ce(N__26379),
            .sr(N__49476));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__25983),
            .in2(N__25727),
            .in3(N__25706),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__50272),
            .ce(N__26372),
            .sr(N__49483));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__25947),
            .in2(N__25703),
            .in3(N__26003),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__50272),
            .ce(N__26372),
            .sr(N__49483));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__25999),
            .in2(N__25988),
            .in3(N__25967),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__50272),
            .ce(N__26372),
            .sr(N__49483));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__25963),
            .in2(N__25952),
            .in3(N__25931),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__50272),
            .ce(N__26372),
            .sr(N__49483));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25928),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(N__26372),
            .sr(N__49483));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_8_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__31331),
            .in2(N__25925),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_8_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_8_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_8_11_1  (
            .in0(N__31523),
            .in1(N__26852),
            .in2(_gnd_net_),
            .in3(N__25916),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__50261),
            .ce(),
            .sr(N__49489));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_8_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_8_11_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_8_11_2  (
            .in0(N__31527),
            .in1(N__26831),
            .in2(N__25913),
            .in3(N__25904),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__50261),
            .ce(),
            .sr(N__49489));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_8_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_8_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_8_11_3  (
            .in0(N__31524),
            .in1(N__26810),
            .in2(_gnd_net_),
            .in3(N__25901),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__50261),
            .ce(),
            .sr(N__49489));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_8_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_8_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_8_11_4  (
            .in0(N__31528),
            .in1(N__26777),
            .in2(_gnd_net_),
            .in3(N__25898),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__50261),
            .ce(),
            .sr(N__49489));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_8_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_8_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_8_11_5  (
            .in0(N__31525),
            .in1(N__26756),
            .in2(_gnd_net_),
            .in3(N__26030),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__50261),
            .ce(),
            .sr(N__49489));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_8_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_8_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_8_11_6  (
            .in0(N__31529),
            .in1(N__27128),
            .in2(_gnd_net_),
            .in3(N__26027),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__50261),
            .ce(),
            .sr(N__49489));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_8_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_8_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_8_11_7  (
            .in0(N__31526),
            .in1(N__27107),
            .in2(_gnd_net_),
            .in3(N__26024),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__50261),
            .ce(),
            .sr(N__49489));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_8_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_8_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_8_12_0  (
            .in0(N__31515),
            .in1(N__27089),
            .in2(_gnd_net_),
            .in3(N__26021),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__50249),
            .ce(),
            .sr(N__49493));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_8_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_8_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_8_12_1  (
            .in0(N__31508),
            .in1(N__27058),
            .in2(_gnd_net_),
            .in3(N__26018),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__50249),
            .ce(),
            .sr(N__49493));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_8_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_8_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_8_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_8_12_2  (
            .in0(N__31512),
            .in1(N__27026),
            .in2(_gnd_net_),
            .in3(N__26015),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__50249),
            .ce(),
            .sr(N__49493));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_8_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_8_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_8_12_3  (
            .in0(N__31509),
            .in1(N__26993),
            .in2(_gnd_net_),
            .in3(N__26012),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__50249),
            .ce(),
            .sr(N__49493));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_8_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_8_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_8_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_8_12_4  (
            .in0(N__31513),
            .in1(N__26975),
            .in2(_gnd_net_),
            .in3(N__26009),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__50249),
            .ce(),
            .sr(N__49493));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_8_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_8_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_8_12_5  (
            .in0(N__31510),
            .in1(N__26942),
            .in2(_gnd_net_),
            .in3(N__26006),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__50249),
            .ce(),
            .sr(N__49493));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_8_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_8_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_8_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_8_12_6  (
            .in0(N__31514),
            .in1(N__27248),
            .in2(_gnd_net_),
            .in3(N__26057),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__50249),
            .ce(),
            .sr(N__49493));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_8_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_8_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_8_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_8_12_7  (
            .in0(N__31511),
            .in1(N__29863),
            .in2(_gnd_net_),
            .in3(N__26054),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__50249),
            .ce(),
            .sr(N__49493));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_8_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_8_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_8_13_0  (
            .in0(N__31519),
            .in1(N__29887),
            .in2(_gnd_net_),
            .in3(N__26051),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__50238),
            .ce(),
            .sr(N__49497));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_8_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_8_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_8_13_1  (
            .in0(N__31537),
            .in1(N__29362),
            .in2(_gnd_net_),
            .in3(N__26048),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__50238),
            .ce(),
            .sr(N__49497));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_8_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_8_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_8_13_2  (
            .in0(N__31520),
            .in1(N__29338),
            .in2(_gnd_net_),
            .in3(N__26045),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__50238),
            .ce(),
            .sr(N__49497));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_8_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_8_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_8_13_3  (
            .in0(N__31538),
            .in1(N__29517),
            .in2(_gnd_net_),
            .in3(N__26042),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__50238),
            .ce(),
            .sr(N__49497));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_8_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_8_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_8_13_4  (
            .in0(N__31521),
            .in1(N__29496),
            .in2(_gnd_net_),
            .in3(N__26039),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__50238),
            .ce(),
            .sr(N__49497));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_8_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_8_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_8_13_5  (
            .in0(N__31539),
            .in1(N__26485),
            .in2(_gnd_net_),
            .in3(N__26036),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__50238),
            .ce(),
            .sr(N__49497));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_8_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_8_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_8_13_6  (
            .in0(N__31522),
            .in1(N__26506),
            .in2(_gnd_net_),
            .in3(N__26033),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__50238),
            .ce(),
            .sr(N__49497));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_8_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_8_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_8_13_7  (
            .in0(N__31540),
            .in1(N__26628),
            .in2(_gnd_net_),
            .in3(N__26165),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__50238),
            .ce(),
            .sr(N__49497));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_8_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_8_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_8_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_8_14_0  (
            .in0(N__31530),
            .in1(N__26649),
            .in2(_gnd_net_),
            .in3(N__26162),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__50226),
            .ce(),
            .sr(N__49501));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_8_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_8_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_8_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_8_14_1  (
            .in0(N__31534),
            .in1(N__26158),
            .in2(_gnd_net_),
            .in3(N__26141),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__50226),
            .ce(),
            .sr(N__49501));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_8_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_8_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_8_14_2  (
            .in0(N__31531),
            .in1(N__26138),
            .in2(_gnd_net_),
            .in3(N__26123),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__50226),
            .ce(),
            .sr(N__49501));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_8_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_8_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_8_14_3  (
            .in0(N__31535),
            .in1(N__26120),
            .in2(_gnd_net_),
            .in3(N__26105),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__50226),
            .ce(),
            .sr(N__49501));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_8_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_8_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_8_14_4  (
            .in0(N__31532),
            .in1(N__26101),
            .in2(_gnd_net_),
            .in3(N__26084),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__50226),
            .ce(),
            .sr(N__49501));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_8_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_8_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_8_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_8_14_5  (
            .in0(N__31536),
            .in1(N__26922),
            .in2(_gnd_net_),
            .in3(N__26081),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__50226),
            .ce(),
            .sr(N__49501));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_8_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_8_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_8_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_8_14_6  (
            .in0(N__31533),
            .in1(N__26884),
            .in2(_gnd_net_),
            .in3(N__26078),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50226),
            .ce(),
            .sr(N__49501));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_8_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_8_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_8_15_4 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_8_15_4  (
            .in0(N__26074),
            .in1(N__31380),
            .in2(N__31615),
            .in3(N__27408),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50216),
            .ce(),
            .sr(N__49505));
    defparam \phase_controller_inst2.stoper_tr.running_LC_8_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_8_15_6 .LUT_INIT=16'b1010111000101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_8_15_6  (
            .in0(N__26447),
            .in1(N__31379),
            .in2(N__31616),
            .in3(N__27409),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50216),
            .ce(),
            .sr(N__49505));
    defparam \phase_controller_inst2.start_timer_hc_LC_8_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_8_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_8_15_7 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_8_15_7  (
            .in0(N__26435),
            .in1(N__26429),
            .in2(N__46931),
            .in3(N__31280),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50216),
            .ce(),
            .sr(N__49505));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_8_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_8_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(N__26405),
            .in2(_gnd_net_),
            .in3(N__26298),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_200_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_8_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_8_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_8_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26328),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26282),
            .ce(),
            .sr(N__49513));
    defparam \delay_measurement_inst.stop_timer_tr_LC_8_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_8_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_8_17_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_8_17_5  (
            .in0(N__26329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26282),
            .ce(),
            .sr(N__49513));
    defparam \phase_controller_inst2.S1_LC_8_29_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_8_29_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_8_29_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_8_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26273),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50170),
            .ce(),
            .sr(N__49550));
    defparam \phase_controller_inst2.S2_LC_8_29_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_8_29_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_8_29_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_8_29_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26225),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50170),
            .ce(),
            .sr(N__49550));
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_4.C_ON=1'b0;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_4 (
            .in0(N__50324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clock_output_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_9_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_9_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_9_5_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_23_LC_9_5_4  (
            .in0(N__34710),
            .in1(N__28962),
            .in2(_gnd_net_),
            .in3(N__28946),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50316),
            .ce(N__29758),
            .sr(N__49437));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_9_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_9_6_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_9_6_0  (
            .in0(N__26492),
            .in1(N__26528),
            .in2(N__26519),
            .in3(N__26470),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_9_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_9_6_1 .LUT_INIT=16'b1011001010111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_9_6_1  (
            .in0(N__26527),
            .in1(N__26518),
            .in2(N__26471),
            .in3(N__26491),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_2  (
            .in0(N__34613),
            .in1(N__28618),
            .in2(_gnd_net_),
            .in3(N__28639),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50308),
            .ce(N__29759),
            .sr(N__49447));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_9_6_7  (
            .in0(N__28699),
            .in1(N__28681),
            .in2(_gnd_net_),
            .in3(N__34614),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50308),
            .ce(N__29759),
            .sr(N__49447));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_9_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_9_7_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_9_7_0  (
            .in0(N__29105),
            .in1(N__31164),
            .in2(_gnd_net_),
            .in3(N__26459),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_9_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_9_7_1 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_9_7_1  (
            .in0(N__32253),
            .in1(N__26555),
            .in2(N__26453),
            .in3(N__26564),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_9_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_9_7_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_9_7_2  (
            .in0(N__29025),
            .in1(_gnd_net_),
            .in2(N__26450),
            .in3(N__29005),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_9_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_9_7_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__34364),
            .in2(_gnd_net_),
            .in3(N__34871),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_9_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_9_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_9_7_5  (
            .in0(N__28721),
            .in1(N__28740),
            .in2(_gnd_net_),
            .in3(N__34612),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_9_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_9_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_9_7_6  (
            .in0(N__28818),
            .in1(N__28770),
            .in2(N__28679),
            .in3(N__29578),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_9_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_9_7_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_9_7_7  (
            .in0(N__29441),
            .in1(N__28739),
            .in2(N__26573),
            .in3(N__26570),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_9_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_9_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_9_8_0  (
            .in0(N__28877),
            .in1(N__31104),
            .in2(N__29006),
            .in3(N__33860),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_9_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_9_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_9_8_1  (
            .in0(N__26537),
            .in1(N__26549),
            .in2(N__26558),
            .in3(N__26543),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_9_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_9_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_9_8_2  (
            .in0(N__29270),
            .in1(N__26690),
            .in2(N__33399),
            .in3(N__29631),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_9_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_9_8_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_9_8_3  (
            .in0(N__33022),
            .in1(N__29803),
            .in2(N__33267),
            .in3(N__26722),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_9_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_9_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_9_8_4  (
            .in0(N__28928),
            .in1(N__29678),
            .in2(N__28607),
            .in3(N__34938),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_9_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_9_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_9_8_5  (
            .in0(N__29679),
            .in1(N__29656),
            .in2(_gnd_net_),
            .in3(N__34604),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(elapsed_time_ns_1_RNIV9PBB_0_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_9_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_9_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_9_8_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_21_LC_9_8_6  (
            .in0(N__34605),
            .in1(_gnd_net_),
            .in2(N__26531),
            .in3(N__29680),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50286),
            .ce(N__34321),
            .sr(N__49462));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_9_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_9_9_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_9_9_0  (
            .in0(N__26597),
            .in1(N__32966),
            .in2(N__32993),
            .in3(N__26585),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_9_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_9_1  (
            .in0(N__26691),
            .in1(N__26671),
            .in2(N__34765),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_9_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_9_9_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__34684),
            .in2(N__26600),
            .in3(N__26692),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50273),
            .ce(N__34276),
            .sr(N__49470));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_9_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_9_9_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_9_9_3  (
            .in0(N__34685),
            .in1(N__29308),
            .in2(N__29286),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50273),
            .ce(N__34276),
            .sr(N__49470));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_9_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_9_9_4 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_9_9_4  (
            .in0(N__26596),
            .in1(N__32965),
            .in2(N__32992),
            .in3(N__26584),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_9_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_9_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_9_9_5  (
            .in0(N__34679),
            .in1(N__26734),
            .in2(_gnd_net_),
            .in3(N__26717),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_9_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_9_9_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_9_9_6  (
            .in0(N__26718),
            .in1(_gnd_net_),
            .in2(N__26576),
            .in3(N__34683),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50273),
            .ce(N__34276),
            .sr(N__49470));
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_9_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_9_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_24_LC_9_10_0  (
            .in0(N__34948),
            .in1(N__33830),
            .in2(_gnd_net_),
            .in3(N__34772),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(N__29762),
            .sr(N__49477));
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_9_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_9_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_9_10_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_30_LC_9_10_1  (
            .in0(N__29026),
            .in1(N__34767),
            .in2(_gnd_net_),
            .in3(N__28994),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(N__29762),
            .sr(N__49477));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_9_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_9_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_9_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_9_10_2  (
            .in0(N__28799),
            .in1(N__28782),
            .in2(_gnd_net_),
            .in3(N__34770),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(N__29762),
            .sr(N__49477));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_9_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_9_10_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_9_10_3  (
            .in0(N__34769),
            .in1(N__28748),
            .in2(_gnd_net_),
            .in3(N__28720),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(N__29762),
            .sr(N__49477));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_9_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_9_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_9_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_9_10_4  (
            .in0(N__26735),
            .in1(N__26723),
            .in2(_gnd_net_),
            .in3(N__34771),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(N__29762),
            .sr(N__49477));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_9_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_9_10_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_9_10_5  (
            .in0(N__28829),
            .in1(N__34766),
            .in2(_gnd_net_),
            .in3(N__28844),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(N__29762),
            .sr(N__49477));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_9_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_9_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_9_10_6  (
            .in0(N__34913),
            .in1(N__34885),
            .in2(_gnd_net_),
            .in3(N__34773),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(N__29762),
            .sr(N__49477));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_9_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_9_10_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_9_10_7  (
            .in0(N__34768),
            .in1(N__26696),
            .in2(_gnd_net_),
            .in3(N__26672),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(N__29762),
            .sr(N__49477));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_11_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_11_0  (
            .in0(N__26651),
            .in1(N__26629),
            .in2(N__26612),
            .in3(N__26660),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_9_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_9_11_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_9_11_1  (
            .in0(N__26659),
            .in1(N__26650),
            .in2(N__26633),
            .in3(N__26608),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_9_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_9_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_25_LC_9_11_3  (
            .in0(N__33901),
            .in1(N__33874),
            .in2(_gnd_net_),
            .in3(N__34775),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50250),
            .ce(N__29764),
            .sr(N__49484));
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_11_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_31_LC_9_11_4  (
            .in0(N__34774),
            .in1(N__32243),
            .in2(_gnd_net_),
            .in3(N__32219),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50250),
            .ce(N__29764),
            .sr(N__49484));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_9_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_9_11_5 .LUT_INIT=16'b1101010011011101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_9_11_5  (
            .in0(N__26869),
            .in1(N__26893),
            .in2(N__26906),
            .in3(N__26923),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_9_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_9_11_6 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_9_11_6  (
            .in0(N__26924),
            .in1(N__26905),
            .in2(N__26894),
            .in3(N__26870),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_9_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_9_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__29543),
            .in2(N__26861),
            .in3(N__31327),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_9_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_9_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__29237),
            .in2(N__26840),
            .in3(N__26851),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_9_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_9_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__29174),
            .in2(N__26819),
            .in3(N__26830),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_9_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_9_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__29168),
            .in2(N__26798),
            .in3(N__26809),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_9_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_9_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__26765),
            .in2(N__26789),
            .in3(N__26776),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_9_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_9_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__29399),
            .in2(N__26744),
            .in3(N__26755),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_9_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_9_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__27137),
            .in2(N__27116),
            .in3(N__27127),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_9_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_9_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__27095),
            .in2(N__29147),
            .in3(N__27106),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_9_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_9_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__27077),
            .in2(N__29552),
            .in3(N__27088),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_9_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_9_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__27071),
            .in2(N__27044),
            .in3(N__27062),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_9_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_9_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__27035),
            .in2(N__27014),
            .in3(N__27025),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_9_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_9_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__26981),
            .in2(N__27005),
            .in3(N__26992),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_9_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_9_13_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_9_13_4  (
            .in0(N__26974),
            .in1(N__29693),
            .in2(N__26963),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_9_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_9_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__26930),
            .in2(N__26954),
            .in3(N__26941),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_9_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_9_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__27236),
            .in2(N__29777),
            .in3(N__27247),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_9_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_9_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__29849),
            .in2(N__29906),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_9_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_9_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__29324),
            .in2(N__29393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_9_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_9_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__29468),
            .in2(N__29537),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_9_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_9_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__27230),
            .in2(N__27221),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_9_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_9_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__27209),
            .in2(N__27200),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_9_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_9_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__27185),
            .in2(N__27176),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_9_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_9_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__27164),
            .in2(N__27152),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_9_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_9_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__27440),
            .in2(N__27431),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_9_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_9_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27416),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_9_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_9_15_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_9_15_0  (
            .in0(N__31748),
            .in1(N__27392),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_9_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_9_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_9_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__31739),
            .in2(_gnd_net_),
            .in3(N__27362),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__50205),
            .ce(),
            .sr(N__49502));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_9_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_9_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_9_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__31727),
            .in2(_gnd_net_),
            .in3(N__27332),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__50205),
            .ce(),
            .sr(N__49502));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_9_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_9_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_9_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__31715),
            .in2(_gnd_net_),
            .in3(N__27302),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__50205),
            .ce(),
            .sr(N__49502));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_9_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_9_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_9_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__31703),
            .in2(_gnd_net_),
            .in3(N__27278),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__50205),
            .ce(),
            .sr(N__49502));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_9_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_9_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_9_15_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31691),
            .in3(N__27251),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__50205),
            .ce(),
            .sr(N__49502));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_9_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_9_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_9_15_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31676),
            .in3(N__27683),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__50205),
            .ce(),
            .sr(N__49502));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_9_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_9_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_9_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31661),
            .in3(N__27653),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__50205),
            .ce(),
            .sr(N__49502));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_9_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_9_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_9_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__31928),
            .in2(_gnd_net_),
            .in3(N__27629),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__50196),
            .ce(),
            .sr(N__49506));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_9_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_9_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_9_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__31910),
            .in2(_gnd_net_),
            .in3(N__27596),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__50196),
            .ce(),
            .sr(N__49506));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_9_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_9_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_9_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__31889),
            .in2(_gnd_net_),
            .in3(N__27560),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__50196),
            .ce(),
            .sr(N__49506));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_9_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_9_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_9_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__31874),
            .in2(_gnd_net_),
            .in3(N__27530),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__50196),
            .ce(),
            .sr(N__49506));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_9_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_9_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_9_16_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31862),
            .in3(N__27500),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__50196),
            .ce(),
            .sr(N__49506));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_9_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_9_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_9_16_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31847),
            .in3(N__27473),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__50196),
            .ce(),
            .sr(N__49506));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_9_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_9_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_9_16_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31832),
            .in3(N__27443),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .clk(N__50196),
            .ce(),
            .sr(N__49506));
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_9_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_9_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_9_16_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_15_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31817),
            .in3(N__27932),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .clk(N__50196),
            .ce(),
            .sr(N__49506));
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_9_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_9_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_9_17_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_16_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32048),
            .in3(N__27902),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_16 ),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .clk(N__50190),
            .ce(),
            .sr(N__49508));
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_9_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_9_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_9_17_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_17_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32033),
            .in3(N__27866),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .clk(N__50190),
            .ce(),
            .sr(N__49508));
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_9_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_9_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_9_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_18_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__32018),
            .in2(_gnd_net_),
            .in3(N__27836),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .clk(N__50190),
            .ce(),
            .sr(N__49508));
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_9_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_9_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_9_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_19_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__31997),
            .in2(_gnd_net_),
            .in3(N__27803),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .clk(N__50190),
            .ce(),
            .sr(N__49508));
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_9_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_9_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_9_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_20_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__31985),
            .in2(_gnd_net_),
            .in3(N__27767),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .clk(N__50190),
            .ce(),
            .sr(N__49508));
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_9_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_9_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_9_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_21_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__31973),
            .in2(_gnd_net_),
            .in3(N__27740),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .clk(N__50190),
            .ce(),
            .sr(N__49508));
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_9_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_9_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_9_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_22_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(N__31961),
            .in2(_gnd_net_),
            .in3(N__27707),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .clk(N__50190),
            .ce(),
            .sr(N__49508));
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_9_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_9_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_9_17_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_23_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31949),
            .in3(N__28178),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .clk(N__50190),
            .ce(),
            .sr(N__49508));
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_9_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_9_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_9_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_24_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__32150),
            .in2(_gnd_net_),
            .in3(N__28145),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_24 ),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .clk(N__50186),
            .ce(),
            .sr(N__49514));
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_9_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_9_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_9_18_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_25_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32138),
            .in3(N__28118),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .clk(N__50186),
            .ce(),
            .sr(N__49514));
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_9_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_9_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_9_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_26_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__32123),
            .in2(_gnd_net_),
            .in3(N__28085),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .clk(N__50186),
            .ce(),
            .sr(N__49514));
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_9_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_9_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_9_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_27_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__32111),
            .in2(_gnd_net_),
            .in3(N__28058),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .clk(N__50186),
            .ce(),
            .sr(N__49514));
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_9_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_9_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_9_18_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_28_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32099),
            .in3(N__28028),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .clk(N__50186),
            .ce(),
            .sr(N__49514));
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_9_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_9_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_9_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_29_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__32084),
            .in2(_gnd_net_),
            .in3(N__28001),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .clk(N__50186),
            .ce(),
            .sr(N__49514));
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_9_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_9_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_9_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_30_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__30107),
            .in2(_gnd_net_),
            .in3(N__27965),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ),
            .clk(N__50186),
            .ce(),
            .sr(N__49514));
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_9_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_9_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_9_18_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_31_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__32069),
            .in2(_gnd_net_),
            .in3(N__28490),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50186),
            .ce(),
            .sr(N__49514));
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_9_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_9_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_9_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_31_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28487),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50181),
            .ce(),
            .sr(N__49521));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_9_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_9_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_9_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28466),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50174),
            .ce(),
            .sr(N__49533));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_9_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_9_26_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_9_26_0  (
            .in0(_gnd_net_),
            .in1(N__28403),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_26_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_9_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_9_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_9_26_1  (
            .in0(_gnd_net_),
            .in1(N__28379),
            .in2(_gnd_net_),
            .in3(N__28337),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_9_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_9_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_9_26_2  (
            .in0(_gnd_net_),
            .in1(N__28334),
            .in2(_gnd_net_),
            .in3(N__28298),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_9_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_9_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_9_26_3  (
            .in0(_gnd_net_),
            .in1(N__28295),
            .in2(_gnd_net_),
            .in3(N__28259),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_9_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_9_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_9_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_9_26_4  (
            .in0(_gnd_net_),
            .in1(N__30062),
            .in2(_gnd_net_),
            .in3(N__28235),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_9_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_9_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_9_26_5  (
            .in0(_gnd_net_),
            .in1(N__48431),
            .in2(N__30017),
            .in3(N__28211),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_9_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_9_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_9_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_9_26_6  (
            .in0(_gnd_net_),
            .in1(N__29966),
            .in2(N__48440),
            .in3(N__28538),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_9_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_9_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_9_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_9_26_7  (
            .in0(_gnd_net_),
            .in1(N__48435),
            .in2(N__29921),
            .in3(N__28511),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_9_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_9_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_9_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_9_27_0  (
            .in0(_gnd_net_),
            .in1(N__30374),
            .in2(_gnd_net_),
            .in3(N__28493),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_9_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_9_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_9_27_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_9_27_1  (
            .in0(_gnd_net_),
            .in1(N__30329),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_9_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_9_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_9_27_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_9_27_2  (
            .in0(_gnd_net_),
            .in1(N__30284),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_9_27_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_9_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_9_27_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_9_27_3  (
            .in0(_gnd_net_),
            .in1(N__30242),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_9_27_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_9_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_9_27_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_9_27_4  (
            .in0(_gnd_net_),
            .in1(N__30197),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_9_27_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_9_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_9_27_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_9_27_5  (
            .in0(_gnd_net_),
            .in1(N__30146),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_9_27_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_9_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_9_27_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_9_27_6  (
            .in0(_gnd_net_),
            .in1(N__30116),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_9_27_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_9_27_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_9_27_7  (
            .in0(_gnd_net_),
            .in1(N__30659),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_9_28_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_9_28_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_9_28_0  (
            .in0(_gnd_net_),
            .in1(N__30629),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_28_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_9_28_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_9_28_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_9_28_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_9_28_1  (
            .in0(_gnd_net_),
            .in1(N__30599),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_9_28_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_9_28_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_9_28_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_9_28_2  (
            .in0(_gnd_net_),
            .in1(N__30569),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_9_28_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_9_28_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_9_28_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_9_28_3  (
            .in0(_gnd_net_),
            .in1(N__30548),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_9_28_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_9_28_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_9_28_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_9_28_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28580),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_4_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_4_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_10_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28565),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50309),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_4_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_4_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_10_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28577),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50309),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_6_0  (
            .in0(N__28640),
            .in1(N__28617),
            .in2(_gnd_net_),
            .in3(N__34603),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_6_2  (
            .in0(N__28906),
            .in1(N__28885),
            .in2(_gnd_net_),
            .in3(N__34601),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_6_3  (
            .in0(N__34599),
            .in1(N__29307),
            .in2(_gnd_net_),
            .in3(N__29287),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_6_4  (
            .in0(N__29419),
            .in1(N__29458),
            .in2(_gnd_net_),
            .in3(N__34600),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_10_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_10_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_10_6_6  (
            .in0(N__28700),
            .in1(N__28680),
            .in2(_gnd_net_),
            .in3(N__34602),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_10_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_10_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_10_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_10_7_0  (
            .in0(N__29454),
            .in1(N__29415),
            .in2(_gnd_net_),
            .in3(N__34672),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(N__34312),
            .sr(N__49438));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_10_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_10_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_10_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_10_7_1  (
            .in0(N__34669),
            .in1(N__28747),
            .in2(_gnd_net_),
            .in3(N__28719),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(N__34312),
            .sr(N__49438));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_10_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_10_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_10_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_10_7_2  (
            .in0(N__28698),
            .in1(N__28682),
            .in2(_gnd_net_),
            .in3(N__34670),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(N__34312),
            .sr(N__49438));
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_10_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_10_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_10_7_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_22_LC_10_7_3  (
            .in0(N__34666),
            .in1(N__28638),
            .in2(N__28622),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(N__34312),
            .sr(N__49438));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_10_7_5  (
            .in0(N__34668),
            .in1(N__29224),
            .in2(_gnd_net_),
            .in3(N__29197),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(N__34312),
            .sr(N__49438));
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_10_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_10_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_10_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_23_LC_10_7_6  (
            .in0(N__28970),
            .in1(N__28945),
            .in2(_gnd_net_),
            .in3(N__34671),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(N__34312),
            .sr(N__49438));
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_10_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_10_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_10_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_29_LC_10_7_7  (
            .in0(N__34667),
            .in1(N__28902),
            .in2(_gnd_net_),
            .in3(N__28884),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(N__34312),
            .sr(N__49438));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_8_0  (
            .in0(N__34608),
            .in1(N__28827),
            .in2(_gnd_net_),
            .in3(N__28840),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(elapsed_time_ns_1_RNIU7OBB_0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_10_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_10_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_10_8_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_10_8_1  (
            .in0(N__28828),
            .in1(_gnd_net_),
            .in2(N__28802),
            .in3(N__34611),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50263),
            .ce(N__34316),
            .sr(N__49448));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_10_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_10_8_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_10_8_2  (
            .in0(N__34606),
            .in1(N__28783),
            .in2(_gnd_net_),
            .in3(N__28795),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_10_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_10_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_10_8_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_10_8_3  (
            .in0(N__28784),
            .in1(_gnd_net_),
            .in2(N__28754),
            .in3(N__34610),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50263),
            .ce(N__34316),
            .sr(N__49448));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_8_5  (
            .in0(N__29592),
            .in1(N__29563),
            .in2(_gnd_net_),
            .in3(N__34607),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(elapsed_time_ns_1_RNILK91B_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_10_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_10_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_10_8_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_10_8_6  (
            .in0(N__34609),
            .in1(_gnd_net_),
            .in2(N__28751),
            .in3(N__29593),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50263),
            .ce(N__34316),
            .sr(N__49448));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_9_0 .LUT_INIT=16'b0101000011010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_9_0  (
            .in0(N__32920),
            .in1(N__29132),
            .in2(N__29123),
            .in3(N__32944),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_9_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_9_1  (
            .in0(N__29640),
            .in1(N__29611),
            .in2(_gnd_net_),
            .in3(N__34733),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_10_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_10_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_10_9_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_20_LC_10_9_2  (
            .in0(N__34735),
            .in1(_gnd_net_),
            .in2(N__29138),
            .in3(N__29641),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50252),
            .ce(N__34263),
            .sr(N__49455));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_10_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_10_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_10_9_3  (
            .in0(N__29817),
            .in1(N__29788),
            .in2(_gnd_net_),
            .in3(N__34732),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(elapsed_time_ns_1_RNI2COBB_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_10_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_10_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_10_9_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_10_9_4  (
            .in0(N__34734),
            .in1(_gnd_net_),
            .in2(N__29135),
            .in3(N__29818),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50252),
            .ce(N__34263),
            .sr(N__49455));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_10_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_10_9_5 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_10_9_5  (
            .in0(N__29131),
            .in1(N__32921),
            .in2(N__32945),
            .in3(N__29122),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_10_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_10_0  (
            .in0(N__29054),
            .in1(N__33134),
            .in2(N__29045),
            .in3(N__33155),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_28_LC_10_10_2  (
            .in0(N__29107),
            .in1(N__29075),
            .in2(_gnd_net_),
            .in3(N__34839),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50240),
            .ce(N__34254),
            .sr(N__49463));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_10_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_10_4  (
            .in0(N__29053),
            .in1(N__33133),
            .in2(N__29044),
            .in3(N__33154),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_10_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_10_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_10_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_30_LC_10_10_6  (
            .in0(N__29027),
            .in1(N__29001),
            .in2(_gnd_net_),
            .in3(N__34840),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50240),
            .ce(N__34254),
            .sr(N__49463));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_10_7 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_10_7  (
            .in0(N__31646),
            .in1(N__33112),
            .in2(N__33083),
            .in3(N__31634),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_11_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_11_0  (
            .in0(N__29368),
            .in1(N__29347),
            .in2(N__29249),
            .in3(N__29378),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_10_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_10_11_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_10_11_1  (
            .in0(N__29377),
            .in1(N__29369),
            .in2(N__29348),
            .in3(N__29245),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_10_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_10_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_10_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_10_11_3  (
            .in0(N__29312),
            .in1(N__29288),
            .in2(_gnd_net_),
            .in3(N__34830),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50228),
            .ce(N__29761),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_10_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_10_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_10_11_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_10_11_4  (
            .in0(N__34828),
            .in1(N__34001),
            .in2(_gnd_net_),
            .in3(N__34043),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50228),
            .ce(N__29761),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_10_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_10_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_10_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_10_11_5  (
            .in0(N__29231),
            .in1(N__29201),
            .in2(_gnd_net_),
            .in3(N__34831),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50228),
            .ce(N__29761),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_10_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_10_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_10_11_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_10_11_6  (
            .in0(N__34829),
            .in1(N__30845),
            .in2(_gnd_net_),
            .in3(N__30814),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50228),
            .ce(N__29761),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_10_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_10_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_10_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_26_LC_10_12_0  (
            .in0(N__34833),
            .in1(N__31121),
            .in2(_gnd_net_),
            .in3(N__31136),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(N__29763),
            .sr(N__49478));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_10_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_10_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_10_12_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_10_12_1  (
            .in0(N__34412),
            .in1(N__34838),
            .in2(_gnd_net_),
            .in3(N__34384),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(N__29763),
            .sr(N__49478));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_12_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_10_12_3  (
            .in0(N__33041),
            .in1(N__34835),
            .in2(_gnd_net_),
            .in3(N__33059),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(N__29763),
            .sr(N__49478));
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_10_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_10_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_10_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_21_LC_10_12_4  (
            .in0(N__34832),
            .in1(N__29687),
            .in2(_gnd_net_),
            .in3(N__29663),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(N__29763),
            .sr(N__49478));
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_10_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_10_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_10_12_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_20_LC_10_12_5  (
            .in0(N__29645),
            .in1(N__34837),
            .in2(_gnd_net_),
            .in3(N__29615),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(N__29763),
            .sr(N__49478));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_10_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_10_12_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_10_12_6  (
            .in0(N__34834),
            .in1(N__29600),
            .in2(_gnd_net_),
            .in3(N__29567),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(N__29763),
            .sr(N__49478));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_10_12_7  (
            .in0(N__32744),
            .in1(N__34836),
            .in2(_gnd_net_),
            .in3(N__32186),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(N__29763),
            .sr(N__49478));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_13_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_13_0  (
            .in0(N__29518),
            .in1(N__29528),
            .in2(N__29480),
            .in3(N__29500),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_10_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_10_13_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_10_13_1  (
            .in0(N__29527),
            .in1(N__29519),
            .in2(N__29501),
            .in3(N__29479),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_10_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_10_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_10_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_10_13_4  (
            .in0(N__29462),
            .in1(N__29423),
            .in2(_gnd_net_),
            .in3(N__34844),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50207),
            .ce(N__29765),
            .sr(N__49485));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_14_0 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_14_0  (
            .in0(N__29843),
            .in1(N__29869),
            .in2(N__29834),
            .in3(N__29894),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_10_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_10_14_1 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_10_14_1  (
            .in0(N__29893),
            .in1(N__29842),
            .in2(N__29873),
            .in3(N__29830),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_10_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_10_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_10_14_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_10_14_2  (
            .in0(N__33281),
            .in1(N__33299),
            .in2(_gnd_net_),
            .in3(N__34843),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50197),
            .ce(N__29766),
            .sr(N__49490));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_10_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_10_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_10_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_10_14_3  (
            .in0(N__34841),
            .in1(N__33412),
            .in2(_gnd_net_),
            .in3(N__33434),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50197),
            .ce(N__29766),
            .sr(N__49490));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_10_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_10_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_10_14_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_10_14_6  (
            .in0(N__29822),
            .in1(N__29792),
            .in2(_gnd_net_),
            .in3(N__34842),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50197),
            .ce(N__29766),
            .sr(N__49490));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_10_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_10_15_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_10_15_0  (
            .in0(N__36464),
            .in1(N__33707),
            .in2(_gnd_net_),
            .in3(N__43574),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_10_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_10_15_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_10_15_2  (
            .in0(N__36386),
            .in1(N__33653),
            .in2(_gnd_net_),
            .in3(N__43572),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(\current_shift_inst.control_input_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_15_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29729),
            .in3(N__31768),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50191),
            .ce(),
            .sr(N__49494));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43573),
            .lcout(\current_shift_inst.N_1269_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_10_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_10_15_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_10_15_7  (
            .in0(N__43575),
            .in1(N__36449),
            .in2(_gnd_net_),
            .in3(N__33692),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_10_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_10_16_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_10_16_0  (
            .in0(N__33677),
            .in1(N__36434),
            .in2(_gnd_net_),
            .in3(N__43591),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_10_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_10_17_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_10_17_0  (
            .in0(N__33746),
            .in1(N__36530),
            .in2(_gnd_net_),
            .in3(N__43592),
            .lcout(\current_shift_inst.control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_10_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_10_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32065),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_10_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_10_23_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_10_23_3  (
            .in0(N__32522),
            .in1(N__32551),
            .in2(_gnd_net_),
            .in3(N__32367),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_10_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_10_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_10_26_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_10_26_0  (
            .in0(_gnd_net_),
            .in1(N__30101),
            .in2(N__30083),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_10_26_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_10_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_10_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_10_26_1  (
            .in0(_gnd_net_),
            .in1(N__30056),
            .in2(N__30038),
            .in3(N__30008),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_10_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_10_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_10_26_2  (
            .in0(_gnd_net_),
            .in1(N__30005),
            .in2(N__29987),
            .in3(N__29960),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_10_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_10_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_10_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_10_26_3  (
            .in0(_gnd_net_),
            .in1(N__29957),
            .in2(N__29942),
            .in3(N__29909),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_10_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_10_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_10_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_10_26_4  (
            .in0(_gnd_net_),
            .in1(N__30413),
            .in2(N__30395),
            .in3(N__30368),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_10_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_10_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_10_26_5  (
            .in0(_gnd_net_),
            .in1(N__30365),
            .in2(N__30347),
            .in3(N__30323),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_10_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_10_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_10_26_6  (
            .in0(_gnd_net_),
            .in1(N__30320),
            .in2(N__30302),
            .in3(N__30278),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_10_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_10_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_10_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_10_26_7  (
            .in0(_gnd_net_),
            .in1(N__30275),
            .in2(N__30260),
            .in3(N__30236),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_10_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_10_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_10_27_0  (
            .in0(_gnd_net_),
            .in1(N__30233),
            .in2(N__30218),
            .in3(N__30191),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(bfn_10_27_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_10_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_10_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_10_27_1  (
            .in0(_gnd_net_),
            .in1(N__30188),
            .in2(N__30170),
            .in3(N__30140),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_10_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_10_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_10_27_2  (
            .in0(_gnd_net_),
            .in1(N__32501),
            .in2(N__30137),
            .in3(N__30110),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_10_27_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_10_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_10_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_10_27_3  (
            .in0(_gnd_net_),
            .in1(N__32504),
            .in2(N__30683),
            .in3(N__30653),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_10_27_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_10_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_10_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_10_27_4  (
            .in0(_gnd_net_),
            .in1(N__32502),
            .in2(N__30650),
            .in3(N__30623),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_10_27_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_10_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_10_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_10_27_5  (
            .in0(_gnd_net_),
            .in1(N__32505),
            .in2(N__30620),
            .in3(N__30593),
            .lcout(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_10_27_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_10_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_10_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_10_27_6  (
            .in0(_gnd_net_),
            .in1(N__32503),
            .in2(N__30590),
            .in3(N__30563),
            .lcout(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_10_27_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_10_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_10_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_10_27_7  (
            .in0(_gnd_net_),
            .in1(N__32506),
            .in2(N__30560),
            .in3(N__30542),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_10_28_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_10_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_10_28_0  (
            .in0(N__30539),
            .in1(N__32291),
            .in2(_gnd_net_),
            .in3(N__30533),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_11_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_11_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_11_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_11_5_4  (
            .in0(N__33997),
            .in1(N__34738),
            .in2(_gnd_net_),
            .in3(N__34039),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50288),
            .ce(N__34337),
            .sr(N__49413));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_11_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_11_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_11_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_11_6_6  (
            .in0(N__34757),
            .in1(N__32733),
            .in2(_gnd_net_),
            .in3(N__32179),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50275),
            .ce(N__34280),
            .sr(N__49418));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_11_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_11_7_0 .LUT_INIT=16'b0111010100010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_11_7_0  (
            .in0(N__32879),
            .in1(N__32900),
            .in2(N__30868),
            .in3(N__30854),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_11_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_11_7_4 .LUT_INIT=16'b1111011101010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_11_7_4  (
            .in0(N__32878),
            .in1(N__32899),
            .in2(N__30869),
            .in3(N__30853),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_11_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_11_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_11_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_11_7_7  (
            .in0(N__30838),
            .in1(N__30815),
            .in2(_gnd_net_),
            .in3(N__34673),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50264),
            .ce(N__34322),
            .sr(N__49427));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__30770),
            .in2(N__30782),
            .in3(N__32713),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__30764),
            .in2(N__30755),
            .in3(N__32680),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__30746),
            .in2(N__30740),
            .in3(N__32662),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_8_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_8_3  (
            .in0(N__32647),
            .in1(N__30722),
            .in2(N__30731),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__30716),
            .in2(N__30710),
            .in3(N__32632),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_8_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_8_5  (
            .in0(N__32617),
            .in1(N__30701),
            .in2(N__30695),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__34853),
            .in2(N__30980),
            .in3(N__32602),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__34346),
            .in2(N__30971),
            .in3(N__32587),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__30962),
            .in2(N__30956),
            .in3(N__32851),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__30947),
            .in2(N__30941),
            .in3(N__32836),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__30932),
            .in2(N__30926),
            .in3(N__32821),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_9_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_9_3  (
            .in0(N__32806),
            .in1(N__30914),
            .in2(N__30905),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__30893),
            .in2(N__33008),
            .in3(N__32791),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_9_5  (
            .in0(N__32776),
            .in1(N__30887),
            .in2(N__30878),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_9_6  (
            .in0(N__32761),
            .in1(N__31070),
            .in2(N__31079),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__33308),
            .in2(N__33374),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__31064),
            .in2(N__31052),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__31034),
            .in2(N__31028),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__31019),
            .in2(N__31010),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__33920),
            .in2(N__33971),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__31205),
            .in2(N__31214),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__30998),
            .in2(N__30992),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_11_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_11_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__31622),
            .in2(N__31226),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_11_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_11_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31217),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_11_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_11_11_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_11_11_0  (
            .in0(N__31145),
            .in1(N__31088),
            .in2(N__33197),
            .in3(N__33174),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_11_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_11_11_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_11_11_1  (
            .in0(N__31087),
            .in1(N__33195),
            .in2(N__33176),
            .in3(N__31144),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_11_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_11_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_11_11_2  (
            .in0(N__31173),
            .in1(N__31192),
            .in2(_gnd_net_),
            .in3(N__34746),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_11_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_11_11_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_27_LC_11_11_3  (
            .in0(N__34749),
            .in1(_gnd_net_),
            .in2(N__31181),
            .in3(N__31174),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50219),
            .ce(N__34261),
            .sr(N__49464));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_11_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_11_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_11_11_4  (
            .in0(N__31119),
            .in1(N__31135),
            .in2(_gnd_net_),
            .in3(N__34747),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_11_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_11_11_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_26_LC_11_11_5  (
            .in0(N__34748),
            .in1(_gnd_net_),
            .in2(N__31124),
            .in3(N__31120),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50219),
            .ce(N__34261),
            .sr(N__49464));
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_11_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_11_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_31_LC_11_11_6  (
            .in0(N__32257),
            .in1(N__32215),
            .in2(_gnd_net_),
            .in3(N__34750),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50219),
            .ce(N__34261),
            .sr(N__49464));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_11_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_11_11_7 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_11_11_7  (
            .in0(N__31645),
            .in1(N__33078),
            .in2(N__33113),
            .in3(N__31633),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_11_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_11_12_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__31614),
            .in2(_gnd_net_),
            .in3(N__31574),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_11_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_11_12_3 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_11_12_3  (
            .in0(N__31391),
            .in1(N__31355),
            .in2(N__31334),
            .in3(N__31326),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50208),
            .ce(),
            .sr(N__49472));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_11_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_11_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_11_13_0 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_11_13_0  (
            .in0(N__34141),
            .in1(N__33226),
            .in2(N__35171),
            .in3(N__32712),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50198),
            .ce(),
            .sr(N__49479));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_13_3 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_13_3  (
            .in0(N__31242),
            .in1(N__31303),
            .in2(_gnd_net_),
            .in3(N__31290),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_13_4 .LUT_INIT=16'b1011101000111010;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_11_13_4  (
            .in0(N__31304),
            .in1(N__31243),
            .in2(N__31307),
            .in3(N__37657),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50198),
            .ce(),
            .sr(N__49479));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_11_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_11_13_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__31241),
            .in2(_gnd_net_),
            .in3(N__37656),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_11_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_11_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_11_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31295),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50192),
            .ce(),
            .sr(N__49486));
    defparam \phase_controller_inst1.T45_LC_11_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.T45_LC_11_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T45_LC_11_14_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.T45_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__31786),
            .in2(_gnd_net_),
            .in3(N__33457),
            .lcout(T45_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50192),
            .ce(),
            .sr(N__49486));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_11_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_11_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__31775),
            .in2(N__31769),
            .in3(N__31767),
            .lcout(\current_shift_inst.control_input_1 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_11_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_11_15_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__33506),
            .in2(_gnd_net_),
            .in3(N__31730),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__33500),
            .in2(_gnd_net_),
            .in3(N__31718),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_15_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__33494),
            .in2(_gnd_net_),
            .in3(N__31706),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_15_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__33488),
            .in2(_gnd_net_),
            .in3(N__31694),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_11_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_11_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__33482),
            .in2(_gnd_net_),
            .in3(N__31679),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_15_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__33476),
            .in2(_gnd_net_),
            .in3(N__31664),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_15_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__35201),
            .in2(_gnd_net_),
            .in3(N__31649),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_11_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_11_16_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__31934),
            .in2(_gnd_net_),
            .in3(N__31919),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_16_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__31916),
            .in2(_gnd_net_),
            .in3(N__31901),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_16_2 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31898),
            .in3(N__31877),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_16_3 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35339),
            .in3(N__31865),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_11_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_11_16_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__35321),
            .in2(_gnd_net_),
            .in3(N__31850),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_11_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_11_16_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__35303),
            .in2(_gnd_net_),
            .in3(N__31835),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_12 ),
            .carryout(\current_shift_inst.control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_11_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_11_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__35285),
            .in2(_gnd_net_),
            .in3(N__31820),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_13 ),
            .carryout(\current_shift_inst.control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_11_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_11_16_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__35267),
            .in2(_gnd_net_),
            .in3(N__31805),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_14 ),
            .carryout(\current_shift_inst.control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_11_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_11_17_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__35393),
            .in2(_gnd_net_),
            .in3(N__32036),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\current_shift_inst.control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_11_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_11_17_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__32564),
            .in2(_gnd_net_),
            .in3(N__32021),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_16 ),
            .carryout(\current_shift_inst.control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_11_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_11_17_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__32573),
            .in2(_gnd_net_),
            .in3(N__32006),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_17 ),
            .carryout(\current_shift_inst.control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_11_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_11_17_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__32003),
            .in2(_gnd_net_),
            .in3(N__31988),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_18 ),
            .carryout(\current_shift_inst.control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_11_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_11_17_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__35462),
            .in2(_gnd_net_),
            .in3(N__31976),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_19 ),
            .carryout(\current_shift_inst.control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_11_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_11_17_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__35747),
            .in2(_gnd_net_),
            .in3(N__31964),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_20 ),
            .carryout(\current_shift_inst.control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_17_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__35729),
            .in2(_gnd_net_),
            .in3(N__31952),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_21 ),
            .carryout(\current_shift_inst.control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_11_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_11_17_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__35702),
            .in2(_gnd_net_),
            .in3(N__31937),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_22 ),
            .carryout(\current_shift_inst.control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_11_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_11_18_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__35534),
            .in2(_gnd_net_),
            .in3(N__32141),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\current_shift_inst.control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_11_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_11_18_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__35378),
            .in2(_gnd_net_),
            .in3(N__32126),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_24 ),
            .carryout(\current_shift_inst.control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_11_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_11_18_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__35480),
            .in2(_gnd_net_),
            .in3(N__32114),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_25 ),
            .carryout(\current_shift_inst.control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_11_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_11_18_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__32054),
            .in2(_gnd_net_),
            .in3(N__32102),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_26 ),
            .carryout(\current_shift_inst.control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_11_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_11_18_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__33788),
            .in2(_gnd_net_),
            .in3(N__32087),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_27 ),
            .carryout(\current_shift_inst.control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_11_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_11_18_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__33782),
            .in2(_gnd_net_),
            .in3(N__32075),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_28 ),
            .carryout(\current_shift_inst.control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_11_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_11_18_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_11_18_6  (
            .in0(N__43516),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32072),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_11_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_11_18_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_11_18_7  (
            .in0(N__36638),
            .in1(N__33800),
            .in2(_gnd_net_),
            .in3(N__43515),
            .lcout(\current_shift_inst.control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_11_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_11_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_11_19_0  (
            .in0(N__45376),
            .in1(N__41055),
            .in2(N__42785),
            .in3(N__41017),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_11_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_11_19_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_11_19_5  (
            .in0(N__43560),
            .in1(N__33755),
            .in2(_gnd_net_),
            .in3(N__36554),
            .lcout(\current_shift_inst.control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_19_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_19_6  (
            .in0(N__33764),
            .in1(N__36569),
            .in2(_gnd_net_),
            .in3(N__43559),
            .lcout(\current_shift_inst.control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_11_23_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_11_23_0 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_11_23_0  (
            .in0(N__32555),
            .in1(N__32521),
            .in2(N__32411),
            .in3(N__32309),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_4_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_4_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_12_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32264),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50287),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_12_4_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_12_4_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_12_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_12_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32279),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50287),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_12_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_5_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35852),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34054),
            .ce(),
            .sr(N__49405));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_6_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__35170),
            .in2(_gnd_net_),
            .in3(N__33230),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_12_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_12_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_12_6_3  (
            .in0(N__32258),
            .in1(N__32208),
            .in2(_gnd_net_),
            .in3(N__34737),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_12_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_12_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_12_6_7  (
            .in0(N__32178),
            .in1(N__32737),
            .in2(_gnd_net_),
            .in3(N__34736),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_12_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_12_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__32717),
            .in2(N__32690),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_12_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_12_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_12_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_12_7_1  (
            .in0(N__34234),
            .in1(N__32681),
            .in2(_gnd_net_),
            .in3(N__32669),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__50251),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_12_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_12_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_12_7_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_12_7_2  (
            .in0(N__34331),
            .in1(N__33209),
            .in2(N__32666),
            .in3(N__32651),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__50251),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_12_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_12_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_12_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_12_7_3  (
            .in0(N__34235),
            .in1(N__32648),
            .in2(_gnd_net_),
            .in3(N__32636),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__50251),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_12_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_12_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_12_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_12_7_4  (
            .in0(N__34332),
            .in1(N__32633),
            .in2(_gnd_net_),
            .in3(N__32621),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__50251),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_12_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_12_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_12_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_12_7_5  (
            .in0(N__34236),
            .in1(N__32618),
            .in2(_gnd_net_),
            .in3(N__32606),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__50251),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_12_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_12_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_12_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_12_7_6  (
            .in0(N__34333),
            .in1(N__32603),
            .in2(_gnd_net_),
            .in3(N__32591),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__50251),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_7_7  (
            .in0(N__34237),
            .in1(N__32588),
            .in2(_gnd_net_),
            .in3(N__32576),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__50251),
            .ce(),
            .sr(N__49419));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_8_0  (
            .in0(N__34330),
            .in1(N__32852),
            .in2(_gnd_net_),
            .in3(N__32840),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__50239),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_12_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_12_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_12_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_12_8_1  (
            .in0(N__34317),
            .in1(N__32837),
            .in2(_gnd_net_),
            .in3(N__32825),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__50239),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_12_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_12_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_12_8_2  (
            .in0(N__34327),
            .in1(N__32822),
            .in2(_gnd_net_),
            .in3(N__32810),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__50239),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_12_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_12_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_12_8_3  (
            .in0(N__34318),
            .in1(N__32807),
            .in2(_gnd_net_),
            .in3(N__32795),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__50239),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_12_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_12_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_12_8_4  (
            .in0(N__34328),
            .in1(N__32792),
            .in2(_gnd_net_),
            .in3(N__32780),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__50239),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_12_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_12_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_12_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_12_8_5  (
            .in0(N__34319),
            .in1(N__32777),
            .in2(_gnd_net_),
            .in3(N__32765),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__50239),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_12_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_12_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_12_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_12_8_6  (
            .in0(N__34329),
            .in1(N__32762),
            .in2(_gnd_net_),
            .in3(N__32750),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__50239),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_12_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_12_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_12_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_12_8_7  (
            .in0(N__34320),
            .in1(N__33354),
            .in2(_gnd_net_),
            .in3(N__32747),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__50239),
            .ce(),
            .sr(N__49428));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_12_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_12_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_12_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_12_9_0  (
            .in0(N__34230),
            .in1(N__33324),
            .in2(_gnd_net_),
            .in3(N__32996),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__50227),
            .ce(),
            .sr(N__49439));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_12_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_12_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_12_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_12_9_1  (
            .in0(N__34323),
            .in1(N__32985),
            .in2(_gnd_net_),
            .in3(N__32969),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__50227),
            .ce(),
            .sr(N__49439));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_12_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_12_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_12_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_12_9_2  (
            .in0(N__34231),
            .in1(N__32964),
            .in2(_gnd_net_),
            .in3(N__32948),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__50227),
            .ce(),
            .sr(N__49439));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_12_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_12_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_12_9_3  (
            .in0(N__34324),
            .in1(N__32940),
            .in2(_gnd_net_),
            .in3(N__32924),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__50227),
            .ce(),
            .sr(N__49439));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_12_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_12_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_12_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_12_9_4  (
            .in0(N__34232),
            .in1(N__32919),
            .in2(_gnd_net_),
            .in3(N__32903),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__50227),
            .ce(),
            .sr(N__49439));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_12_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_12_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_12_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_12_9_5  (
            .in0(N__34325),
            .in1(N__32898),
            .in2(_gnd_net_),
            .in3(N__32882),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__50227),
            .ce(),
            .sr(N__49439));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_12_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_12_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_12_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_12_9_6  (
            .in0(N__34233),
            .in1(N__32877),
            .in2(_gnd_net_),
            .in3(N__32861),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__50227),
            .ce(),
            .sr(N__49439));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_12_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_12_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_12_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_12_9_7  (
            .in0(N__34326),
            .in1(N__33956),
            .in2(_gnd_net_),
            .in3(N__32858),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__50227),
            .ce(),
            .sr(N__49439));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_12_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_12_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_12_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_12_10_0  (
            .in0(N__34226),
            .in1(N__33936),
            .in2(_gnd_net_),
            .in3(N__32855),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__50217),
            .ce(),
            .sr(N__49449));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_12_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_12_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_12_10_1  (
            .in0(N__34309),
            .in1(N__33196),
            .in2(_gnd_net_),
            .in3(N__33179),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__50217),
            .ce(),
            .sr(N__49449));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_12_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_12_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_12_10_2  (
            .in0(N__34227),
            .in1(N__33175),
            .in2(_gnd_net_),
            .in3(N__33158),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__50217),
            .ce(),
            .sr(N__49449));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_12_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_12_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_12_10_3  (
            .in0(N__34310),
            .in1(N__33153),
            .in2(_gnd_net_),
            .in3(N__33137),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__50217),
            .ce(),
            .sr(N__49449));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_12_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_12_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_12_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_12_10_4  (
            .in0(N__34228),
            .in1(N__33132),
            .in2(_gnd_net_),
            .in3(N__33116),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__50217),
            .ce(),
            .sr(N__49449));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_12_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_12_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_12_10_5  (
            .in0(N__34311),
            .in1(N__33111),
            .in2(_gnd_net_),
            .in3(N__33089),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__50217),
            .ce(),
            .sr(N__49449));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_12_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_12_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_12_10_6  (
            .in0(N__34229),
            .in1(N__33079),
            .in2(_gnd_net_),
            .in3(N__33086),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50217),
            .ce(),
            .sr(N__49449));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_12_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_12_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_12_11_0  (
            .in0(N__34752),
            .in1(N__33036),
            .in2(_gnd_net_),
            .in3(N__33055),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_12_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_12_11_1 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_12_11_1  (
            .in0(N__33037),
            .in1(N__34754),
            .in2(N__33011),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50206),
            .ce(N__34202),
            .sr(N__49456));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_12_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_12_11_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_12_11_2  (
            .in0(N__34753),
            .in1(_gnd_net_),
            .in2(N__33413),
            .in3(N__33427),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(elapsed_time_ns_1_RNI4EOBB_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_12_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_12_11_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__34756),
            .in2(N__33416),
            .in3(N__33411),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50206),
            .ce(N__34202),
            .sr(N__49456));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_12_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_12_11_4 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_12_11_4  (
            .in0(N__33325),
            .in1(N__33238),
            .in2(N__33359),
            .in3(N__33334),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_11_5 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_11_5  (
            .in0(N__33239),
            .in1(N__33355),
            .in2(N__33338),
            .in3(N__33326),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_12_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_12_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_12_11_6  (
            .in0(N__34751),
            .in1(N__33276),
            .in2(_gnd_net_),
            .in3(N__33292),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_12_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_12_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_12_11_7 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_12_11_7  (
            .in0(N__33277),
            .in1(N__34755),
            .in2(N__33242),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50206),
            .ce(N__34202),
            .sr(N__49456));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_12_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_12_12_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__35011),
            .in2(_gnd_net_),
            .in3(N__35127),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_12_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_12_12_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33212),
            .in3(N__35164),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_12_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_12_13_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_12_13_0  (
            .in0(N__34986),
            .in1(N__39839),
            .in2(N__48065),
            .in3(N__48013),
            .lcout(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_12_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_12_13_1 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_12_13_1  (
            .in0(N__35107),
            .in1(N__35012),
            .in2(_gnd_net_),
            .in3(N__35036),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_12_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_12_13_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_12_13_2  (
            .in0(N__36885),
            .in1(N__38405),
            .in2(_gnd_net_),
            .in3(N__48910),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_12_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_12_13_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__35013),
            .in2(_gnd_net_),
            .in3(N__35037),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__35066),
            .in2(_gnd_net_),
            .in3(N__35091),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_12_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_12_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__35067),
            .in2(_gnd_net_),
            .in3(N__35092),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_0_LC_12_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_12_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_12_14_0 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \phase_controller_inst1.state_0_LC_12_14_0  (
            .in0(N__34988),
            .in1(N__33469),
            .in2(N__33458),
            .in3(N__39846),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50187),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_14_1 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_12_14_1  (
            .in0(N__33470),
            .in1(N__35169),
            .in2(N__35020),
            .in3(N__35134),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50187),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_12_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_12_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__33468),
            .in2(_gnd_net_),
            .in3(N__33453),
            .lcout(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ),
            .ltout(\phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_12_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_12_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_12_14_3 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst1.state_3_LC_12_14_3  (
            .in0(N__35602),
            .in1(N__35680),
            .in2(N__33437),
            .in3(N__33571),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50187),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__35601),
            .in2(_gnd_net_),
            .in3(N__35676),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_12_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_12_14_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a3_1_LC_12_14_5  (
            .in0(N__33546),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46894),
            .lcout(state_ns_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_4_LC_12_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_12_14_6 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_12_14_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.state_4_LC_12_14_6  (
            .in0(N__46895),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33545),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50187),
            .ce(),
            .sr(N__49480));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_12_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_12_15_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_12_15_0  (
            .in0(N__45440),
            .in1(N__41519),
            .in2(N__42882),
            .in3(N__41483),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_12_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_12_15_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_12_15_2  (
            .in0(N__43576),
            .in1(N__33629),
            .in2(_gnd_net_),
            .in3(N__36374),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_15_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_15_3  (
            .in0(N__43577),
            .in1(N__36362),
            .in2(_gnd_net_),
            .in3(N__33620),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_12_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_12_15_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_12_15_4  (
            .in0(N__36335),
            .in1(N__33611),
            .in2(_gnd_net_),
            .in3(N__43578),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_12_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_12_15_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_12_15_5  (
            .in0(N__43579),
            .in1(N__36323),
            .in2(_gnd_net_),
            .in3(N__33602),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_12_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_12_15_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_12_15_6  (
            .in0(N__36311),
            .in1(N__33593),
            .in2(_gnd_net_),
            .in3(N__43580),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_15_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_15_7  (
            .in0(N__43581),
            .in1(N__36296),
            .in2(_gnd_net_),
            .in3(N__33722),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_12_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_12_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__41179),
            .in2(N__41552),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_12_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_12_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__40886),
            .in2(N__37877),
            .in3(N__45041),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_12_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_12_16_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_12_16_2  (
            .in0(N__45042),
            .in1(N__42431),
            .in2(N__36767),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_12_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_12_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__36611),
            .in2(N__42605),
            .in3(N__33641),
            .lcout(\current_shift_inst.un38_control_input_0_s0_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_12_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_12_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__42435),
            .in2(N__33638),
            .in3(N__33623),
            .lcout(\current_shift_inst.un38_control_input_0_s0_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_12_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_12_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__35369),
            .in2(N__42606),
            .in3(N__33614),
            .lcout(\current_shift_inst.un38_control_input_0_s0_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_12_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_12_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__42439),
            .in2(N__35192),
            .in3(N__33605),
            .lcout(\current_shift_inst.un38_control_input_0_s0_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_12_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_12_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__35363),
            .in2(N__42607),
            .in3(N__33596),
            .lcout(\current_shift_inst.un38_control_input_0_s0_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_12_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_12_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__42482),
            .in2(N__35432),
            .in3(N__33584),
            .lcout(\current_shift_inst.un38_control_input_0_s0_8 ),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_12_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_12_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__40793),
            .in2(N__42716),
            .in3(N__33713),
            .lcout(\current_shift_inst.un38_control_input_0_s0_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_12_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_12_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__42486),
            .in2(N__35450),
            .in3(N__33710),
            .lcout(\current_shift_inst.un38_control_input_0_s0_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_12_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_12_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__35546),
            .in2(N__42717),
            .in3(N__33695),
            .lcout(\current_shift_inst.un38_control_input_0_s0_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_12_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_12_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__42490),
            .in2(N__35357),
            .in3(N__33680),
            .lcout(\current_shift_inst.un38_control_input_0_s0_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_12_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_12_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__37760),
            .in2(N__42718),
            .in3(N__33665),
            .lcout(\current_shift_inst.un38_control_input_0_s0_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_12_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_12_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(N__42494),
            .in2(N__35420),
            .in3(N__33662),
            .lcout(\current_shift_inst.un38_control_input_0_s0_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_12_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_12_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__35258),
            .in2(N__42719),
            .in3(N__33659),
            .lcout(\current_shift_inst.un38_control_input_0_s0_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_12_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_12_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__42563),
            .in2(N__35510),
            .in3(N__33656),
            .lcout(\current_shift_inst.un38_control_input_0_s0_16 ),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_12_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_12_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__35411),
            .in2(N__42778),
            .in3(N__33773),
            .lcout(\current_shift_inst.un38_control_input_0_s0_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_12_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_12_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__42567),
            .in2(N__35519),
            .in3(N__33770),
            .lcout(\current_shift_inst.un38_control_input_0_s0_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_12_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_12_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__35405),
            .in2(N__42779),
            .in3(N__33767),
            .lcout(\current_shift_inst.un38_control_input_0_s0_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_12_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_12_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__42571),
            .in2(N__37796),
            .in3(N__33758),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_12_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_12_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__37832),
            .in2(N__42780),
            .in3(N__33749),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_12_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_12_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__42575),
            .in2(N__35441),
            .in3(N__33734),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_12_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_12_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__35525),
            .in2(N__42781),
            .in3(N__33731),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_12_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_12_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__42579),
            .in2(N__35495),
            .in3(N__33728),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_12_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_12_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__42224),
            .in2(N__42782),
            .in3(N__33725),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_12_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_12_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__42583),
            .in2(N__35717),
            .in3(N__33812),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_12_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_12_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__37859),
            .in2(N__42783),
            .in3(N__33809),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_12_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_12_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__42587),
            .in2(N__37889),
            .in3(N__33806),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_12_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_12_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__35501),
            .in2(N__42784),
            .in3(N__33803),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_12_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_12_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__42591),
            .in2(N__41321),
            .in3(N__33794),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_12_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_12_19_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_12_19_7  (
            .in0(N__40766),
            .in1(N__36623),
            .in2(N__43590),
            .in3(N__33791),
            .lcout(\current_shift_inst.control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_12_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_12_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43571),
            .lcout(\current_shift_inst.control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.start_timer_s1_LC_12_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_12_21_3 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_12_21_3  (
            .in0(N__35574),
            .in1(N__36749),
            .in2(_gnd_net_),
            .in3(N__35628),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50171),
            .ce(),
            .sr(N__49509));
    defparam \phase_controller_inst1.S1_LC_12_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_12_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_12_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35629),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50171),
            .ce(),
            .sr(N__49509));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_0 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_0 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49571),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35853),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34055),
            .ce(),
            .sr(N__49406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_13_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_13_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_13_7_2  (
            .in0(N__34739),
            .in1(N__34404),
            .in2(_gnd_net_),
            .in3(N__34374),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_13_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_13_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_13_7_3  (
            .in0(N__33996),
            .in1(N__34038),
            .in2(_gnd_net_),
            .in3(N__34740),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_13_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_13_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_13_7_6  (
            .in0(N__34741),
            .in1(N__34909),
            .in2(_gnd_net_),
            .in3(N__34881),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_13_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_13_8_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_13_8_0  (
            .in0(N__33954),
            .in1(N__33937),
            .in2(N__33842),
            .in3(N__34922),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_13_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_13_8_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_13_8_1  (
            .in0(N__34921),
            .in1(N__33955),
            .in2(N__33941),
            .in3(N__33838),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_13_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_13_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_25_LC_13_8_3  (
            .in0(N__34778),
            .in1(N__33908),
            .in2(_gnd_net_),
            .in3(N__33878),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50253),
            .ce(N__34262),
            .sr(N__49420));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_13_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_13_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_13_8_4  (
            .in0(N__34954),
            .in1(N__33823),
            .in2(_gnd_net_),
            .in3(N__34776),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(elapsed_time_ns_1_RNI2DPBB_0_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_13_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_13_8_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_24_LC_13_8_5  (
            .in0(N__34777),
            .in1(_gnd_net_),
            .in2(N__34958),
            .in3(N__34955),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50253),
            .ce(N__34262),
            .sr(N__49420));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_13_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_13_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_13_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_13_8_6  (
            .in0(N__34905),
            .in1(N__34889),
            .in2(_gnd_net_),
            .in3(N__34780),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50253),
            .ce(N__34262),
            .sr(N__49420));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_13_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_13_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_13_8_7  (
            .in0(N__34779),
            .in1(N__34408),
            .in2(_gnd_net_),
            .in3(N__34385),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50253),
            .ce(N__34262),
            .sr(N__49420));
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_13_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_13_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_31_LC_13_9_7  (
            .in0(N__40277),
            .in1(N__36685),
            .in2(_gnd_net_),
            .in3(N__48856),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50241),
            .ce(N__49832),
            .sr(N__49429));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_10_1 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_10_1  (
            .in0(N__46988),
            .in1(N__43991),
            .in2(N__44296),
            .in3(N__49833),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50229),
            .ce(),
            .sr(N__49440));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_13_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_13_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_13_11_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_13_11_0  (
            .in0(N__38345),
            .in1(N__48921),
            .in2(_gnd_net_),
            .in3(N__36788),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50220),
            .ce(N__47862),
            .sr(N__49450));
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_13_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_13_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_13_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_22_LC_13_11_5  (
            .in0(N__48920),
            .in1(N__47756),
            .in2(_gnd_net_),
            .in3(N__47727),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50220),
            .ce(N__47862),
            .sr(N__49450));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_12_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_12_0  (
            .in0(N__35180),
            .in1(N__34076),
            .in2(N__36023),
            .in3(N__36000),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_12_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_12_1  (
            .in0(N__34075),
            .in1(N__36021),
            .in2(N__36002),
            .in3(N__35179),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_13_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_13_12_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_23_LC_13_12_3  (
            .in0(N__47655),
            .in1(N__48922),
            .in2(_gnd_net_),
            .in3(N__47675),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50209),
            .ce(N__47861),
            .sr(N__49457));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_13_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_13_12_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_13_12_4  (
            .in0(N__36987),
            .in1(N__38285),
            .in2(_gnd_net_),
            .in3(N__48880),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_LC_13_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_13_13_2 .LUT_INIT=16'b1010111000101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_13_13_2  (
            .in0(N__35108),
            .in1(N__35168),
            .in2(N__35021),
            .in3(N__35135),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(),
            .sr(N__49465));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_13_3 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_13_13_3  (
            .in0(N__35817),
            .in1(N__35801),
            .in2(_gnd_net_),
            .in3(N__35864),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(),
            .sr(N__49465));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_13_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_13_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_13_13_4 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_13_13_4  (
            .in0(N__36169),
            .in1(N__35096),
            .in2(N__35078),
            .in3(N__37116),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(),
            .sr(N__49465));
    defparam \phase_controller_inst1.start_timer_tr_LC_13_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_13_5 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_13_13_5  (
            .in0(N__35051),
            .in1(N__35045),
            .in2(N__46916),
            .in3(N__35038),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(),
            .sr(N__49465));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_13_13_6  (
            .in0(N__35039),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(),
            .sr(N__49465));
    defparam \phase_controller_inst1.state_1_LC_13_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_13_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_13_13_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst1.state_1_LC_13_13_7  (
            .in0(N__34987),
            .in1(N__39845),
            .in2(_gnd_net_),
            .in3(N__47969),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(),
            .sr(N__49465));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_13_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_13_14_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_13_14_0  (
            .in0(N__36277),
            .in1(N__35976),
            .in2(N__35243),
            .in3(N__35252),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_13_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_13_14_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_13_14_1  (
            .in0(N__35251),
            .in1(N__36276),
            .in2(N__35981),
            .in3(N__35239),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_13_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_13_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_13_14_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_24_LC_13_14_2  (
            .in0(N__40586),
            .in1(N__40628),
            .in2(_gnd_net_),
            .in3(N__48935),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50193),
            .ce(N__47860),
            .sr(N__49473));
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_13_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_13_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_13_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_25_LC_13_14_3  (
            .in0(N__48931),
            .in1(N__40678),
            .in2(_gnd_net_),
            .in3(N__40697),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50193),
            .ce(N__47860),
            .sr(N__49473));
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_13_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_13_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_13_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_31_LC_13_14_4  (
            .in0(N__40276),
            .in1(N__36692),
            .in2(_gnd_net_),
            .in3(N__48936),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50193),
            .ce(N__47860),
            .sr(N__49473));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_13_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_13_14_5 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_13_14_5  (
            .in0(N__35218),
            .in1(N__36247),
            .in2(N__36062),
            .in3(N__35227),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_13_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_13_14_6 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_13_14_6  (
            .in0(N__36246),
            .in1(N__36057),
            .in2(N__35231),
            .in3(N__35219),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_13_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_13_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_13_14_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_30_LC_13_14_7  (
            .in0(N__35777),
            .in1(_gnd_net_),
            .in2(N__48938),
            .in3(N__39175),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50193),
            .ce(N__47860),
            .sr(N__49473));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_15_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_15_0  (
            .in0(N__36473),
            .in1(N__35210),
            .in2(_gnd_net_),
            .in3(N__43582),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_13_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_13_15_2 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_13_15_2  (
            .in0(N__41060),
            .in1(N__42771),
            .in2(N__41018),
            .in3(N__45442),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_13_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_13_15_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_13_15_5  (
            .in0(N__45441),
            .in1(N__41141),
            .in2(N__42883),
            .in3(N__41108),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_15_6 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_15_6  (
            .in0(N__43073),
            .in1(N__45443),
            .in2(N__43034),
            .in3(N__42772),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_13_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_13_16_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_13_16_0  (
            .in0(N__41377),
            .in1(N__45438),
            .in2(N__42720),
            .in3(N__41345),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_13_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_13_16_1 .LUT_INIT=16'b0001101100011011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_13_16_1  (
            .in0(N__43551),
            .in1(N__36422),
            .in2(N__35348),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_13_16_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_13_16_2  (
            .in0(N__36413),
            .in1(N__35327),
            .in2(_gnd_net_),
            .in3(N__43552),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_13_16_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_13_16_3  (
            .in0(N__43553),
            .in1(N__35312),
            .in2(_gnd_net_),
            .in3(N__36404),
            .lcout(\current_shift_inst.control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_13_16_4 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_13_16_4  (
            .in0(N__35294),
            .in1(N__43554),
            .in2(_gnd_net_),
            .in3(N__36395),
            .lcout(\current_shift_inst.control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_13_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_13_16_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_13_16_5  (
            .in0(N__43555),
            .in1(N__36587),
            .in2(_gnd_net_),
            .in3(N__35276),
            .lcout(\current_shift_inst.control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_13_16_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_13_16_6  (
            .in0(N__42502),
            .in1(N__45439),
            .in2(N__41440),
            .in3(N__41405),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_13_16_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_13_16_7  (
            .in0(N__45437),
            .in1(N__42498),
            .in2(N__40949),
            .in3(N__40984),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_17_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_17_0  (
            .in0(N__45435),
            .in1(N__42504),
            .in2(N__39980),
            .in3(N__40009),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_17_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_17_1  (
            .in0(N__42503),
            .in1(N__45431),
            .in2(N__41615),
            .in3(N__41573),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_13_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_13_17_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_13_17_2  (
            .in0(N__45432),
            .in1(N__42511),
            .in2(N__41974),
            .in3(N__41927),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_13_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_13_17_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_13_17_3  (
            .in0(N__40010),
            .in1(N__45436),
            .in2(N__42721),
            .in3(N__39978),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_13_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_13_17_4 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_13_17_4  (
            .in0(N__45433),
            .in1(N__41897),
            .in2(N__41087),
            .in3(N__42512),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_13_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_13_17_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_13_17_5  (
            .in0(N__41857),
            .in1(N__45434),
            .in2(N__42722),
            .in3(N__41813),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_17_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_17_6  (
            .in0(N__35399),
            .in1(N__36578),
            .in2(_gnd_net_),
            .in3(N__43556),
            .lcout(\current_shift_inst.control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_18_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_18_0  (
            .in0(N__36656),
            .in1(N__35384),
            .in2(_gnd_net_),
            .in3(N__43558),
            .lcout(\current_shift_inst.control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_13_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_13_18_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_13_18_1  (
            .in0(N__45277),
            .in1(N__44777),
            .in2(N__42861),
            .in3(N__44816),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_18_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_18_2  (
            .in0(N__36665),
            .in1(N__35540),
            .in2(_gnd_net_),
            .in3(N__43557),
            .lcout(\current_shift_inst.control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_13_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_13_18_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_13_18_3  (
            .in0(N__45279),
            .in1(N__43138),
            .in2(N__42862),
            .in3(N__43097),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_13_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_13_18_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_13_18_4  (
            .in0(N__45280),
            .in1(N__42723),
            .in2(N__41792),
            .in3(N__41753),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_13_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_13_18_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_13_18_5  (
            .in0(N__45278),
            .in1(N__41252),
            .in2(N__42863),
            .in3(N__41210),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_18_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_18_7  (
            .in0(N__42730),
            .in1(N__45281),
            .in2(N__42209),
            .in3(N__42170),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_13_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_13_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_13_19_0  (
            .in0(N__45282),
            .in1(N__39949),
            .in2(N__42864),
            .in3(N__39908),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_19_1 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_19_1  (
            .in0(N__35486),
            .in1(N__36647),
            .in2(_gnd_net_),
            .in3(N__43567),
            .lcout(\current_shift_inst.control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_19_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_19_2  (
            .in0(N__43561),
            .in1(N__35468),
            .in2(_gnd_net_),
            .in3(N__36518),
            .lcout(\current_shift_inst.control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_19_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_19_3  (
            .in0(N__35753),
            .in1(N__36506),
            .in2(_gnd_net_),
            .in3(N__43562),
            .lcout(\current_shift_inst.control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_19_4 .LUT_INIT=16'b0011010100110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_19_4  (
            .in0(N__36491),
            .in1(N__35735),
            .in2(N__43589),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_13_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_13_19_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_13_19_6  (
            .in0(N__45283),
            .in1(N__41303),
            .in2(N__42865),
            .in3(N__39599),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_19_7 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_19_7  (
            .in0(N__35708),
            .in1(N__36482),
            .in2(_gnd_net_),
            .in3(N__43566),
            .lcout(\current_shift_inst.control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_2_LC_13_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_13_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_13_20_2 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_2_LC_13_20_2  (
            .in0(N__35623),
            .in1(N__48047),
            .in2(N__35690),
            .in3(N__48020),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50175),
            .ce(),
            .sr(N__49503));
    defparam \phase_controller_inst1.T01_LC_13_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_LC_13_20_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.T01_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__35641),
            .in2(_gnd_net_),
            .in3(N__35624),
            .lcout(T01_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50175),
            .ce(),
            .sr(N__49503));
    defparam \current_shift_inst.timer_s1.running_LC_13_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_21_6 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_21_6  (
            .in0(N__36727),
            .in1(N__36752),
            .in2(_gnd_net_),
            .in3(N__37948),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50172),
            .ce(),
            .sr(N__49507));
    defparam \current_shift_inst.stop_timer_s1_LC_13_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_13_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_13_21_7 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_13_21_7  (
            .in0(N__36751),
            .in1(N__36728),
            .in2(N__35630),
            .in3(N__35575),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50172),
            .ce(),
            .sr(N__49507));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__37943),
            .in2(_gnd_net_),
            .in3(N__36725),
            .lcout(\current_shift_inst.timer_s1.N_162_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_13_30_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_30_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_30_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_30_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39856),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50165),
            .ce(),
            .sr(N__49539));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_14_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_14_6_6 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_14_6_6  (
            .in0(N__35796),
            .in1(N__35831),
            .in2(_gnd_net_),
            .in3(N__35860),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_199_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_14_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_14_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_14_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_30_LC_14_7_2  (
            .in0(N__35769),
            .in1(N__39179),
            .in2(_gnd_net_),
            .in3(N__48908),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50276),
            .ce(N__49806),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_14_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_14_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35826),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_14_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_14_8_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_14_8_1  (
            .in0(N__47448),
            .in1(N__50354),
            .in2(N__40679),
            .in3(N__39173),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_14_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_14_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_14_8_2  (
            .in0(N__35932),
            .in1(N__38814),
            .in2(_gnd_net_),
            .in3(N__48877),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_8_3  (
            .in0(N__35827),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35797),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_198_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_14_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_14_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_14_8_7  (
            .in0(N__48876),
            .in1(N__35773),
            .in2(_gnd_net_),
            .in3(N__39174),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_14_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_14_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_14_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_14_9_4  (
            .in0(N__48855),
            .in1(N__38512),
            .in2(_gnd_net_),
            .in3(N__37152),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50254),
            .ce(N__49805),
            .sr(N__49421));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_14_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_14_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_14_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_14_9_6  (
            .in0(N__48854),
            .in1(N__35928),
            .in2(_gnd_net_),
            .in3(N__38816),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50254),
            .ce(N__49805),
            .sr(N__49421));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_14_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_14_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_14_10_2  (
            .in0(N__48888),
            .in1(N__35933),
            .in2(_gnd_net_),
            .in3(N__38815),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50242),
            .ce(N__47866),
            .sr(N__49430));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_14_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_14_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_14_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_14_10_5  (
            .in0(N__36991),
            .in1(N__38284),
            .in2(_gnd_net_),
            .in3(N__48890),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50242),
            .ce(N__47866),
            .sr(N__49430));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_14_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_14_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_14_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_14_10_6  (
            .in0(N__48889),
            .in1(N__44055),
            .in2(_gnd_net_),
            .in3(N__44035),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50242),
            .ce(N__47866),
            .sr(N__49430));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(N__35912),
            .in2(N__37124),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_11_1  (
            .in0(N__36223),
            .in1(N__37087),
            .in2(_gnd_net_),
            .in3(N__35900),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__50230),
            .ce(),
            .sr(N__49441));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_11_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_11_2  (
            .in0(N__36227),
            .in1(N__37054),
            .in2(N__35897),
            .in3(N__35882),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__50230),
            .ce(),
            .sr(N__49441));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_11_3  (
            .in0(N__36224),
            .in1(N__37027),
            .in2(_gnd_net_),
            .in3(N__35879),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__50230),
            .ce(),
            .sr(N__49441));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_11_4  (
            .in0(N__36228),
            .in1(N__37399),
            .in2(_gnd_net_),
            .in3(N__35876),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__50230),
            .ce(),
            .sr(N__49441));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_11_5  (
            .in0(N__36225),
            .in1(N__37369),
            .in2(_gnd_net_),
            .in3(N__35873),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__50230),
            .ce(),
            .sr(N__49441));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_11_6  (
            .in0(N__36229),
            .in1(N__37327),
            .in2(_gnd_net_),
            .in3(N__35960),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__50230),
            .ce(),
            .sr(N__49441));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_11_7  (
            .in0(N__36226),
            .in1(N__37306),
            .in2(_gnd_net_),
            .in3(N__35957),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__50230),
            .ce(),
            .sr(N__49441));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_12_0  (
            .in0(N__36196),
            .in1(N__37258),
            .in2(_gnd_net_),
            .in3(N__35954),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__50221),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_12_1  (
            .in0(N__36173),
            .in1(N__37219),
            .in2(_gnd_net_),
            .in3(N__35951),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__50221),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_12_2  (
            .in0(N__36193),
            .in1(N__37180),
            .in2(_gnd_net_),
            .in3(N__35948),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__50221),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_12_3  (
            .in0(N__36174),
            .in1(N__37594),
            .in2(_gnd_net_),
            .in3(N__35945),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__50221),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_12_4  (
            .in0(N__36194),
            .in1(N__37570),
            .in2(_gnd_net_),
            .in3(N__35942),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__50221),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_12_5  (
            .in0(N__36175),
            .in1(N__37534),
            .in2(_gnd_net_),
            .in3(N__35939),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__50221),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_12_6  (
            .in0(N__36195),
            .in1(N__37495),
            .in2(_gnd_net_),
            .in3(N__35936),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__50221),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_12_7  (
            .in0(N__36176),
            .in1(N__39115),
            .in2(_gnd_net_),
            .in3(N__36041),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__50221),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_13_0  (
            .in0(N__36161),
            .in1(N__39100),
            .in2(_gnd_net_),
            .in3(N__36038),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__50210),
            .ce(),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_13_1  (
            .in0(N__36165),
            .in1(N__36833),
            .in2(_gnd_net_),
            .in3(N__36035),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__50210),
            .ce(),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_13_2  (
            .in0(N__36162),
            .in1(N__36850),
            .in2(_gnd_net_),
            .in3(N__36032),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__50210),
            .ce(),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_13_3  (
            .in0(N__36166),
            .in1(N__36933),
            .in2(_gnd_net_),
            .in3(N__36029),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__50210),
            .ce(),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_13_4  (
            .in0(N__36163),
            .in1(N__36960),
            .in2(_gnd_net_),
            .in3(N__36026),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__50210),
            .ce(),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_13_5  (
            .in0(N__36167),
            .in1(N__36022),
            .in2(_gnd_net_),
            .in3(N__36005),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__50210),
            .ce(),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_13_6  (
            .in0(N__36164),
            .in1(N__36001),
            .in2(_gnd_net_),
            .in3(N__35984),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__50210),
            .ce(),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_13_7  (
            .in0(N__36168),
            .in1(N__35980),
            .in2(_gnd_net_),
            .in3(N__35963),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__50210),
            .ce(),
            .sr(N__49458));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_14_0  (
            .in0(N__36220),
            .in1(N__36278),
            .in2(_gnd_net_),
            .in3(N__36263),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__50200),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_14_1  (
            .in0(N__36216),
            .in1(N__44614),
            .in2(_gnd_net_),
            .in3(N__36260),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__50200),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_14_2  (
            .in0(N__36221),
            .in1(N__44589),
            .in2(_gnd_net_),
            .in3(N__36257),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__50200),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_14_3  (
            .in0(N__36217),
            .in1(N__45526),
            .in2(_gnd_net_),
            .in3(N__36254),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__50200),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_14_4  (
            .in0(N__36222),
            .in1(N__45505),
            .in2(_gnd_net_),
            .in3(N__36251),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__50200),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_14_5  (
            .in0(N__36218),
            .in1(N__36248),
            .in2(_gnd_net_),
            .in3(N__36233),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__50200),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_14_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_14_6  (
            .in0(N__36061),
            .in1(N__36219),
            .in2(_gnd_net_),
            .in3(N__36065),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50200),
            .ce(),
            .sr(N__49466));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__45083),
            .in2(N__41180),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__40899),
            .in2(N__40862),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__42745),
            .in2(N__36707),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_14_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__36599),
            .in2(N__42876),
            .in3(N__36377),
            .lcout(\current_shift_inst.un38_control_input_0_s1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__42749),
            .in2(N__41456),
            .in3(N__36365),
            .lcout(\current_shift_inst.un38_control_input_0_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__39245),
            .in2(N__42877),
            .in3(N__36353),
            .lcout(\current_shift_inst.un38_control_input_0_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__42753),
            .in2(N__36350),
            .in3(N__36326),
            .lcout(\current_shift_inst.un38_control_input_0_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__37781),
            .in2(N__42878),
            .in3(N__36314),
            .lcout(\current_shift_inst.un38_control_input_0_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__42608),
            .in2(N__41156),
            .in3(N__36299),
            .lcout(\current_shift_inst.un38_control_input_0_s1_8 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__40778),
            .in2(N__42792),
            .in3(N__36281),
            .lcout(\current_shift_inst.un38_control_input_0_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__42612),
            .in2(N__37628),
            .in3(N__36467),
            .lcout(\current_shift_inst.un38_control_input_0_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_14_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__37766),
            .in2(N__42793),
            .in3(N__36452),
            .lcout(\current_shift_inst.un38_control_input_0_s1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__42616),
            .in2(N__37775),
            .in3(N__36437),
            .lcout(\current_shift_inst.un38_control_input_0_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_14_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__37634),
            .in2(N__42794),
            .in3(N__36425),
            .lcout(\current_shift_inst.un38_control_input_0_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_14_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_14_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__42620),
            .in2(N__37619),
            .in3(N__36416),
            .lcout(\current_shift_inst.un38_control_input_0_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_14_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_14_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__37610),
            .in2(N__42795),
            .in3(N__36407),
            .lcout(\current_shift_inst.un38_control_input_0_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_14_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__42796),
            .in2(N__39881),
            .in3(N__36398),
            .lcout(\current_shift_inst.un38_control_input_0_s1_16 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_14_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__37850),
            .in2(N__42889),
            .in3(N__36389),
            .lcout(\current_shift_inst.un38_control_input_0_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_14_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__42800),
            .in2(N__37739),
            .in3(N__36581),
            .lcout(\current_shift_inst.un38_control_input_0_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_14_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_14_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__37745),
            .in2(N__42890),
            .in3(N__36572),
            .lcout(\current_shift_inst.un38_control_input_0_s1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__42804),
            .in2(N__37805),
            .in3(N__36557),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__37751),
            .in2(N__42891),
            .in3(N__36542),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__42808),
            .in2(N__36539),
            .in3(N__36521),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__37724),
            .in2(N__42892),
            .in3(N__36509),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__39260),
            .in2(N__42893),
            .in3(N__36494),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__42815),
            .in2(N__37907),
            .in3(N__36485),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__37895),
            .in2(N__42894),
            .in3(N__36476),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__42819),
            .in2(N__37823),
            .in3(N__36659),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__37811),
            .in2(N__42895),
            .in3(N__36650),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__42823),
            .in2(N__37844),
            .in3(N__36641),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_14_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_14_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__42825),
            .in2(N__42968),
            .in3(N__36629),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_14_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_14_18_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_14_18_7  (
            .in0(N__45284),
            .in1(N__42824),
            .in2(_gnd_net_),
            .in3(N__36626),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_14_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_14_19_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_14_19_4  (
            .in0(N__42786),
            .in1(N__45223),
            .in2(N__42034),
            .in3(N__41998),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44997),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50178),
            .ce(N__44954),
            .sr(N__49495));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_14_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_14_19_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_14_19_6  (
            .in0(N__42787),
            .in1(N__45224),
            .in2(N__42035),
            .in3(N__41999),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_19_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_19_7  (
            .in0(N__45222),
            .in1(N__42788),
            .in2(N__42146),
            .in3(N__42109),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_21_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_21_3  (
            .in0(N__36750),
            .in1(N__37947),
            .in2(_gnd_net_),
            .in3(N__36726),
            .lcout(\current_shift_inst.timer_s1.N_163_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_22_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_22_4  (
            .in0(N__45335),
            .in1(N__42145),
            .in2(N__42910),
            .in3(N__42113),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_15_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_15_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_15_6_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_15_6_4  (
            .in0(N__44105),
            .in1(N__48906),
            .in2(_gnd_net_),
            .in3(N__44126),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50299),
            .ce(N__47872),
            .sr(N__49398));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_15_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_15_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_15_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_15_7_0  (
            .in0(N__46487),
            .in1(N__46340),
            .in2(_gnd_net_),
            .in3(N__48907),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50289),
            .ce(N__47871),
            .sr(N__49402));
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_15_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_15_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_21_LC_15_8_4  (
            .in0(N__39770),
            .in1(N__39799),
            .in2(_gnd_net_),
            .in3(N__48879),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(N__47869),
            .sr(N__49408));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_15_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_15_8_6  (
            .in0(N__40043),
            .in1(N__40073),
            .in2(_gnd_net_),
            .in3(N__48878),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(N__47869),
            .sr(N__49408));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_15_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_15_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_15_9_0  (
            .in0(N__40275),
            .in1(N__36684),
            .in2(_gnd_net_),
            .in3(N__48776),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_15_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_15_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_15_9_2  (
            .in0(N__38796),
            .in1(N__44027),
            .in2(N__47792),
            .in3(N__47079),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_15_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_15_9_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_15_9_3  (
            .in0(N__47720),
            .in1(N__47643),
            .in2(N__40627),
            .in3(N__39767),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_15_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_15_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_15_9_4  (
            .in0(N__36818),
            .in1(N__36803),
            .in2(N__36812),
            .in3(N__36809),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_15_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_15_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_15_9_5  (
            .in0(N__44094),
            .in1(N__47907),
            .in2(N__43938),
            .in3(N__47199),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_15_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_15_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_15_9_6  (
            .in0(N__44059),
            .in1(N__44028),
            .in2(_gnd_net_),
            .in3(N__48777),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_9_7  (
            .in0(N__48778),
            .in1(N__38505),
            .in2(_gnd_net_),
            .in3(N__37156),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_15_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_15_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_15_10_0  (
            .in0(N__38273),
            .in1(N__38336),
            .in2(N__38400),
            .in3(N__40064),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_15_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_15_10_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_15_10_1  (
            .in0(N__40322),
            .in1(N__38504),
            .in2(N__36797),
            .in3(N__36794),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_15_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_15_10_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_15_10_2  (
            .in0(N__47508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40118),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_15_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_15_10_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_15_10_4  (
            .in0(N__38337),
            .in1(N__48884),
            .in2(_gnd_net_),
            .in3(N__36781),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(elapsed_time_ns_1_RNITUBN9_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_15_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_15_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_15_10_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_15_10_5  (
            .in0(N__48885),
            .in1(_gnd_net_),
            .in2(N__36770),
            .in3(N__38338),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50255),
            .ce(N__49791),
            .sr(N__49422));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_15_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_15_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_15_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_15_10_6  (
            .in0(N__36893),
            .in1(N__38399),
            .in2(_gnd_net_),
            .in3(N__48887),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50255),
            .ce(N__49791),
            .sr(N__49422));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_15_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_15_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_15_10_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_15_10_7  (
            .in0(N__48886),
            .in1(_gnd_net_),
            .in2(N__36995),
            .in3(N__38274),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50255),
            .ce(N__49791),
            .sr(N__49422));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_15_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_15_11_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_15_11_0  (
            .in0(N__36940),
            .in1(N__36917),
            .in2(N__36965),
            .in3(N__36902),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_15_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_15_11_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_15_11_1  (
            .in0(N__36901),
            .in1(N__36964),
            .in2(N__36944),
            .in3(N__36916),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_15_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_15_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_15_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_20_LC_15_11_2  (
            .in0(N__43889),
            .in1(N__43919),
            .in2(_gnd_net_),
            .in3(N__48905),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50243),
            .ce(N__47867),
            .sr(N__49431));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_15_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_15_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_15_11_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_15_11_5  (
            .in0(N__40124),
            .in1(N__48891),
            .in2(_gnd_net_),
            .in3(N__40097),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50243),
            .ce(N__47867),
            .sr(N__49431));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_15_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_15_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_15_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_15_11_6  (
            .in0(N__48893),
            .in1(N__47520),
            .in2(_gnd_net_),
            .in3(N__47543),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50243),
            .ce(N__47867),
            .sr(N__49431));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_15_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_15_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_15_11_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_15_11_7  (
            .in0(N__38404),
            .in1(N__48892),
            .in2(_gnd_net_),
            .in3(N__36892),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50243),
            .ce(N__47867),
            .sr(N__49431));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_12_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_12_0  (
            .in0(N__36832),
            .in1(N__47891),
            .in2(N__36869),
            .in3(N__36849),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_12_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_12_1  (
            .in0(N__47890),
            .in1(N__36868),
            .in2(N__36851),
            .in3(N__36831),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_15_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_15_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_15_12_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_15_12_4  (
            .in0(N__43724),
            .in1(N__46460),
            .in2(_gnd_net_),
            .in3(N__48903),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50231),
            .ce(N__47863),
            .sr(N__49442));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_15_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_15_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_15_12_5  (
            .in0(N__48901),
            .in1(N__43700),
            .in2(_gnd_net_),
            .in3(N__46384),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50231),
            .ce(N__47863),
            .sr(N__49442));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_15_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_15_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_15_12_6  (
            .in0(N__40331),
            .in1(N__40301),
            .in2(_gnd_net_),
            .in3(N__48904),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50231),
            .ce(N__47863),
            .sr(N__49442));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_15_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_15_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_15_12_7  (
            .in0(N__48902),
            .in1(N__38516),
            .in2(_gnd_net_),
            .in3(N__37157),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50231),
            .ce(N__47863),
            .sr(N__49442));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_15_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_15_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__37094),
            .in2(N__37136),
            .in3(N__37117),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_15_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_15_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__39056),
            .in2(N__37073),
            .in3(N__37088),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_15_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_15_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__37064),
            .in2(N__37040),
            .in3(N__37058),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_15_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_15_13_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_15_13_3  (
            .in0(N__37031),
            .in1(N__37013),
            .in2(N__37007),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_15_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_15_13_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_15_13_4  (
            .in0(N__37400),
            .in1(N__37376),
            .in2(N__37385),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_15_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_15_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_15_13_5  (
            .in0(N__37370),
            .in1(N__37355),
            .in2(N__37349),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_15_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_15_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__37313),
            .in2(N__37340),
            .in3(N__37328),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_15_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_15_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_15_13_7  (
            .in0(N__37307),
            .in1(N__37292),
            .in2(N__37283),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_15_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_15_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__37274),
            .in2(N__37244),
            .in3(N__37262),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_15_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_15_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__37232),
            .in2(N__37205),
            .in3(N__37220),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_15_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_15_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__37196),
            .in2(N__37166),
            .in3(N__37184),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_15_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_15_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__37604),
            .in2(N__37580),
            .in3(N__37595),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_15_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_15_14_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_15_14_4  (
            .in0(N__37571),
            .in1(N__37556),
            .in2(N__37544),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_15_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_15_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_15_14_5  (
            .in0(N__37535),
            .in1(N__39062),
            .in2(N__37520),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_15_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_15_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__37508),
            .in2(N__37481),
            .in3(N__37496),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_15_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_15_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__39131),
            .in2(N__39080),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_15_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_15_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__37472),
            .in2(N__37463),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_15_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_15_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__37451),
            .in2(N__37442),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_15_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_15_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__37427),
            .in2(N__37415),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_15_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_15_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__37718),
            .in2(N__37706),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_15_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_15_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__44573),
            .in2(N__44639),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_15_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_15_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(N__45491),
            .in2(N__44564),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_15_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_15_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__37691),
            .in2(N__37679),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_15_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_15_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37664),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_15_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_15_16_0 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_15_16_0  (
            .in0(N__41537),
            .in1(N__42857),
            .in2(N__42083),
            .in3(N__45383),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_15_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_15_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_15_16_1  (
            .in0(N__45378),
            .in1(N__40985),
            .in2(N__42902),
            .in3(N__40948),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_16_2 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_16_2  (
            .in0(N__41926),
            .in1(N__42858),
            .in2(N__41975),
            .in3(N__45384),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_15_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_15_16_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_15_16_3  (
            .in0(N__45385),
            .in1(N__42859),
            .in2(N__41441),
            .in3(N__41401),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_15_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_15_16_4 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_15_16_4  (
            .in0(N__43069),
            .in1(N__45377),
            .in2(N__43029),
            .in3(N__42854),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41048),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_15_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_15_16_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_15_16_6  (
            .in0(N__41344),
            .in1(N__42856),
            .in2(N__41381),
            .in3(N__45382),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_15_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_15_16_7 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_15_16_7  (
            .in0(N__42855),
            .in1(N__44776),
            .in2(N__45447),
            .in3(N__44812),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_17_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_17_0  (
            .in0(N__42076),
            .in1(N__45407),
            .in2(N__42896),
            .in3(N__41536),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_15_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_15_17_1 .LUT_INIT=16'b1010000010101111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_15_17_1  (
            .in0(N__41638),
            .in1(N__42827),
            .in2(N__45451),
            .in3(N__41675),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_15_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_15_17_2 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_15_17_2  (
            .in0(N__42831),
            .in1(N__41809),
            .in2(N__41858),
            .in3(N__45410),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_15_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_15_17_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_15_17_3  (
            .in0(N__45409),
            .in1(N__42826),
            .in2(N__41752),
            .in3(N__41791),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_17_4 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_17_4  (
            .in0(N__42832),
            .in1(N__43090),
            .in2(N__43139),
            .in3(N__45414),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_15_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_15_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41369),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_17_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_17_6  (
            .in0(N__41896),
            .in1(N__45408),
            .in2(N__42897),
            .in3(N__41079),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_17_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_17_7  (
            .in0(N__45415),
            .in1(N__42833),
            .in2(N__42169),
            .in3(N__42208),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_18_0 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_18_0  (
            .in0(N__41671),
            .in1(N__45390),
            .in2(N__41639),
            .in3(N__42839),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_18_1 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_18_1  (
            .in0(N__42837),
            .in1(N__39656),
            .in2(N__45449),
            .in3(N__39619),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_18_2 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_18_2  (
            .in0(N__39443),
            .in1(N__42838),
            .in2(N__39710),
            .in3(N__45396),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_18_3 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_18_3  (
            .in0(N__42841),
            .in1(N__41725),
            .in2(N__45448),
            .in3(N__41708),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_18_4 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_18_4  (
            .in0(N__41707),
            .in1(N__45386),
            .in2(N__41726),
            .in3(N__42840),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40002),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_18_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_18_6  (
            .in0(N__42285),
            .in1(N__42842),
            .in2(N__42263),
            .in3(N__45391),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_15_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_15_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_15_18_7  (
            .in0(N__45392),
            .in1(N__41302),
            .in2(N__42898),
            .in3(N__39597),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41948),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_19_1 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_19_1  (
            .in0(N__45221),
            .in1(N__42847),
            .in2(N__39442),
            .in3(N__39700),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_15_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_15_19_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_15_19_2  (
            .in0(N__39699),
            .in1(N__45219),
            .in2(_gnd_net_),
            .in3(N__39435),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_19_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_19_5  (
            .in0(N__45218),
            .in1(N__40817),
            .in2(N__40909),
            .in3(N__40847),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40964),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_19_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_19_7  (
            .in0(N__45220),
            .in1(N__42846),
            .in2(N__39655),
            .in3(N__39618),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41418),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41231),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42245),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_15_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_15_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41771),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_21_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__37949),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_15_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_15_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41660),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_5_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_5_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_5_0  (
            .in0(N__38178),
            .in1(N__43854),
            .in2(_gnd_net_),
            .in3(N__37922),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_5_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__50317),
            .ce(N__38055),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_5_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_5_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_5_1  (
            .in0(N__38162),
            .in1(N__43824),
            .in2(_gnd_net_),
            .in3(N__37919),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__50317),
            .ce(N__38055),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_5_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_5_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_5_2  (
            .in0(N__38179),
            .in1(N__38559),
            .in2(_gnd_net_),
            .in3(N__37916),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__50317),
            .ce(N__38055),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_5_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_5_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_5_3  (
            .in0(N__38163),
            .in1(N__38530),
            .in2(_gnd_net_),
            .in3(N__37913),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__50317),
            .ce(N__38055),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_5_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_5_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_5_4  (
            .in0(N__38180),
            .in1(N__38472),
            .in2(_gnd_net_),
            .in3(N__37910),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__50317),
            .ce(N__38055),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_5_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_5_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_5_5  (
            .in0(N__38164),
            .in1(N__38445),
            .in2(_gnd_net_),
            .in3(N__37976),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__50317),
            .ce(N__38055),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_5_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_5_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_5_6  (
            .in0(N__38181),
            .in1(N__38419),
            .in2(_gnd_net_),
            .in3(N__37973),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__50317),
            .ce(N__38055),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_5_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_5_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_5_7  (
            .in0(N__38165),
            .in1(N__38359),
            .in2(_gnd_net_),
            .in3(N__37970),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__50317),
            .ce(N__38055),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_6_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_6_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_6_0  (
            .in0(N__38161),
            .in1(N__38301),
            .in2(_gnd_net_),
            .in3(N__37967),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_6_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__50310),
            .ce(N__38054),
            .sr(N__49395));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_6_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_6_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_6_1  (
            .in0(N__38173),
            .in1(N__38238),
            .in2(_gnd_net_),
            .in3(N__37964),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__50310),
            .ce(N__38054),
            .sr(N__49395));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_6_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_6_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_6_2  (
            .in0(N__38158),
            .in1(N__38212),
            .in2(_gnd_net_),
            .in3(N__37961),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__50310),
            .ce(N__38054),
            .sr(N__49395));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_6_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_6_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_6_3  (
            .in0(N__38170),
            .in1(N__38773),
            .in2(_gnd_net_),
            .in3(N__37958),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__50310),
            .ce(N__38054),
            .sr(N__49395));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_6_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_6_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_6_4  (
            .in0(N__38159),
            .in1(N__38748),
            .in2(_gnd_net_),
            .in3(N__37955),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__50310),
            .ce(N__38054),
            .sr(N__49395));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_6_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_6_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_6_5  (
            .in0(N__38171),
            .in1(N__38721),
            .in2(_gnd_net_),
            .in3(N__37952),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__50310),
            .ce(N__38054),
            .sr(N__49395));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_6_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_6_6  (
            .in0(N__38160),
            .in1(N__38695),
            .in2(_gnd_net_),
            .in3(N__38006),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__50310),
            .ce(N__38054),
            .sr(N__49395));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_6_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_6_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_6_7  (
            .in0(N__38172),
            .in1(N__38673),
            .in2(_gnd_net_),
            .in3(N__38003),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__50310),
            .ce(N__38054),
            .sr(N__49395));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_7_0  (
            .in0(N__38154),
            .in1(N__38640),
            .in2(_gnd_net_),
            .in3(N__38000),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__50300),
            .ce(N__38056),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_7_1  (
            .in0(N__38166),
            .in1(N__38616),
            .in2(_gnd_net_),
            .in3(N__37997),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__50300),
            .ce(N__38056),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_7_2  (
            .in0(N__38155),
            .in1(N__38586),
            .in2(_gnd_net_),
            .in3(N__37994),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__50300),
            .ce(N__38056),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_7_3  (
            .in0(N__38167),
            .in1(N__39048),
            .in2(_gnd_net_),
            .in3(N__37991),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__50300),
            .ce(N__38056),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_7_4  (
            .in0(N__38156),
            .in1(N__39024),
            .in2(_gnd_net_),
            .in3(N__37988),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__50300),
            .ce(N__38056),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_7_5  (
            .in0(N__38168),
            .in1(N__38991),
            .in2(_gnd_net_),
            .in3(N__37985),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__50300),
            .ce(N__38056),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_7_6  (
            .in0(N__38157),
            .in1(N__38962),
            .in2(_gnd_net_),
            .in3(N__37982),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__50300),
            .ce(N__38056),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_7_7  (
            .in0(N__38169),
            .in1(N__38932),
            .in2(_gnd_net_),
            .in3(N__37979),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__50300),
            .ce(N__38056),
            .sr(N__49399));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_8_0  (
            .in0(N__38174),
            .in1(N__38901),
            .in2(_gnd_net_),
            .in3(N__38198),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__50290),
            .ce(N__38057),
            .sr(N__49403));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_8_1  (
            .in0(N__38182),
            .in1(N__38877),
            .in2(_gnd_net_),
            .in3(N__38195),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__50290),
            .ce(N__38057),
            .sr(N__49403));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_8_2  (
            .in0(N__38175),
            .in1(N__38853),
            .in2(_gnd_net_),
            .in3(N__38192),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__50290),
            .ce(N__38057),
            .sr(N__49403));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_8_3  (
            .in0(N__38183),
            .in1(N__39198),
            .in2(_gnd_net_),
            .in3(N__38189),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__50290),
            .ce(N__38057),
            .sr(N__49403));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_8_4  (
            .in0(N__38176),
            .in1(N__38833),
            .in2(_gnd_net_),
            .in3(N__38186),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__50290),
            .ce(N__38057),
            .sr(N__49403));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_8_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_8_5  (
            .in0(N__39217),
            .in1(N__38177),
            .in2(_gnd_net_),
            .in3(N__38060),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50290),
            .ce(N__38057),
            .sr(N__49403));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__43861),
            .in2(N__38566),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__50278),
            .ce(N__43792),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__38536),
            .in2(N__43838),
            .in3(N__38009),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__50278),
            .ce(N__43792),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(N__38567),
            .in2(N__38479),
            .in3(N__38540),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__50278),
            .ce(N__43792),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__38537),
            .in2(N__38452),
            .in3(N__38483),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__50278),
            .ce(N__43792),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__38425),
            .in2(N__38480),
            .in3(N__38456),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__50278),
            .ce(N__43792),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__38365),
            .in2(N__38453),
            .in3(N__38429),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__50278),
            .ce(N__43792),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__38426),
            .in2(N__38314),
            .in3(N__38369),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__50278),
            .ce(N__43792),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(N__38366),
            .in2(N__38251),
            .in3(N__38318),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__50278),
            .ce(N__43792),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__38218),
            .in2(N__38315),
            .in3(N__38255),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__50265),
            .ce(N__43801),
            .sr(N__49414));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__38779),
            .in2(N__38252),
            .in3(N__38222),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__50265),
            .ce(N__43801),
            .sr(N__49414));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__38219),
            .in2(N__38755),
            .in3(N__38783),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__50265),
            .ce(N__43801),
            .sr(N__49414));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__38780),
            .in2(N__38728),
            .in3(N__38759),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__50265),
            .ce(N__43801),
            .sr(N__49414));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(N__38701),
            .in2(N__38756),
            .in3(N__38732),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__50265),
            .ce(N__43801),
            .sr(N__49414));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__38674),
            .in2(N__38729),
            .in3(N__38705),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__50265),
            .ce(N__43801),
            .sr(N__49414));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__38702),
            .in2(N__38651),
            .in3(N__38681),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__50265),
            .ce(N__43801),
            .sr(N__49414));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(N__38617),
            .in2(N__38678),
            .in3(N__38654),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__50265),
            .ce(N__43801),
            .sr(N__49414));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__38650),
            .in2(N__38593),
            .in3(N__38624),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__50256),
            .ce(N__43800),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__39049),
            .in2(N__38621),
            .in3(N__38597),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__50256),
            .ce(N__43800),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__39025),
            .in2(N__38594),
            .in3(N__38570),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__50256),
            .ce(N__43800),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__39050),
            .in2(N__39002),
            .in3(N__39032),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__50256),
            .ce(N__43800),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__38968),
            .in2(N__39029),
            .in3(N__39005),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__50256),
            .ce(N__43800),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__39001),
            .in2(N__38944),
            .in3(N__38972),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__50256),
            .ce(N__43800),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__38969),
            .in2(N__38914),
            .in3(N__38948),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__50256),
            .ce(N__43800),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__38878),
            .in2(N__38945),
            .in3(N__38918),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__50256),
            .ce(N__43800),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__38854),
            .in2(N__38915),
            .in3(N__38885),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__50244),
            .ce(N__43805),
            .sr(N__49432));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__39199),
            .in2(N__38882),
            .in3(N__38858),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__50244),
            .ce(N__43805),
            .sr(N__49432));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__38855),
            .in2(N__38837),
            .in3(N__38819),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__50244),
            .ce(N__43805),
            .sr(N__49432));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__39221),
            .in2(N__39203),
            .in3(N__39137),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__50244),
            .ce(N__43805),
            .sr(N__49432));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39134),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50244),
            .ce(N__43805),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_13_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_13_0  (
            .in0(N__39071),
            .in1(N__47048),
            .in2(N__39125),
            .in3(N__39099),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_13_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_13_1  (
            .in0(N__47047),
            .in1(N__39124),
            .in2(N__39101),
            .in3(N__39070),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_16_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_16_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_16_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_16_13_3  (
            .in0(N__48926),
            .in1(N__47209),
            .in2(_gnd_net_),
            .in3(N__47234),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50232),
            .ce(N__47864),
            .sr(N__49443));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_16_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_16_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_16_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_16_13_4  (
            .in0(N__47111),
            .in1(N__47091),
            .in2(_gnd_net_),
            .in3(N__48930),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50232),
            .ce(N__47864),
            .sr(N__49443));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_16_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_16_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_16_13_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_16_13_7  (
            .in0(N__43748),
            .in1(_gnd_net_),
            .in2(N__48937),
            .in3(N__46421),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50232),
            .ce(N__47864),
            .sr(N__49443));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43068),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_16_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_16_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41598),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_14_2 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_14_2  (
            .in0(N__42887),
            .in1(N__39904),
            .in2(N__39953),
            .in3(N__45455),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42021),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_14_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_14_4  (
            .in0(N__41518),
            .in1(N__44898),
            .in2(_gnd_net_),
            .in3(N__41472),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41517),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_14_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_14_6  (
            .in0(N__41133),
            .in1(N__45454),
            .in2(N__42909),
            .in3(N__41104),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41132),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__40916),
            .in2(N__45482),
            .in3(N__45480),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__39509),
            .in2(_gnd_net_),
            .in3(N__39233),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__39230),
            .in2(_gnd_net_),
            .in3(N__39224),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__39335),
            .in2(_gnd_net_),
            .in3(N__39329),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__39326),
            .in2(_gnd_net_),
            .in3(N__39320),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__39317),
            .in2(_gnd_net_),
            .in3(N__39311),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__39308),
            .in2(_gnd_net_),
            .in3(N__39302),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__39299),
            .in2(_gnd_net_),
            .in3(N__39293),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_16_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42923),
            .in3(N__39290),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__39287),
            .in2(_gnd_net_),
            .in3(N__39275),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__44741),
            .in2(_gnd_net_),
            .in3(N__39272),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__39269),
            .in2(_gnd_net_),
            .in3(N__39263),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(N__42047),
            .in2(_gnd_net_),
            .in3(N__39416),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(N__39413),
            .in2(_gnd_net_),
            .in3(N__39404),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(N__39401),
            .in2(_gnd_net_),
            .in3(N__39389),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_16_7  (
            .in0(_gnd_net_),
            .in1(N__39386),
            .in2(_gnd_net_),
            .in3(N__39374),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(N__41864),
            .in2(_gnd_net_),
            .in3(N__39371),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__39368),
            .in2(_gnd_net_),
            .in3(N__39359),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(N__40019),
            .in2(_gnd_net_),
            .in3(N__39356),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_17_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41684),
            .in3(N__39353),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__39350),
            .in2(_gnd_net_),
            .in3(N__39338),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__39476),
            .in2(_gnd_net_),
            .in3(N__39470),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__41903),
            .in2(_gnd_net_),
            .in3(N__39467),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(N__39500),
            .in2(_gnd_net_),
            .in3(N__39464),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(N__39461),
            .in2(_gnd_net_),
            .in3(N__39452),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__41258),
            .in2(_gnd_net_),
            .in3(N__39449),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(N__39719),
            .in2(_gnd_net_),
            .in3(N__39446),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__39674),
            .in2(_gnd_net_),
            .in3(N__39422),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__39665),
            .in2(_gnd_net_),
            .in3(N__39419),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39512),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42131),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39938),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__44732),
            .in2(N__45760),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__50184),
            .ce(N__44957),
            .sr(N__49487));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__45791),
            .in2(N__45730),
            .in3(N__39494),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__50184),
            .ce(N__44957),
            .sr(N__49487));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__45697),
            .in2(N__45761),
            .in3(N__39491),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__50184),
            .ce(N__44957),
            .sr(N__49487));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__45667),
            .in2(N__45731),
            .in3(N__39488),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__50184),
            .ce(N__44957),
            .sr(N__49487));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__45637),
            .in2(N__45701),
            .in3(N__39485),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__50184),
            .ce(N__44957),
            .sr(N__49487));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__45607),
            .in2(N__45671),
            .in3(N__39482),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__50184),
            .ce(N__44957),
            .sr(N__49487));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__45577),
            .in2(N__45641),
            .in3(N__39479),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__50184),
            .ce(N__44957),
            .sr(N__49487));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_19_7  (
            .in0(_gnd_net_),
            .in1(N__46057),
            .in2(N__45611),
            .in3(N__39539),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__50184),
            .ce(N__44957),
            .sr(N__49487));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__46024),
            .in2(N__45581),
            .in3(N__39536),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__50182),
            .ce(N__44956),
            .sr(N__49491));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(N__46000),
            .in2(N__46061),
            .in3(N__39533),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__50182),
            .ce(N__44956),
            .sr(N__49491));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__46025),
            .in2(N__45976),
            .in3(N__39530),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__50182),
            .ce(N__44956),
            .sr(N__49491));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(N__46001),
            .in2(N__45946),
            .in3(N__39527),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__50182),
            .ce(N__44956),
            .sr(N__49491));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__45916),
            .in2(N__45977),
            .in3(N__39524),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__50182),
            .ce(N__44956),
            .sr(N__49491));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(N__45889),
            .in2(N__45947),
            .in3(N__39521),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__50182),
            .ce(N__44956),
            .sr(N__49491));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__45917),
            .in2(N__45862),
            .in3(N__39518),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__50182),
            .ce(N__44956),
            .sr(N__49491));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(N__45820),
            .in2(N__45893),
            .in3(N__39515),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__50182),
            .ce(N__44956),
            .sr(N__49491));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(N__46297),
            .in2(N__45863),
            .in3(N__39566),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__50179),
            .ce(N__44955),
            .sr(N__49496));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(N__46270),
            .in2(N__45824),
            .in3(N__39563),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__50179),
            .ce(N__44955),
            .sr(N__49496));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(N__46243),
            .in2(N__46301),
            .in3(N__39560),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__50179),
            .ce(N__44955),
            .sr(N__49496));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__46271),
            .in2(N__46216),
            .in3(N__39557),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__50179),
            .ce(N__44955),
            .sr(N__49496));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__46186),
            .in2(N__46247),
            .in3(N__39554),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__50179),
            .ce(N__44955),
            .sr(N__49496));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(N__46162),
            .in2(N__46217),
            .in3(N__39551),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__50179),
            .ce(N__44955),
            .sr(N__49496));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(N__46187),
            .in2(N__46138),
            .in3(N__39548),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__50179),
            .ce(N__44955),
            .sr(N__49496));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_21_7  (
            .in0(_gnd_net_),
            .in1(N__46163),
            .in2(N__46099),
            .in3(N__39545),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__50179),
            .ce(N__44955),
            .sr(N__49496));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(N__46777),
            .in2(N__46139),
            .in3(N__39542),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__50177),
            .ce(N__44953),
            .sr(N__49498));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_22_1  (
            .in0(_gnd_net_),
            .in1(N__46747),
            .in2(N__46100),
            .in3(N__39731),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__50177),
            .ce(N__44953),
            .sr(N__49498));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(N__46721),
            .in2(N__46781),
            .in3(N__39728),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__50177),
            .ce(N__44953),
            .sr(N__49498));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(N__46571),
            .in2(N__46751),
            .in3(N__39725),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__50177),
            .ce(N__44953),
            .sr(N__49498));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39722),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39641),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39690),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42188),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_23_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_23_0  (
            .in0(N__39642),
            .in1(N__45399),
            .in2(_gnd_net_),
            .in3(N__39623),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_23_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_23_2  (
            .in0(N__41274),
            .in1(N__45398),
            .in2(_gnd_net_),
            .in3(N__39598),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_16_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_16_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41843),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_23_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_23_4  (
            .in0(N__44929),
            .in1(N__40008),
            .in2(_gnd_net_),
            .in3(N__39979),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_23_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_23_5  (
            .in0(N__39939),
            .in1(N__44930),
            .in2(_gnd_net_),
            .in3(N__39903),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_16_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_16_23_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_16_23_6  (
            .in0(N__41209),
            .in1(N__42888),
            .in2(N__41251),
            .in3(N__45400),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_23_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_23_7  (
            .in0(N__45397),
            .in1(N__42255),
            .in2(_gnd_net_),
            .in3(N__42286),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.T23_LC_16_30_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.T23_LC_16_30_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T23_LC_16_30_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.T23_LC_16_30_6  (
            .in0(_gnd_net_),
            .in1(N__39811),
            .in2(_gnd_net_),
            .in3(N__39863),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50169),
            .ce(),
            .sr(N__49529));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_17_5_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_17_5_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_17_5_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_17_5_1  (
            .in0(N__39792),
            .in1(N__39768),
            .in2(_gnd_net_),
            .in3(N__48689),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_17_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_17_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_17_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_21_LC_17_7_0  (
            .in0(N__39800),
            .in1(N__39769),
            .in2(_gnd_net_),
            .in3(N__48827),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50311),
            .ce(N__49834),
            .sr(N__49396));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_17_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_17_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_17_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_17_7_4  (
            .in0(N__46379),
            .in1(N__43692),
            .in2(_gnd_net_),
            .in3(N__48828),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50311),
            .ce(N__49834),
            .sr(N__49396));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_17_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_17_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_17_8_0  (
            .in0(N__40035),
            .in1(N__40072),
            .in2(_gnd_net_),
            .in3(N__48674),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50301),
            .ce(N__49792),
            .sr(N__49400));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_17_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_17_8_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_17_8_1  (
            .in0(N__48673),
            .in1(N__40089),
            .in2(_gnd_net_),
            .in3(N__40120),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50301),
            .ce(N__49792),
            .sr(N__49400));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_17_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_17_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_17_8_2  (
            .in0(N__40324),
            .in1(N__40293),
            .in2(_gnd_net_),
            .in3(N__48677),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50301),
            .ce(N__49792),
            .sr(N__49400));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_17_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_17_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_17_8_3  (
            .in0(N__48672),
            .in1(N__46483),
            .in2(_gnd_net_),
            .in3(N__46335),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50301),
            .ce(N__49792),
            .sr(N__49400));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_17_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_17_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_17_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_17_8_4  (
            .in0(N__43716),
            .in1(N__46448),
            .in2(_gnd_net_),
            .in3(N__48676),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50301),
            .ce(N__49792),
            .sr(N__49400));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_17_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_17_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_17_8_6  (
            .in0(N__46413),
            .in1(N__43740),
            .in2(_gnd_net_),
            .in3(N__48675),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50301),
            .ce(N__49792),
            .sr(N__49400));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_17_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_17_9_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_17_9_0  (
            .in0(N__40093),
            .in1(N__40119),
            .in2(_gnd_net_),
            .in3(N__48667),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_17_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_17_9_1 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_17_9_1  (
            .in0(N__40358),
            .in1(N__44660),
            .in2(N__44692),
            .in3(N__40343),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_9_2  (
            .in0(N__40039),
            .in1(N__40065),
            .in2(_gnd_net_),
            .in3(N__48665),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_17_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_17_9_3 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_17_9_3  (
            .in0(N__40357),
            .in1(N__44659),
            .in2(N__44693),
            .in3(N__40342),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_9_4  (
            .in0(N__40297),
            .in1(N__40323),
            .in2(_gnd_net_),
            .in3(N__48666),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_17_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_17_9_5 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_17_9_5  (
            .in0(N__40265),
            .in1(N__40232),
            .in2(N__40220),
            .in3(N__47012),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_17_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_17_9_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_17_9_6  (
            .in0(N__40578),
            .in1(_gnd_net_),
            .in2(N__40208),
            .in3(N__40622),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_17_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_17_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__40193),
            .in2(N__40205),
            .in3(N__44292),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_17_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_17_10_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_17_10_1  (
            .in0(N__44266),
            .in1(N__40187),
            .in2(N__40178),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_17_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_17_10_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_17_10_2  (
            .in0(N__44242),
            .in1(N__40169),
            .in2(N__40160),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_17_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_17_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__40139),
            .in2(N__40151),
            .in3(N__44227),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_17_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_17_10_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_17_10_4  (
            .in0(N__44212),
            .in1(N__40133),
            .in2(N__40508),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_17_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_17_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_17_10_5  (
            .in0(N__44197),
            .in1(N__40496),
            .in2(N__40484),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_17_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_17_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(N__47489),
            .in2(N__40472),
            .in3(N__44182),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_17_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_17_10_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_17_10_7  (
            .in0(N__44167),
            .in1(N__40463),
            .in2(N__40451),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_17_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_17_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__40439),
            .in2(N__40427),
            .in3(N__44152),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_17_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_17_11_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_17_11_1  (
            .in0(N__44407),
            .in1(N__40418),
            .in2(N__40406),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_17_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_17_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__40397),
            .in2(N__40385),
            .in3(N__44392),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_17_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_17_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__40376),
            .in2(N__40367),
            .in3(N__44378),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_17_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_17_11_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_17_11_4  (
            .in0(N__44356),
            .in1(N__40532),
            .in2(N__40547),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_17_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_17_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__47060),
            .in2(N__40526),
            .in3(N__44341),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_17_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_17_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__44012),
            .in2(N__40517),
            .in3(N__44326),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_17_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_17_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__47123),
            .in2(N__46802),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_17_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_17_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__44138),
            .in2(N__43676),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_17_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_17_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__43952),
            .in2(N__43412),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_17_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_17_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__47552),
            .in2(N__47690),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_17_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_17_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__40712),
            .in2(N__40706),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_17_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_17_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__48995),
            .in2(N__49070),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_17_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_17_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_17_12_5  (
            .in0(_gnd_net_),
            .in1(N__47408),
            .in2(N__47345),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_17_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_17_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__40736),
            .in2(N__40727),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40715),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_17_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_17_13_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_17_13_0  (
            .in0(N__44449),
            .in1(N__40556),
            .in2(N__40640),
            .in3(N__44430),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_17_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_17_13_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_17_13_1  (
            .in0(N__40555),
            .in1(N__40639),
            .in2(N__44432),
            .in3(N__44448),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_17_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_17_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_17_13_2  (
            .in0(N__48690),
            .in1(N__40670),
            .in2(_gnd_net_),
            .in3(N__40690),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(elapsed_time_ns_1_RNI36DN9_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_17_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_17_13_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_25_LC_17_13_3  (
            .in0(N__40671),
            .in1(_gnd_net_),
            .in2(N__40643),
            .in3(N__48692),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50245),
            .ce(N__49799),
            .sr(N__49433));
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_17_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_17_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_24_LC_17_13_5  (
            .in0(N__40626),
            .in1(N__40582),
            .in2(_gnd_net_),
            .in3(N__48691),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50245),
            .ce(N__49799),
            .sr(N__49433));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_17_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_17_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_17_14_1  (
            .in0(N__45790),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50233),
            .ce(N__44960),
            .sr(N__49444));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_17_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_17_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40835),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_17_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_17_14_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_17_14_3  (
            .in0(N__40836),
            .in1(N__45452),
            .in2(N__40910),
            .in3(N__40810),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_17_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_17_14_4 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_17_14_4  (
            .in0(N__40837),
            .in1(N__40809),
            .in2(_gnd_net_),
            .in3(N__44865),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_17_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_17_14_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(N__45453),
            .in2(_gnd_net_),
            .in3(N__43000),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_17_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_17_15_0 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_17_15_0  (
            .in0(N__42952),
            .in1(N__45444),
            .in2(N__40751),
            .in3(N__42880),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_17_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_17_15_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_17_15_1  (
            .in0(N__45445),
            .in1(N__42881),
            .in2(N__42953),
            .in3(N__40750),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_17_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_17_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__45446),
            .in2(_gnd_net_),
            .in3(N__42879),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_15_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_15_3  (
            .in0(N__42948),
            .in1(N__44864),
            .in2(_gnd_net_),
            .in3(N__40746),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45101),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_17_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_17_15_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_17_15_5  (
            .in0(N__45102),
            .in1(_gnd_net_),
            .in2(N__41183),
            .in3(N__44863),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45001),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50222),
            .ce(N__44958),
            .sr(N__49452));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_15_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__44731),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50222),
            .ce(N__44958),
            .sr(N__49452));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_17_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_17_16_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_17_16_0  (
            .in0(N__48150),
            .in1(N__45033),
            .in2(_gnd_net_),
            .in3(N__45076),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_17_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_17_16_1 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_17_16_1  (
            .in0(N__41566),
            .in1(N__45417),
            .in2(N__41614),
            .in3(N__42860),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_16_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_16_2  (
            .in0(N__44899),
            .in1(N__41134),
            .in2(_gnd_net_),
            .in3(N__41103),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_16_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_16_3  (
            .in0(N__41895),
            .in1(N__44903),
            .in2(_gnd_net_),
            .in3(N__41080),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_16_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_16_4  (
            .in0(N__44900),
            .in1(_gnd_net_),
            .in2(N__41059),
            .in3(N__40998),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_16_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_16_5  (
            .in0(N__40983),
            .in1(N__44902),
            .in2(_gnd_net_),
            .in3(N__40932),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_16_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_16_6  (
            .in0(N__44901),
            .in1(N__41607),
            .in2(_gnd_net_),
            .in3(N__41565),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_16_7 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_16_7  (
            .in0(N__45461),
            .in1(N__45416),
            .in2(_gnd_net_),
            .in3(N__45103),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_17_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_17_0  (
            .in0(N__42075),
            .in1(N__44909),
            .in2(_gnd_net_),
            .in3(N__41535),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_17_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_17_17_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_17_17_1  (
            .in0(N__41513),
            .in1(N__45424),
            .in2(N__42911),
            .in3(N__41479),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_17_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_17_2  (
            .in0(N__41427),
            .in1(N__44911),
            .in2(_gnd_net_),
            .in3(N__41397),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_17_3  (
            .in0(N__44908),
            .in1(N__41376),
            .in2(_gnd_net_),
            .in3(N__41337),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_17_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_17_17_4 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_17_17_4  (
            .in0(N__45425),
            .in1(N__42906),
            .in2(N__43001),
            .in3(N__45034),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41301),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_17_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_17_6  (
            .in0(N__41250),
            .in1(N__44912),
            .in2(_gnd_net_),
            .in3(N__41199),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_17_7  (
            .in0(N__44910),
            .in1(N__41958),
            .in2(_gnd_net_),
            .in3(N__41916),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43136),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41885),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_18_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_18_2  (
            .in0(N__41856),
            .in1(N__44914),
            .in2(_gnd_net_),
            .in3(N__41808),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_18_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_18_3  (
            .in0(N__44913),
            .in1(N__41781),
            .in2(_gnd_net_),
            .in3(N__41742),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_18_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_18_4  (
            .in0(N__41706),
            .in1(N__44915),
            .in2(_gnd_net_),
            .in3(N__41721),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41705),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_18_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_18_6  (
            .in0(N__41670),
            .in1(N__44916),
            .in2(_gnd_net_),
            .in3(N__41631),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_18_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_18_7  (
            .in0(N__43137),
            .in1(N__44928),
            .in2(_gnd_net_),
            .in3(N__43089),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_19_0  (
            .in0(N__44907),
            .in1(N__43055),
            .in2(_gnd_net_),
            .in3(N__43033),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_17_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_17_19_1 .LUT_INIT=16'b1111001111110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_17_19_1  (
            .in0(N__42908),
            .in1(N__45406),
            .in2(N__42996),
            .in3(N__45044),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_17_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_17_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42934),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_17_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_17_19_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_17_19_3  (
            .in0(N__42907),
            .in1(N__45405),
            .in2(N__42287),
            .in3(N__42256),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_4  (
            .in0(N__45404),
            .in1(N__42198),
            .in2(_gnd_net_),
            .in3(N__42162),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_19_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_19_5  (
            .in0(N__42132),
            .in1(N__44905),
            .in2(_gnd_net_),
            .in3(N__42108),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42065),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_19_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_19_7  (
            .in0(N__42022),
            .in1(N__44906),
            .in2(_gnd_net_),
            .in3(N__41992),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_17_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_17_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__45043),
            .in2(N__45062),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_17_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_17_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(N__48151),
            .in2(N__43211),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_17_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_17_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(N__43196),
            .in2(N__48248),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_17_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_17_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__48155),
            .in2(N__43190),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_17_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_17_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(N__43181),
            .in2(N__48249),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_17_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_17_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(N__48159),
            .in2(N__43169),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_17_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_17_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__43157),
            .in2(N__48250),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_17_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_17_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(N__48163),
            .in2(N__43148),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_17_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_17_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(N__48263),
            .in2(N__43307),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_17_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_17_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(N__43292),
            .in2(N__48337),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_17_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_17_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(N__48251),
            .in2(N__43283),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_17_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_17_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(N__44789),
            .in2(N__48334),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_17_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_17_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(N__48255),
            .in2(N__43268),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_17_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_17_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_17_21_5  (
            .in0(_gnd_net_),
            .in1(N__43253),
            .in2(N__48335),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_17_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_17_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(N__48259),
            .in2(N__43244),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_17_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_17_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(N__43232),
            .in2(N__48336),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_17_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_17_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(N__48267),
            .in2(N__43223),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_22_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_17_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_17_22_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_17_22_1  (
            .in0(_gnd_net_),
            .in1(N__43397),
            .in2(N__48338),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_17_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_17_22_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_17_22_2  (
            .in0(_gnd_net_),
            .in1(N__48271),
            .in2(N__43388),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_17_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_17_22_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_17_22_3  (
            .in0(_gnd_net_),
            .in1(N__43373),
            .in2(N__48339),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_17_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_17_22_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_17_22_4  (
            .in0(_gnd_net_),
            .in1(N__48275),
            .in2(N__43361),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_17_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_17_22_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(N__43346),
            .in2(N__48340),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_17_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_17_22_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_17_22_6  (
            .in0(_gnd_net_),
            .in1(N__48279),
            .in2(N__43337),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_17_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_17_22_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_17_22_7  (
            .in0(_gnd_net_),
            .in1(N__43325),
            .in2(N__48341),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_17_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_17_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_17_23_0  (
            .in0(_gnd_net_),
            .in1(N__48283),
            .in2(N__43316),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_17_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_17_23_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_17_23_1  (
            .in0(_gnd_net_),
            .in1(N__43661),
            .in2(N__48342),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_17_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_17_23_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_17_23_2  (
            .in0(_gnd_net_),
            .in1(N__48287),
            .in2(N__43655),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_17_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_17_23_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_17_23_3  (
            .in0(_gnd_net_),
            .in1(N__43646),
            .in2(N__48343),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_17_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_17_23_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_17_23_4  (
            .in0(_gnd_net_),
            .in1(N__48291),
            .in2(N__43640),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_17_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_17_23_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_17_23_5  (
            .in0(_gnd_net_),
            .in1(N__43622),
            .in2(N__48344),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_17_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_17_23_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_17_23_6  (
            .in0(_gnd_net_),
            .in1(N__48295),
            .in2(N__43610),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_23_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_23_7  (
            .in0(_gnd_net_),
            .in1(N__45450),
            .in2(_gnd_net_),
            .in3(N__43595),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_18_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_18_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_18_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_20_LC_18_6_4  (
            .in0(N__43881),
            .in1(N__43940),
            .in2(_gnd_net_),
            .in3(N__48829),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50320),
            .ce(N__49807),
            .sr(N__49393));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_7_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_7_0  (
            .in0(N__44479),
            .in1(N__43964),
            .in2(N__44507),
            .in3(N__43973),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_18_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_18_7_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_18_7_1  (
            .in0(N__43972),
            .in1(N__43963),
            .in2(N__44483),
            .in3(N__44506),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_18_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_18_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_18_7_4  (
            .in0(N__43885),
            .in1(N__43939),
            .in2(_gnd_net_),
            .in3(N__48826),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43865),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50312),
            .ce(N__43793),
            .sr(N__49397));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43837),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50312),
            .ce(N__43793),
            .sr(N__49397));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_18_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_18_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_18_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_18_8_5  (
            .in0(N__43744),
            .in1(N__46409),
            .in2(_gnd_net_),
            .in3(N__48651),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_18_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_18_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_18_8_6  (
            .in0(N__48652),
            .in1(N__43720),
            .in2(_gnd_net_),
            .in3(N__46459),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_18_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_18_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_18_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_18_8_7  (
            .in0(N__43696),
            .in1(N__46383),
            .in2(_gnd_net_),
            .in3(N__48653),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_9_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_9_0  (
            .in0(N__44528),
            .in1(N__44071),
            .in2(N__44552),
            .in3(N__44003),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_18_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_18_9_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_18_9_1  (
            .in0(N__44002),
            .in1(N__44527),
            .in2(N__44072),
            .in3(N__44548),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_18_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_18_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_18_9_2  (
            .in0(N__44103),
            .in1(N__48668),
            .in2(_gnd_net_),
            .in3(N__44119),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(elapsed_time_ns_1_RNI68CN9_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_18_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_18_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_18_9_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_18_9_3  (
            .in0(N__48670),
            .in1(_gnd_net_),
            .in2(N__44108),
            .in3(N__44104),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50302),
            .ce(N__49835),
            .sr(N__49401));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_18_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_18_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_18_9_6  (
            .in0(N__44060),
            .in1(N__44039),
            .in2(_gnd_net_),
            .in3(N__48671),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50302),
            .ce(N__49835),
            .sr(N__49401));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_18_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_18_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_18_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_18_9_7  (
            .in0(N__48669),
            .in1(N__47945),
            .in2(_gnd_net_),
            .in3(N__47924),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50302),
            .ce(N__49835),
            .sr(N__49401));
    defparam \phase_controller_inst1.stoper_hc.running_LC_18_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_18_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_18_10_2 .LUT_INIT=16'b1101010111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_18_10_2  (
            .in0(N__46835),
            .in1(N__47002),
            .in2(N__46957),
            .in3(N__46987),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50291),
            .ce(),
            .sr(N__49404));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_18_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_18_10_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_18_10_3  (
            .in0(_gnd_net_),
            .in1(N__46834),
            .in2(_gnd_net_),
            .in3(N__46950),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_18_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_18_10_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_18_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43994),
            .in3(N__46985),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_18_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_18_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_18_10_6  (
            .in0(_gnd_net_),
            .in1(N__46986),
            .in2(_gnd_net_),
            .in3(N__43984),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_18_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_18_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__44306),
            .in2(N__44300),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_18_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_18_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_18_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_18_11_1  (
            .in0(N__49744),
            .in1(N__44267),
            .in2(_gnd_net_),
            .in3(N__44255),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__50279),
            .ce(),
            .sr(N__49410));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_18_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_18_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_18_11_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_18_11_2  (
            .in0(N__49788),
            .in1(N__44243),
            .in2(N__44252),
            .in3(N__44231),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__50279),
            .ce(),
            .sr(N__49410));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_18_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_18_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_18_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_18_11_3  (
            .in0(N__49745),
            .in1(N__44228),
            .in2(_gnd_net_),
            .in3(N__44216),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__50279),
            .ce(),
            .sr(N__49410));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_18_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_18_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_18_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_18_11_4  (
            .in0(N__49789),
            .in1(N__44213),
            .in2(_gnd_net_),
            .in3(N__44201),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__50279),
            .ce(),
            .sr(N__49410));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_18_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_18_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_18_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_18_11_5  (
            .in0(N__49746),
            .in1(N__44198),
            .in2(_gnd_net_),
            .in3(N__44186),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__50279),
            .ce(),
            .sr(N__49410));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_18_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_18_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_18_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_18_11_6  (
            .in0(N__49790),
            .in1(N__44183),
            .in2(_gnd_net_),
            .in3(N__44171),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__50279),
            .ce(),
            .sr(N__49410));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_18_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_18_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_18_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_18_11_7  (
            .in0(N__49747),
            .in1(N__44168),
            .in2(_gnd_net_),
            .in3(N__44156),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__50279),
            .ce(),
            .sr(N__49410));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_18_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_18_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_18_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_18_12_0  (
            .in0(N__49850),
            .in1(N__44153),
            .in2(_gnd_net_),
            .in3(N__44141),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49415));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_18_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_18_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_18_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_18_12_1  (
            .in0(N__49774),
            .in1(N__44408),
            .in2(_gnd_net_),
            .in3(N__44396),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49415));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_18_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_18_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_18_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_18_12_2  (
            .in0(N__49847),
            .in1(N__44393),
            .in2(_gnd_net_),
            .in3(N__44381),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49415));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_18_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_18_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_18_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_18_12_3  (
            .in0(N__49775),
            .in1(N__44374),
            .in2(_gnd_net_),
            .in3(N__44360),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49415));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_18_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_18_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_18_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_18_12_4  (
            .in0(N__49848),
            .in1(N__44357),
            .in2(_gnd_net_),
            .in3(N__44345),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49415));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_18_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_18_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_18_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_18_12_5  (
            .in0(N__49776),
            .in1(N__44342),
            .in2(_gnd_net_),
            .in3(N__44330),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49415));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_18_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_18_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_18_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_18_12_6  (
            .in0(N__49849),
            .in1(N__44327),
            .in2(_gnd_net_),
            .in3(N__44315),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49415));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_18_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_18_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_18_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_18_12_7  (
            .in0(N__49777),
            .in1(N__47180),
            .in2(_gnd_net_),
            .in3(N__44312),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49415));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_18_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_18_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_18_13_0  (
            .in0(N__49766),
            .in1(N__47149),
            .in2(_gnd_net_),
            .in3(N__44309),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__50257),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_18_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_18_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_18_13_1  (
            .in0(N__49836),
            .in1(N__44547),
            .in2(_gnd_net_),
            .in3(N__44531),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__50257),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_18_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_18_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_18_13_2  (
            .in0(N__49767),
            .in1(N__44526),
            .in2(_gnd_net_),
            .in3(N__44510),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__50257),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_18_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_18_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_18_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_18_13_3  (
            .in0(N__49837),
            .in1(N__44502),
            .in2(_gnd_net_),
            .in3(N__44486),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__50257),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_18_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_18_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_18_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_18_13_4  (
            .in0(N__49768),
            .in1(N__44478),
            .in2(_gnd_net_),
            .in3(N__44459),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__50257),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_18_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_18_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_18_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_18_13_5  (
            .in0(N__49838),
            .in1(N__47575),
            .in2(_gnd_net_),
            .in3(N__44456),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__50257),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_18_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_18_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_18_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_18_13_6  (
            .in0(N__49769),
            .in1(N__47602),
            .in2(_gnd_net_),
            .in3(N__44453),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__50257),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_18_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_18_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_18_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_18_13_7  (
            .in0(N__49839),
            .in1(N__44450),
            .in2(_gnd_net_),
            .in3(N__44435),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__50257),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_18_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_18_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_18_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_18_14_0  (
            .in0(N__49770),
            .in1(N__44431),
            .in2(_gnd_net_),
            .in3(N__44414),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__50246),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_18_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_18_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_18_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_18_14_1  (
            .in0(N__49851),
            .in1(N__49020),
            .in2(_gnd_net_),
            .in3(N__44411),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__50246),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_18_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_18_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_18_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_18_14_2  (
            .in0(N__49771),
            .in1(N__49044),
            .in2(_gnd_net_),
            .in3(N__44702),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__50246),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_18_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_18_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_18_14_3  (
            .in0(N__49852),
            .in1(N__47373),
            .in2(_gnd_net_),
            .in3(N__44699),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__50246),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_18_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_18_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_18_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_18_14_4  (
            .in0(N__49772),
            .in1(N__47394),
            .in2(_gnd_net_),
            .in3(N__44696),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__50246),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_18_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_18_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_18_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_18_14_5  (
            .in0(N__49853),
            .in1(N__44680),
            .in2(_gnd_net_),
            .in3(N__44666),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__50246),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_18_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_18_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_18_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_18_14_6  (
            .in0(N__49773),
            .in1(N__44653),
            .in2(_gnd_net_),
            .in3(N__44663),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50246),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_15_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_15_0  (
            .in0(N__44596),
            .in1(N__47249),
            .in2(N__44624),
            .in3(N__47261),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_15_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_15_1  (
            .in0(N__47260),
            .in1(N__44623),
            .in2(N__44600),
            .in3(N__47248),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_18_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_18_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_18_15_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_28_LC_18_15_4  (
            .in0(N__48839),
            .in1(N__47305),
            .in2(_gnd_net_),
            .in3(N__47330),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50234),
            .ce(N__47865),
            .sr(N__49445));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_18_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_18_15_5 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_18_15_5  (
            .in0(N__45511),
            .in1(N__45544),
            .in2(N__45536),
            .in3(N__47032),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_18_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_18_15_6 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_18_15_6  (
            .in0(N__45545),
            .in1(N__45532),
            .in2(N__47036),
            .in3(N__45512),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_18_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_18_16_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_18_16_0  (
            .in0(N__45481),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_18_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_18_16_1 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__45418),
            .in2(N__45107),
            .in3(N__45104),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_18_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_18_16_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_18_16_3  (
            .in0(N__48333),
            .in1(N__44966),
            .in2(_gnd_net_),
            .in3(N__45058),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_18_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_18_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_18_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45002),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50223),
            .ce(N__44959),
            .sr(N__49453));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_18_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_18_16_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_18_16_6  (
            .in0(N__44775),
            .in1(N__44904),
            .in2(_gnd_net_),
            .in3(N__44811),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44774),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_18_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_18_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_18_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_18_17_0  (
            .in0(N__46693),
            .in1(N__44724),
            .in2(_gnd_net_),
            .in3(N__44705),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__50211),
            .ce(N__46551),
            .sr(N__49459));
    defparam \current_shift_inst.timer_s1.counter_1_LC_18_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_18_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_18_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_18_17_1  (
            .in0(N__46697),
            .in1(N__45783),
            .in2(_gnd_net_),
            .in3(N__45764),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__50211),
            .ce(N__46551),
            .sr(N__49459));
    defparam \current_shift_inst.timer_s1.counter_2_LC_18_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_18_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_18_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_18_17_2  (
            .in0(N__46694),
            .in1(N__45753),
            .in2(_gnd_net_),
            .in3(N__45734),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__50211),
            .ce(N__46551),
            .sr(N__49459));
    defparam \current_shift_inst.timer_s1.counter_3_LC_18_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_18_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_18_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_18_17_3  (
            .in0(N__46698),
            .in1(N__45718),
            .in2(_gnd_net_),
            .in3(N__45704),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__50211),
            .ce(N__46551),
            .sr(N__49459));
    defparam \current_shift_inst.timer_s1.counter_4_LC_18_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_18_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_18_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_18_17_4  (
            .in0(N__46695),
            .in1(N__45690),
            .in2(_gnd_net_),
            .in3(N__45674),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__50211),
            .ce(N__46551),
            .sr(N__49459));
    defparam \current_shift_inst.timer_s1.counter_5_LC_18_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_18_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_18_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_18_17_5  (
            .in0(N__46699),
            .in1(N__45660),
            .in2(_gnd_net_),
            .in3(N__45644),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__50211),
            .ce(N__46551),
            .sr(N__49459));
    defparam \current_shift_inst.timer_s1.counter_6_LC_18_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_18_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_18_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_18_17_6  (
            .in0(N__46696),
            .in1(N__45630),
            .in2(_gnd_net_),
            .in3(N__45614),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__50211),
            .ce(N__46551),
            .sr(N__49459));
    defparam \current_shift_inst.timer_s1.counter_7_LC_18_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_18_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_18_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_18_17_7  (
            .in0(N__46700),
            .in1(N__45600),
            .in2(_gnd_net_),
            .in3(N__45584),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__50211),
            .ce(N__46551),
            .sr(N__49459));
    defparam \current_shift_inst.timer_s1.counter_8_LC_18_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_18_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_18_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_18_18_0  (
            .in0(N__46664),
            .in1(N__45570),
            .in2(_gnd_net_),
            .in3(N__45548),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__50201),
            .ce(N__46552),
            .sr(N__49467));
    defparam \current_shift_inst.timer_s1.counter_9_LC_18_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_18_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_18_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_18_18_1  (
            .in0(N__46674),
            .in1(N__46050),
            .in2(_gnd_net_),
            .in3(N__46028),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__50201),
            .ce(N__46552),
            .sr(N__49467));
    defparam \current_shift_inst.timer_s1.counter_10_LC_18_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_18_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_18_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_18_18_2  (
            .in0(N__46661),
            .in1(N__46023),
            .in2(_gnd_net_),
            .in3(N__46004),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__50201),
            .ce(N__46552),
            .sr(N__49467));
    defparam \current_shift_inst.timer_s1.counter_11_LC_18_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_18_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_18_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_18_18_3  (
            .in0(N__46671),
            .in1(N__45994),
            .in2(_gnd_net_),
            .in3(N__45980),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__50201),
            .ce(N__46552),
            .sr(N__49467));
    defparam \current_shift_inst.timer_s1.counter_12_LC_18_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_18_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_18_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_18_18_4  (
            .in0(N__46662),
            .in1(N__45964),
            .in2(_gnd_net_),
            .in3(N__45950),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__50201),
            .ce(N__46552),
            .sr(N__49467));
    defparam \current_shift_inst.timer_s1.counter_13_LC_18_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_18_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_18_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_18_18_5  (
            .in0(N__46672),
            .in1(N__45934),
            .in2(_gnd_net_),
            .in3(N__45920),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__50201),
            .ce(N__46552),
            .sr(N__49467));
    defparam \current_shift_inst.timer_s1.counter_14_LC_18_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_18_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_18_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_18_18_6  (
            .in0(N__46663),
            .in1(N__45910),
            .in2(_gnd_net_),
            .in3(N__45896),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__50201),
            .ce(N__46552),
            .sr(N__49467));
    defparam \current_shift_inst.timer_s1.counter_15_LC_18_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_18_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_18_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_18_18_7  (
            .in0(N__46673),
            .in1(N__45882),
            .in2(_gnd_net_),
            .in3(N__45866),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__50201),
            .ce(N__46552),
            .sr(N__49467));
    defparam \current_shift_inst.timer_s1.counter_16_LC_18_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_18_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_18_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_18_19_0  (
            .in0(N__46657),
            .in1(N__45849),
            .in2(_gnd_net_),
            .in3(N__45827),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__50194),
            .ce(N__46553),
            .sr(N__49474));
    defparam \current_shift_inst.timer_s1.counter_17_LC_18_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_18_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_18_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_18_19_1  (
            .in0(N__46665),
            .in1(N__45813),
            .in2(_gnd_net_),
            .in3(N__46304),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__50194),
            .ce(N__46553),
            .sr(N__49474));
    defparam \current_shift_inst.timer_s1.counter_18_LC_18_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_18_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_18_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_18_19_2  (
            .in0(N__46658),
            .in1(N__46296),
            .in2(_gnd_net_),
            .in3(N__46274),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__50194),
            .ce(N__46553),
            .sr(N__49474));
    defparam \current_shift_inst.timer_s1.counter_19_LC_18_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_18_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_18_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_18_19_3  (
            .in0(N__46666),
            .in1(N__46264),
            .in2(_gnd_net_),
            .in3(N__46250),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__50194),
            .ce(N__46553),
            .sr(N__49474));
    defparam \current_shift_inst.timer_s1.counter_20_LC_18_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_18_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_18_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_18_19_4  (
            .in0(N__46659),
            .in1(N__46236),
            .in2(_gnd_net_),
            .in3(N__46220),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__50194),
            .ce(N__46553),
            .sr(N__49474));
    defparam \current_shift_inst.timer_s1.counter_21_LC_18_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_18_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_18_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_18_19_5  (
            .in0(N__46667),
            .in1(N__46204),
            .in2(_gnd_net_),
            .in3(N__46190),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__50194),
            .ce(N__46553),
            .sr(N__49474));
    defparam \current_shift_inst.timer_s1.counter_22_LC_18_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_18_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_18_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_18_19_6  (
            .in0(N__46660),
            .in1(N__46180),
            .in2(_gnd_net_),
            .in3(N__46166),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__50194),
            .ce(N__46553),
            .sr(N__49474));
    defparam \current_shift_inst.timer_s1.counter_23_LC_18_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_18_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_18_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_18_19_7  (
            .in0(N__46668),
            .in1(N__46156),
            .in2(_gnd_net_),
            .in3(N__46142),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__50194),
            .ce(N__46553),
            .sr(N__49474));
    defparam \current_shift_inst.timer_s1.counter_24_LC_18_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_18_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_18_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_18_20_0  (
            .in0(N__46653),
            .in1(N__46125),
            .in2(_gnd_net_),
            .in3(N__46103),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__50188),
            .ce(N__46544),
            .sr(N__49481));
    defparam \current_shift_inst.timer_s1.counter_25_LC_18_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_18_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_18_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_18_20_1  (
            .in0(N__46669),
            .in1(N__46086),
            .in2(_gnd_net_),
            .in3(N__46064),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__50188),
            .ce(N__46544),
            .sr(N__49481));
    defparam \current_shift_inst.timer_s1.counter_26_LC_18_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_18_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_18_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_18_20_2  (
            .in0(N__46654),
            .in1(N__46776),
            .in2(_gnd_net_),
            .in3(N__46754),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__50188),
            .ce(N__46544),
            .sr(N__49481));
    defparam \current_shift_inst.timer_s1.counter_27_LC_18_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_18_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_18_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_18_20_3  (
            .in0(N__46670),
            .in1(N__46740),
            .in2(_gnd_net_),
            .in3(N__46724),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__50188),
            .ce(N__46544),
            .sr(N__49481));
    defparam \current_shift_inst.timer_s1.counter_28_LC_18_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_18_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_18_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_18_20_4  (
            .in0(N__46655),
            .in1(N__46717),
            .in2(_gnd_net_),
            .in3(N__46703),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__50188),
            .ce(N__46544),
            .sr(N__49481));
    defparam \current_shift_inst.timer_s1.counter_29_LC_18_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_18_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_18_20_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_18_20_5  (
            .in0(N__46567),
            .in1(N__46656),
            .in2(_gnd_net_),
            .in3(N__46574),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50188),
            .ce(N__46544),
            .sr(N__49481));
    defparam \phase_controller_inst1.T12_LC_18_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.T12_LC_18_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T12_LC_18_22_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.T12_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(N__46498),
            .in2(_gnd_net_),
            .in3(N__48063),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50183),
            .ce(),
            .sr(N__49492));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_20_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_20_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_20_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_20_7_0  (
            .in0(N__46476),
            .in1(N__46339),
            .in2(_gnd_net_),
            .in3(N__48835),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_20_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_20_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_20_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_20_8_2  (
            .in0(N__46458),
            .in1(N__46414),
            .in2(N__46385),
            .in3(N__46331),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_20_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_20_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_20_9_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_20_9_0  (
            .in0(N__47944),
            .in1(N__47923),
            .in2(_gnd_net_),
            .in3(N__48759),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_20_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_20_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_20_9_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_20_9_5  (
            .in0(N__47301),
            .in1(N__48968),
            .in2(_gnd_net_),
            .in3(N__47018),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_20_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_20_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_20_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_20_9_6  (
            .in0(N__47748),
            .in1(N__47728),
            .in2(_gnd_net_),
            .in3(N__48757),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_20_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_20_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_20_9_7  (
            .in0(N__48758),
            .in1(N__47475),
            .in2(_gnd_net_),
            .in3(N__47447),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_20_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_20_10_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_20_10_1  (
            .in0(N__46821),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46851),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_20_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_20_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_20_10_4  (
            .in0(N__48859),
            .in1(N__50385),
            .in2(_gnd_net_),
            .in3(N__50355),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_20_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_20_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_20_10_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_20_10_5  (
            .in0(N__46820),
            .in1(N__47003),
            .in2(_gnd_net_),
            .in3(N__46850),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_20_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_20_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_20_11_0 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_20_11_0  (
            .in0(N__47996),
            .in1(N__46981),
            .in2(N__46833),
            .in3(N__46958),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50303),
            .ce(),
            .sr(N__49411));
    defparam \phase_controller_inst1.start_timer_hc_LC_20_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_20_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_20_11_2 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_20_11_2  (
            .in0(N__46930),
            .in1(N__47962),
            .in2(N__46856),
            .in3(N__46871),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50303),
            .ce(),
            .sr(N__49411));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_20_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_20_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_20_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_20_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46852),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50303),
            .ce(),
            .sr(N__49411));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_20_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_20_12_0 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_20_12_0  (
            .in0(N__47765),
            .in1(N__47178),
            .in2(N__47161),
            .in3(N__47132),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_20_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_20_12_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_20_12_1  (
            .in0(N__47825),
            .in1(N__47802),
            .in2(_gnd_net_),
            .in3(N__48862),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_20_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_20_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_20_12_2  (
            .in0(N__48861),
            .in1(N__47215),
            .in2(_gnd_net_),
            .in3(N__47227),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(elapsed_time_ns_1_RNI46CN9_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_20_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_20_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_20_12_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_20_12_3  (
            .in0(N__47216),
            .in1(_gnd_net_),
            .in2(N__47183),
            .in3(N__48863),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50292),
            .ce(N__49735),
            .sr(N__49416));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_20_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_20_12_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_20_12_4  (
            .in0(N__47764),
            .in1(N__47179),
            .in2(N__47162),
            .in3(N__47131),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_20_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_20_12_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_20_12_5  (
            .in0(N__47107),
            .in1(N__48860),
            .in2(_gnd_net_),
            .in3(N__47092),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(elapsed_time_ns_1_RNI13CN9_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_20_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_20_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_20_12_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_20_12_6  (
            .in0(N__47093),
            .in1(_gnd_net_),
            .in2(N__47063),
            .in3(N__48925),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50292),
            .ce(N__49735),
            .sr(N__49416));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_20_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_20_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_20_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_20_13_5  (
            .in0(N__47823),
            .in1(N__47803),
            .in2(_gnd_net_),
            .in3(N__48870),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50280),
            .ce(N__47870),
            .sr(N__49425));
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_20_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_20_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_20_13_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_29_LC_20_13_6  (
            .in0(N__48869),
            .in1(N__47476),
            .in2(_gnd_net_),
            .in3(N__47456),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50280),
            .ce(N__47870),
            .sr(N__49425));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_20_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_20_14_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_20_14_0  (
            .in0(N__48830),
            .in1(N__47521),
            .in2(_gnd_net_),
            .in3(N__47533),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_20_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_20_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_20_14_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_20_14_1  (
            .in0(N__47522),
            .in1(_gnd_net_),
            .in2(N__47492),
            .in3(N__48834),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50268),
            .ce(N__49734),
            .sr(N__49435));
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_20_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_20_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_20_14_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_29_LC_20_14_3  (
            .in0(N__47477),
            .in1(N__47455),
            .in2(_gnd_net_),
            .in3(N__48833),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50268),
            .ce(N__49734),
            .sr(N__49435));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_20_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_20_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_20_14_4 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_20_14_4  (
            .in0(N__47269),
            .in1(N__47395),
            .in2(N__47378),
            .in3(N__47353),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_20_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_20_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_20_14_5 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_20_14_5  (
            .in0(N__47396),
            .in1(N__47374),
            .in2(N__47357),
            .in3(N__47270),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_20_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_20_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_20_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_20_14_6  (
            .in0(N__48831),
            .in1(N__47311),
            .in2(_gnd_net_),
            .in3(N__47323),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(elapsed_time_ns_1_RNI69DN9_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_20_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_20_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_20_14_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_28_LC_20_14_7  (
            .in0(N__47312),
            .in1(_gnd_net_),
            .in2(N__47273),
            .in3(N__48832),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50268),
            .ce(N__49734),
            .sr(N__49435));
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_20_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_20_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_20_15_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_26_LC_20_15_2  (
            .in0(N__50390),
            .in1(N__50366),
            .in2(_gnd_net_),
            .in3(N__48924),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50258),
            .ce(N__47868),
            .sr(N__49446));
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_20_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_20_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_20_15_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_27_LC_20_15_7  (
            .in0(N__48923),
            .in1(N__48983),
            .in2(_gnd_net_),
            .in3(N__48467),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50258),
            .ce(N__47868),
            .sr(N__49446));
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_20_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_20_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNIE87F_2_LC_20_16_5  (
            .in0(_gnd_net_),
            .in1(N__48064),
            .in2(_gnd_net_),
            .in3(N__48000),
            .lcout(\phase_controller_inst1.state_RNIE87FZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_21_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_21_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_21_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_21_10_0  (
            .in0(N__47943),
            .in1(N__47922),
            .in2(_gnd_net_),
            .in3(N__48873),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50318),
            .ce(N__47873),
            .sr(N__49412));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_21_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_21_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_21_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_21_11_1  (
            .in0(N__47824),
            .in1(N__47807),
            .in2(_gnd_net_),
            .in3(N__48874),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50313),
            .ce(N__49803),
            .sr(N__49417));
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_21_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_21_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_21_11_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_22_LC_21_11_7  (
            .in0(N__47749),
            .in1(N__47729),
            .in2(_gnd_net_),
            .in3(N__48875),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50313),
            .ce(N__49803),
            .sr(N__49417));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_21_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_21_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_21_12_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_21_12_0  (
            .in0(N__47618),
            .in1(N__47609),
            .in2(N__47588),
            .in3(N__47561),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_21_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_21_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_21_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_21_12_2  (
            .in0(N__48857),
            .in1(N__47656),
            .in2(_gnd_net_),
            .in3(N__47668),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(elapsed_time_ns_1_RNI14DN9_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_21_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_21_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_21_12_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_23_LC_21_12_3  (
            .in0(N__47657),
            .in1(_gnd_net_),
            .in2(N__47621),
            .in3(N__48858),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50304),
            .ce(N__49733),
            .sr(N__49426));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_21_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_21_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_21_12_4 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_21_12_4  (
            .in0(N__47617),
            .in1(N__47608),
            .in2(N__47587),
            .in3(N__47560),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_21_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_21_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_21_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_27_LC_21_13_2  (
            .in0(N__48871),
            .in1(N__48978),
            .in2(_gnd_net_),
            .in3(N__48463),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50293),
            .ce(N__49804),
            .sr(N__49436));
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_21_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_21_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_21_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_26_LC_21_13_3  (
            .in0(N__50386),
            .in1(N__50362),
            .in2(_gnd_net_),
            .in3(N__48872),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50293),
            .ce(N__49804),
            .sr(N__49436));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_21_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_21_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_21_14_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_21_14_0  (
            .in0(N__49055),
            .in1(N__49046),
            .in2(N__49028),
            .in3(N__49004),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_21_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_21_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_21_14_4 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_21_14_4  (
            .in0(N__49054),
            .in1(N__49045),
            .in2(N__49027),
            .in3(N__49003),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_22_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_22_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_22_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_22_11_4  (
            .in0(N__48462),
            .in1(N__48982),
            .in2(_gnd_net_),
            .in3(N__48909),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_24_9_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_24_9_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_24_9_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_24_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // MAIN
