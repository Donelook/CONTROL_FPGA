// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 5 2025 21:16:21

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T45,
    T12,
    s4_phy,
    rgb_g,
    T01,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T45;
    output T12;
    output s4_phy;
    output rgb_g;
    output T01;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__45224;
    wire N__45223;
    wire N__45222;
    wire N__45213;
    wire N__45212;
    wire N__45211;
    wire N__45204;
    wire N__45203;
    wire N__45202;
    wire N__45195;
    wire N__45194;
    wire N__45193;
    wire N__45186;
    wire N__45185;
    wire N__45184;
    wire N__45177;
    wire N__45176;
    wire N__45175;
    wire N__45168;
    wire N__45167;
    wire N__45166;
    wire N__45159;
    wire N__45158;
    wire N__45157;
    wire N__45150;
    wire N__45149;
    wire N__45148;
    wire N__45141;
    wire N__45140;
    wire N__45139;
    wire N__45132;
    wire N__45131;
    wire N__45130;
    wire N__45123;
    wire N__45122;
    wire N__45121;
    wire N__45114;
    wire N__45113;
    wire N__45112;
    wire N__45105;
    wire N__45104;
    wire N__45103;
    wire N__45096;
    wire N__45095;
    wire N__45094;
    wire N__45087;
    wire N__45086;
    wire N__45085;
    wire N__45078;
    wire N__45077;
    wire N__45076;
    wire N__45059;
    wire N__45058;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45044;
    wire N__45041;
    wire N__45040;
    wire N__45037;
    wire N__45034;
    wire N__45031;
    wire N__45026;
    wire N__45023;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45013;
    wire N__45008;
    wire N__45005;
    wire N__45004;
    wire N__45001;
    wire N__44998;
    wire N__44995;
    wire N__44990;
    wire N__44987;
    wire N__44986;
    wire N__44983;
    wire N__44980;
    wire N__44977;
    wire N__44972;
    wire N__44969;
    wire N__44966;
    wire N__44965;
    wire N__44962;
    wire N__44959;
    wire N__44956;
    wire N__44951;
    wire N__44950;
    wire N__44949;
    wire N__44948;
    wire N__44947;
    wire N__44946;
    wire N__44945;
    wire N__44944;
    wire N__44943;
    wire N__44942;
    wire N__44941;
    wire N__44940;
    wire N__44939;
    wire N__44938;
    wire N__44937;
    wire N__44936;
    wire N__44935;
    wire N__44934;
    wire N__44933;
    wire N__44932;
    wire N__44931;
    wire N__44930;
    wire N__44929;
    wire N__44928;
    wire N__44927;
    wire N__44926;
    wire N__44925;
    wire N__44924;
    wire N__44923;
    wire N__44922;
    wire N__44921;
    wire N__44920;
    wire N__44919;
    wire N__44918;
    wire N__44917;
    wire N__44916;
    wire N__44915;
    wire N__44914;
    wire N__44913;
    wire N__44912;
    wire N__44911;
    wire N__44910;
    wire N__44909;
    wire N__44908;
    wire N__44907;
    wire N__44906;
    wire N__44905;
    wire N__44904;
    wire N__44903;
    wire N__44902;
    wire N__44901;
    wire N__44900;
    wire N__44899;
    wire N__44898;
    wire N__44897;
    wire N__44896;
    wire N__44895;
    wire N__44894;
    wire N__44893;
    wire N__44892;
    wire N__44891;
    wire N__44890;
    wire N__44889;
    wire N__44888;
    wire N__44887;
    wire N__44886;
    wire N__44885;
    wire N__44884;
    wire N__44883;
    wire N__44882;
    wire N__44881;
    wire N__44880;
    wire N__44879;
    wire N__44878;
    wire N__44877;
    wire N__44876;
    wire N__44875;
    wire N__44874;
    wire N__44873;
    wire N__44872;
    wire N__44871;
    wire N__44870;
    wire N__44869;
    wire N__44868;
    wire N__44867;
    wire N__44866;
    wire N__44865;
    wire N__44864;
    wire N__44863;
    wire N__44862;
    wire N__44861;
    wire N__44860;
    wire N__44859;
    wire N__44858;
    wire N__44857;
    wire N__44856;
    wire N__44855;
    wire N__44854;
    wire N__44853;
    wire N__44852;
    wire N__44851;
    wire N__44850;
    wire N__44849;
    wire N__44848;
    wire N__44847;
    wire N__44846;
    wire N__44845;
    wire N__44844;
    wire N__44843;
    wire N__44842;
    wire N__44841;
    wire N__44840;
    wire N__44839;
    wire N__44838;
    wire N__44837;
    wire N__44836;
    wire N__44835;
    wire N__44834;
    wire N__44833;
    wire N__44832;
    wire N__44591;
    wire N__44588;
    wire N__44587;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44577;
    wire N__44576;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44561;
    wire N__44556;
    wire N__44553;
    wire N__44546;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44531;
    wire N__44528;
    wire N__44527;
    wire N__44524;
    wire N__44521;
    wire N__44518;
    wire N__44513;
    wire N__44510;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44500;
    wire N__44495;
    wire N__44492;
    wire N__44491;
    wire N__44488;
    wire N__44485;
    wire N__44482;
    wire N__44477;
    wire N__44474;
    wire N__44473;
    wire N__44470;
    wire N__44467;
    wire N__44464;
    wire N__44459;
    wire N__44456;
    wire N__44455;
    wire N__44452;
    wire N__44449;
    wire N__44446;
    wire N__44441;
    wire N__44438;
    wire N__44437;
    wire N__44434;
    wire N__44431;
    wire N__44428;
    wire N__44423;
    wire N__44420;
    wire N__44419;
    wire N__44416;
    wire N__44413;
    wire N__44410;
    wire N__44405;
    wire N__44402;
    wire N__44401;
    wire N__44398;
    wire N__44395;
    wire N__44392;
    wire N__44387;
    wire N__44384;
    wire N__44381;
    wire N__44380;
    wire N__44379;
    wire N__44378;
    wire N__44371;
    wire N__44368;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44357;
    wire N__44354;
    wire N__44351;
    wire N__44346;
    wire N__44339;
    wire N__44338;
    wire N__44337;
    wire N__44336;
    wire N__44335;
    wire N__44334;
    wire N__44333;
    wire N__44332;
    wire N__44331;
    wire N__44328;
    wire N__44327;
    wire N__44326;
    wire N__44323;
    wire N__44322;
    wire N__44321;
    wire N__44320;
    wire N__44319;
    wire N__44318;
    wire N__44317;
    wire N__44316;
    wire N__44315;
    wire N__44314;
    wire N__44313;
    wire N__44312;
    wire N__44311;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44296;
    wire N__44293;
    wire N__44290;
    wire N__44285;
    wire N__44282;
    wire N__44275;
    wire N__44272;
    wire N__44267;
    wire N__44262;
    wire N__44259;
    wire N__44254;
    wire N__44249;
    wire N__44246;
    wire N__44243;
    wire N__44240;
    wire N__44239;
    wire N__44238;
    wire N__44235;
    wire N__44234;
    wire N__44233;
    wire N__44232;
    wire N__44231;
    wire N__44230;
    wire N__44229;
    wire N__44228;
    wire N__44227;
    wire N__44226;
    wire N__44225;
    wire N__44224;
    wire N__44223;
    wire N__44222;
    wire N__44221;
    wire N__44220;
    wire N__44219;
    wire N__44218;
    wire N__44217;
    wire N__44216;
    wire N__44215;
    wire N__44214;
    wire N__44211;
    wire N__44210;
    wire N__44209;
    wire N__44208;
    wire N__44205;
    wire N__44202;
    wire N__44201;
    wire N__44200;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44190;
    wire N__44189;
    wire N__44188;
    wire N__44187;
    wire N__44186;
    wire N__44185;
    wire N__44184;
    wire N__44183;
    wire N__44182;
    wire N__44181;
    wire N__44180;
    wire N__44179;
    wire N__44178;
    wire N__44177;
    wire N__44176;
    wire N__44175;
    wire N__44174;
    wire N__44173;
    wire N__44172;
    wire N__44171;
    wire N__44170;
    wire N__44169;
    wire N__44168;
    wire N__44165;
    wire N__44164;
    wire N__44163;
    wire N__44162;
    wire N__44161;
    wire N__44160;
    wire N__44159;
    wire N__44158;
    wire N__44157;
    wire N__44154;
    wire N__44153;
    wire N__44152;
    wire N__44151;
    wire N__44150;
    wire N__44147;
    wire N__44146;
    wire N__44145;
    wire N__44144;
    wire N__44143;
    wire N__44140;
    wire N__44139;
    wire N__44138;
    wire N__44137;
    wire N__44136;
    wire N__44135;
    wire N__44132;
    wire N__44131;
    wire N__44130;
    wire N__44129;
    wire N__44126;
    wire N__44125;
    wire N__44124;
    wire N__44123;
    wire N__44122;
    wire N__44121;
    wire N__44120;
    wire N__44119;
    wire N__44118;
    wire N__44117;
    wire N__44116;
    wire N__44115;
    wire N__44114;
    wire N__44113;
    wire N__44112;
    wire N__44111;
    wire N__44110;
    wire N__44109;
    wire N__44108;
    wire N__44107;
    wire N__44106;
    wire N__44105;
    wire N__44104;
    wire N__44103;
    wire N__43874;
    wire N__43871;
    wire N__43868;
    wire N__43865;
    wire N__43864;
    wire N__43861;
    wire N__43860;
    wire N__43857;
    wire N__43856;
    wire N__43855;
    wire N__43852;
    wire N__43843;
    wire N__43838;
    wire N__43837;
    wire N__43834;
    wire N__43833;
    wire N__43832;
    wire N__43829;
    wire N__43828;
    wire N__43827;
    wire N__43826;
    wire N__43823;
    wire N__43820;
    wire N__43819;
    wire N__43816;
    wire N__43809;
    wire N__43806;
    wire N__43803;
    wire N__43796;
    wire N__43793;
    wire N__43784;
    wire N__43781;
    wire N__43780;
    wire N__43779;
    wire N__43778;
    wire N__43777;
    wire N__43774;
    wire N__43765;
    wire N__43760;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43750;
    wire N__43745;
    wire N__43744;
    wire N__43743;
    wire N__43740;
    wire N__43737;
    wire N__43736;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43714;
    wire N__43711;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43699;
    wire N__43694;
    wire N__43691;
    wire N__43682;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43671;
    wire N__43668;
    wire N__43665;
    wire N__43662;
    wire N__43659;
    wire N__43656;
    wire N__43651;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43637;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43627;
    wire N__43622;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43610;
    wire N__43607;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43592;
    wire N__43589;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43574;
    wire N__43571;
    wire N__43568;
    wire N__43565;
    wire N__43562;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43541;
    wire N__43538;
    wire N__43535;
    wire N__43532;
    wire N__43529;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43517;
    wire N__43514;
    wire N__43511;
    wire N__43508;
    wire N__43505;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43490;
    wire N__43487;
    wire N__43484;
    wire N__43481;
    wire N__43478;
    wire N__43475;
    wire N__43472;
    wire N__43469;
    wire N__43466;
    wire N__43463;
    wire N__43460;
    wire N__43457;
    wire N__43454;
    wire N__43451;
    wire N__43448;
    wire N__43445;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43433;
    wire N__43430;
    wire N__43427;
    wire N__43424;
    wire N__43421;
    wire N__43418;
    wire N__43415;
    wire N__43412;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43394;
    wire N__43391;
    wire N__43388;
    wire N__43385;
    wire N__43382;
    wire N__43379;
    wire N__43376;
    wire N__43373;
    wire N__43370;
    wire N__43367;
    wire N__43364;
    wire N__43361;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43349;
    wire N__43346;
    wire N__43343;
    wire N__43340;
    wire N__43337;
    wire N__43334;
    wire N__43331;
    wire N__43328;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43310;
    wire N__43307;
    wire N__43304;
    wire N__43301;
    wire N__43298;
    wire N__43295;
    wire N__43292;
    wire N__43289;
    wire N__43286;
    wire N__43283;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43259;
    wire N__43256;
    wire N__43253;
    wire N__43252;
    wire N__43249;
    wire N__43246;
    wire N__43241;
    wire N__43238;
    wire N__43235;
    wire N__43232;
    wire N__43229;
    wire N__43226;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43214;
    wire N__43213;
    wire N__43210;
    wire N__43207;
    wire N__43202;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43189;
    wire N__43188;
    wire N__43185;
    wire N__43182;
    wire N__43181;
    wire N__43180;
    wire N__43179;
    wire N__43178;
    wire N__43175;
    wire N__43174;
    wire N__43171;
    wire N__43168;
    wire N__43155;
    wire N__43148;
    wire N__43145;
    wire N__43144;
    wire N__43143;
    wire N__43140;
    wire N__43139;
    wire N__43136;
    wire N__43133;
    wire N__43132;
    wire N__43131;
    wire N__43128;
    wire N__43119;
    wire N__43116;
    wire N__43111;
    wire N__43106;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43094;
    wire N__43091;
    wire N__43088;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43067;
    wire N__43064;
    wire N__43061;
    wire N__43058;
    wire N__43055;
    wire N__43052;
    wire N__43049;
    wire N__43046;
    wire N__43043;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43019;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42995;
    wire N__42992;
    wire N__42991;
    wire N__42988;
    wire N__42985;
    wire N__42980;
    wire N__42977;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42938;
    wire N__42935;
    wire N__42932;
    wire N__42929;
    wire N__42926;
    wire N__42925;
    wire N__42922;
    wire N__42919;
    wire N__42914;
    wire N__42911;
    wire N__42908;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42848;
    wire N__42845;
    wire N__42842;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42830;
    wire N__42827;
    wire N__42824;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42799;
    wire N__42796;
    wire N__42793;
    wire N__42788;
    wire N__42785;
    wire N__42782;
    wire N__42779;
    wire N__42776;
    wire N__42773;
    wire N__42770;
    wire N__42767;
    wire N__42764;
    wire N__42761;
    wire N__42760;
    wire N__42757;
    wire N__42754;
    wire N__42749;
    wire N__42746;
    wire N__42743;
    wire N__42740;
    wire N__42737;
    wire N__42734;
    wire N__42731;
    wire N__42728;
    wire N__42727;
    wire N__42724;
    wire N__42721;
    wire N__42716;
    wire N__42713;
    wire N__42710;
    wire N__42707;
    wire N__42704;
    wire N__42701;
    wire N__42698;
    wire N__42695;
    wire N__42694;
    wire N__42691;
    wire N__42688;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42674;
    wire N__42671;
    wire N__42668;
    wire N__42665;
    wire N__42662;
    wire N__42661;
    wire N__42658;
    wire N__42655;
    wire N__42650;
    wire N__42647;
    wire N__42644;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42628;
    wire N__42625;
    wire N__42622;
    wire N__42617;
    wire N__42614;
    wire N__42611;
    wire N__42608;
    wire N__42605;
    wire N__42604;
    wire N__42601;
    wire N__42598;
    wire N__42593;
    wire N__42590;
    wire N__42587;
    wire N__42584;
    wire N__42581;
    wire N__42578;
    wire N__42575;
    wire N__42572;
    wire N__42569;
    wire N__42566;
    wire N__42563;
    wire N__42560;
    wire N__42559;
    wire N__42556;
    wire N__42553;
    wire N__42548;
    wire N__42545;
    wire N__42542;
    wire N__42539;
    wire N__42536;
    wire N__42535;
    wire N__42534;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42521;
    wire N__42518;
    wire N__42515;
    wire N__42512;
    wire N__42509;
    wire N__42500;
    wire N__42499;
    wire N__42498;
    wire N__42495;
    wire N__42494;
    wire N__42489;
    wire N__42488;
    wire N__42485;
    wire N__42482;
    wire N__42479;
    wire N__42476;
    wire N__42473;
    wire N__42470;
    wire N__42467;
    wire N__42458;
    wire N__42457;
    wire N__42456;
    wire N__42455;
    wire N__42454;
    wire N__42453;
    wire N__42452;
    wire N__42451;
    wire N__42450;
    wire N__42441;
    wire N__42430;
    wire N__42429;
    wire N__42424;
    wire N__42421;
    wire N__42418;
    wire N__42413;
    wire N__42412;
    wire N__42409;
    wire N__42406;
    wire N__42403;
    wire N__42400;
    wire N__42397;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42380;
    wire N__42379;
    wire N__42376;
    wire N__42373;
    wire N__42372;
    wire N__42371;
    wire N__42366;
    wire N__42365;
    wire N__42362;
    wire N__42359;
    wire N__42356;
    wire N__42351;
    wire N__42344;
    wire N__42343;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42330;
    wire N__42325;
    wire N__42324;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42312;
    wire N__42305;
    wire N__42304;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42290;
    wire N__42289;
    wire N__42286;
    wire N__42281;
    wire N__42276;
    wire N__42269;
    wire N__42268;
    wire N__42267;
    wire N__42266;
    wire N__42265;
    wire N__42264;
    wire N__42261;
    wire N__42260;
    wire N__42257;
    wire N__42256;
    wire N__42253;
    wire N__42252;
    wire N__42251;
    wire N__42250;
    wire N__42249;
    wire N__42248;
    wire N__42247;
    wire N__42246;
    wire N__42245;
    wire N__42244;
    wire N__42233;
    wire N__42228;
    wire N__42227;
    wire N__42222;
    wire N__42215;
    wire N__42204;
    wire N__42199;
    wire N__42198;
    wire N__42197;
    wire N__42196;
    wire N__42195;
    wire N__42194;
    wire N__42191;
    wire N__42190;
    wire N__42189;
    wire N__42188;
    wire N__42187;
    wire N__42186;
    wire N__42185;
    wire N__42184;
    wire N__42183;
    wire N__42182;
    wire N__42181;
    wire N__42180;
    wire N__42179;
    wire N__42176;
    wire N__42171;
    wire N__42168;
    wire N__42167;
    wire N__42166;
    wire N__42165;
    wire N__42158;
    wire N__42141;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42117;
    wire N__42114;
    wire N__42109;
    wire N__42092;
    wire N__42091;
    wire N__42090;
    wire N__42089;
    wire N__42088;
    wire N__42087;
    wire N__42086;
    wire N__42085;
    wire N__42082;
    wire N__42079;
    wire N__42076;
    wire N__42075;
    wire N__42074;
    wire N__42073;
    wire N__42072;
    wire N__42071;
    wire N__42070;
    wire N__42069;
    wire N__42068;
    wire N__42067;
    wire N__42066;
    wire N__42063;
    wire N__42062;
    wire N__42061;
    wire N__42060;
    wire N__42043;
    wire N__42042;
    wire N__42039;
    wire N__42038;
    wire N__42029;
    wire N__42026;
    wire N__42025;
    wire N__42010;
    wire N__42009;
    wire N__42008;
    wire N__42007;
    wire N__42006;
    wire N__42003;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41987;
    wire N__41984;
    wire N__41981;
    wire N__41978;
    wire N__41973;
    wire N__41970;
    wire N__41961;
    wire N__41952;
    wire N__41945;
    wire N__41942;
    wire N__41941;
    wire N__41938;
    wire N__41935;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41911;
    wire N__41906;
    wire N__41903;
    wire N__41900;
    wire N__41897;
    wire N__41894;
    wire N__41891;
    wire N__41888;
    wire N__41885;
    wire N__41882;
    wire N__41881;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41871;
    wire N__41866;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41852;
    wire N__41849;
    wire N__41848;
    wire N__41845;
    wire N__41842;
    wire N__41837;
    wire N__41834;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41819;
    wire N__41816;
    wire N__41815;
    wire N__41814;
    wire N__41813;
    wire N__41812;
    wire N__41811;
    wire N__41810;
    wire N__41809;
    wire N__41808;
    wire N__41807;
    wire N__41806;
    wire N__41805;
    wire N__41804;
    wire N__41803;
    wire N__41802;
    wire N__41801;
    wire N__41800;
    wire N__41799;
    wire N__41798;
    wire N__41797;
    wire N__41796;
    wire N__41795;
    wire N__41794;
    wire N__41793;
    wire N__41792;
    wire N__41791;
    wire N__41790;
    wire N__41789;
    wire N__41788;
    wire N__41787;
    wire N__41778;
    wire N__41769;
    wire N__41764;
    wire N__41755;
    wire N__41746;
    wire N__41737;
    wire N__41728;
    wire N__41719;
    wire N__41714;
    wire N__41711;
    wire N__41704;
    wire N__41699;
    wire N__41696;
    wire N__41693;
    wire N__41686;
    wire N__41681;
    wire N__41678;
    wire N__41675;
    wire N__41672;
    wire N__41671;
    wire N__41668;
    wire N__41665;
    wire N__41662;
    wire N__41657;
    wire N__41656;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41646;
    wire N__41645;
    wire N__41642;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41618;
    wire N__41615;
    wire N__41612;
    wire N__41609;
    wire N__41600;
    wire N__41597;
    wire N__41596;
    wire N__41593;
    wire N__41592;
    wire N__41589;
    wire N__41586;
    wire N__41585;
    wire N__41582;
    wire N__41577;
    wire N__41574;
    wire N__41567;
    wire N__41566;
    wire N__41563;
    wire N__41560;
    wire N__41557;
    wire N__41554;
    wire N__41553;
    wire N__41552;
    wire N__41551;
    wire N__41548;
    wire N__41545;
    wire N__41540;
    wire N__41537;
    wire N__41528;
    wire N__41527;
    wire N__41524;
    wire N__41521;
    wire N__41518;
    wire N__41517;
    wire N__41512;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41502;
    wire N__41495;
    wire N__41492;
    wire N__41491;
    wire N__41488;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41478;
    wire N__41473;
    wire N__41468;
    wire N__41465;
    wire N__41464;
    wire N__41463;
    wire N__41458;
    wire N__41455;
    wire N__41452;
    wire N__41447;
    wire N__41444;
    wire N__41443;
    wire N__41440;
    wire N__41437;
    wire N__41436;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41420;
    wire N__41417;
    wire N__41416;
    wire N__41413;
    wire N__41410;
    wire N__41409;
    wire N__41406;
    wire N__41403;
    wire N__41400;
    wire N__41395;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41383;
    wire N__41380;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41365;
    wire N__41362;
    wire N__41357;
    wire N__41354;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41346;
    wire N__41341;
    wire N__41338;
    wire N__41335;
    wire N__41330;
    wire N__41327;
    wire N__41326;
    wire N__41325;
    wire N__41320;
    wire N__41317;
    wire N__41314;
    wire N__41309;
    wire N__41306;
    wire N__41303;
    wire N__41302;
    wire N__41299;
    wire N__41296;
    wire N__41293;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41281;
    wire N__41278;
    wire N__41277;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41263;
    wire N__41258;
    wire N__41255;
    wire N__41254;
    wire N__41253;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41237;
    wire N__41234;
    wire N__41233;
    wire N__41230;
    wire N__41227;
    wire N__41226;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41210;
    wire N__41207;
    wire N__41206;
    wire N__41203;
    wire N__41200;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41185;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41170;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41157;
    wire N__41154;
    wire N__41147;
    wire N__41144;
    wire N__41143;
    wire N__41140;
    wire N__41137;
    wire N__41136;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41120;
    wire N__41117;
    wire N__41116;
    wire N__41115;
    wire N__41110;
    wire N__41107;
    wire N__41104;
    wire N__41099;
    wire N__41096;
    wire N__41095;
    wire N__41092;
    wire N__41089;
    wire N__41088;
    wire N__41085;
    wire N__41082;
    wire N__41079;
    wire N__41074;
    wire N__41069;
    wire N__41066;
    wire N__41065;
    wire N__41062;
    wire N__41059;
    wire N__41058;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41044;
    wire N__41039;
    wire N__41036;
    wire N__41033;
    wire N__41032;
    wire N__41029;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41014;
    wire N__41009;
    wire N__41006;
    wire N__41005;
    wire N__41004;
    wire N__40999;
    wire N__40996;
    wire N__40993;
    wire N__40988;
    wire N__40985;
    wire N__40984;
    wire N__40981;
    wire N__40978;
    wire N__40977;
    wire N__40972;
    wire N__40969;
    wire N__40966;
    wire N__40961;
    wire N__40958;
    wire N__40957;
    wire N__40954;
    wire N__40951;
    wire N__40950;
    wire N__40947;
    wire N__40944;
    wire N__40941;
    wire N__40936;
    wire N__40931;
    wire N__40928;
    wire N__40925;
    wire N__40924;
    wire N__40921;
    wire N__40920;
    wire N__40917;
    wire N__40914;
    wire N__40911;
    wire N__40906;
    wire N__40903;
    wire N__40898;
    wire N__40895;
    wire N__40894;
    wire N__40891;
    wire N__40888;
    wire N__40887;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40871;
    wire N__40868;
    wire N__40867;
    wire N__40866;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40850;
    wire N__40847;
    wire N__40846;
    wire N__40843;
    wire N__40840;
    wire N__40839;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40825;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40800;
    wire N__40797;
    wire N__40794;
    wire N__40791;
    wire N__40788;
    wire N__40785;
    wire N__40778;
    wire N__40777;
    wire N__40774;
    wire N__40771;
    wire N__40766;
    wire N__40765;
    wire N__40762;
    wire N__40759;
    wire N__40754;
    wire N__40751;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40740;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40724;
    wire N__40721;
    wire N__40720;
    wire N__40717;
    wire N__40714;
    wire N__40713;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40697;
    wire N__40694;
    wire N__40693;
    wire N__40692;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40676;
    wire N__40673;
    wire N__40670;
    wire N__40667;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40655;
    wire N__40652;
    wire N__40649;
    wire N__40646;
    wire N__40643;
    wire N__40640;
    wire N__40637;
    wire N__40634;
    wire N__40631;
    wire N__40628;
    wire N__40625;
    wire N__40622;
    wire N__40621;
    wire N__40620;
    wire N__40619;
    wire N__40618;
    wire N__40617;
    wire N__40616;
    wire N__40615;
    wire N__40614;
    wire N__40613;
    wire N__40612;
    wire N__40611;
    wire N__40610;
    wire N__40609;
    wire N__40608;
    wire N__40607;
    wire N__40606;
    wire N__40603;
    wire N__40602;
    wire N__40599;
    wire N__40598;
    wire N__40595;
    wire N__40594;
    wire N__40591;
    wire N__40590;
    wire N__40587;
    wire N__40586;
    wire N__40583;
    wire N__40582;
    wire N__40579;
    wire N__40578;
    wire N__40577;
    wire N__40576;
    wire N__40575;
    wire N__40574;
    wire N__40573;
    wire N__40572;
    wire N__40571;
    wire N__40564;
    wire N__40561;
    wire N__40552;
    wire N__40551;
    wire N__40548;
    wire N__40547;
    wire N__40532;
    wire N__40515;
    wire N__40514;
    wire N__40511;
    wire N__40510;
    wire N__40507;
    wire N__40506;
    wire N__40503;
    wire N__40502;
    wire N__40499;
    wire N__40498;
    wire N__40495;
    wire N__40494;
    wire N__40491;
    wire N__40490;
    wire N__40487;
    wire N__40486;
    wire N__40485;
    wire N__40482;
    wire N__40477;
    wire N__40470;
    wire N__40469;
    wire N__40468;
    wire N__40467;
    wire N__40466;
    wire N__40465;
    wire N__40464;
    wire N__40463;
    wire N__40462;
    wire N__40461;
    wire N__40458;
    wire N__40455;
    wire N__40438;
    wire N__40423;
    wire N__40420;
    wire N__40413;
    wire N__40410;
    wire N__40403;
    wire N__40394;
    wire N__40391;
    wire N__40382;
    wire N__40379;
    wire N__40378;
    wire N__40377;
    wire N__40376;
    wire N__40373;
    wire N__40366;
    wire N__40363;
    wire N__40360;
    wire N__40357;
    wire N__40354;
    wire N__40351;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40339;
    wire N__40336;
    wire N__40333;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40313;
    wire N__40310;
    wire N__40307;
    wire N__40302;
    wire N__40299;
    wire N__40292;
    wire N__40289;
    wire N__40286;
    wire N__40283;
    wire N__40280;
    wire N__40279;
    wire N__40278;
    wire N__40277;
    wire N__40276;
    wire N__40275;
    wire N__40274;
    wire N__40273;
    wire N__40272;
    wire N__40271;
    wire N__40270;
    wire N__40269;
    wire N__40266;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40256;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40230;
    wire N__40229;
    wire N__40228;
    wire N__40227;
    wire N__40226;
    wire N__40225;
    wire N__40224;
    wire N__40223;
    wire N__40222;
    wire N__40221;
    wire N__40220;
    wire N__40219;
    wire N__40218;
    wire N__40207;
    wire N__40194;
    wire N__40185;
    wire N__40184;
    wire N__40183;
    wire N__40182;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40169;
    wire N__40168;
    wire N__40165;
    wire N__40164;
    wire N__40161;
    wire N__40160;
    wire N__40157;
    wire N__40156;
    wire N__40153;
    wire N__40150;
    wire N__40147;
    wire N__40144;
    wire N__40143;
    wire N__40140;
    wire N__40133;
    wire N__40126;
    wire N__40125;
    wire N__40124;
    wire N__40123;
    wire N__40122;
    wire N__40121;
    wire N__40120;
    wire N__40119;
    wire N__40118;
    wire N__40117;
    wire N__40116;
    wire N__40115;
    wire N__40114;
    wire N__40111;
    wire N__40110;
    wire N__40109;
    wire N__40108;
    wire N__40107;
    wire N__40102;
    wire N__40097;
    wire N__40080;
    wire N__40071;
    wire N__40064;
    wire N__40063;
    wire N__40062;
    wire N__40061;
    wire N__40058;
    wire N__40057;
    wire N__40052;
    wire N__40037;
    wire N__40032;
    wire N__40029;
    wire N__40020;
    wire N__40009;
    wire N__40004;
    wire N__40003;
    wire N__40000;
    wire N__39999;
    wire N__39998;
    wire N__39997;
    wire N__39996;
    wire N__39995;
    wire N__39992;
    wire N__39991;
    wire N__39988;
    wire N__39981;
    wire N__39980;
    wire N__39979;
    wire N__39978;
    wire N__39977;
    wire N__39976;
    wire N__39975;
    wire N__39974;
    wire N__39973;
    wire N__39964;
    wire N__39963;
    wire N__39962;
    wire N__39961;
    wire N__39960;
    wire N__39959;
    wire N__39958;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39940;
    wire N__39937;
    wire N__39934;
    wire N__39929;
    wire N__39926;
    wire N__39911;
    wire N__39908;
    wire N__39893;
    wire N__39886;
    wire N__39869;
    wire N__39866;
    wire N__39865;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39857;
    wire N__39854;
    wire N__39851;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39828;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39809;
    wire N__39806;
    wire N__39803;
    wire N__39800;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39788;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39764;
    wire N__39761;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39749;
    wire N__39746;
    wire N__39743;
    wire N__39740;
    wire N__39737;
    wire N__39734;
    wire N__39731;
    wire N__39728;
    wire N__39725;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39713;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39698;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39686;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39671;
    wire N__39668;
    wire N__39665;
    wire N__39664;
    wire N__39661;
    wire N__39658;
    wire N__39657;
    wire N__39652;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39605;
    wire N__39602;
    wire N__39599;
    wire N__39596;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39584;
    wire N__39581;
    wire N__39578;
    wire N__39575;
    wire N__39572;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39545;
    wire N__39542;
    wire N__39539;
    wire N__39536;
    wire N__39533;
    wire N__39530;
    wire N__39527;
    wire N__39524;
    wire N__39521;
    wire N__39518;
    wire N__39515;
    wire N__39512;
    wire N__39509;
    wire N__39506;
    wire N__39503;
    wire N__39500;
    wire N__39497;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39478;
    wire N__39473;
    wire N__39470;
    wire N__39467;
    wire N__39466;
    wire N__39463;
    wire N__39460;
    wire N__39455;
    wire N__39452;
    wire N__39451;
    wire N__39448;
    wire N__39445;
    wire N__39440;
    wire N__39437;
    wire N__39436;
    wire N__39433;
    wire N__39428;
    wire N__39425;
    wire N__39422;
    wire N__39421;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39406;
    wire N__39403;
    wire N__39400;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39388;
    wire N__39385;
    wire N__39382;
    wire N__39379;
    wire N__39376;
    wire N__39371;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39361;
    wire N__39358;
    wire N__39355;
    wire N__39350;
    wire N__39347;
    wire N__39344;
    wire N__39343;
    wire N__39342;
    wire N__39339;
    wire N__39338;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39313;
    wire N__39308;
    wire N__39303;
    wire N__39296;
    wire N__39295;
    wire N__39294;
    wire N__39293;
    wire N__39292;
    wire N__39291;
    wire N__39278;
    wire N__39275;
    wire N__39272;
    wire N__39269;
    wire N__39268;
    wire N__39265;
    wire N__39262;
    wire N__39261;
    wire N__39256;
    wire N__39253;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39239;
    wire N__39238;
    wire N__39235;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39215;
    wire N__39212;
    wire N__39209;
    wire N__39206;
    wire N__39205;
    wire N__39204;
    wire N__39201;
    wire N__39196;
    wire N__39191;
    wire N__39188;
    wire N__39185;
    wire N__39184;
    wire N__39181;
    wire N__39178;
    wire N__39177;
    wire N__39174;
    wire N__39169;
    wire N__39164;
    wire N__39161;
    wire N__39158;
    wire N__39157;
    wire N__39156;
    wire N__39153;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39119;
    wire N__39116;
    wire N__39113;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39095;
    wire N__39092;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39074;
    wire N__39071;
    wire N__39068;
    wire N__39065;
    wire N__39062;
    wire N__39061;
    wire N__39060;
    wire N__39057;
    wire N__39052;
    wire N__39047;
    wire N__39044;
    wire N__39041;
    wire N__39038;
    wire N__39037;
    wire N__39034;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39024;
    wire N__39021;
    wire N__39014;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39004;
    wire N__39001;
    wire N__39000;
    wire N__38999;
    wire N__38996;
    wire N__38993;
    wire N__38990;
    wire N__38985;
    wire N__38978;
    wire N__38975;
    wire N__38972;
    wire N__38969;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38957;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38936;
    wire N__38933;
    wire N__38930;
    wire N__38927;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38915;
    wire N__38912;
    wire N__38909;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38899;
    wire N__38896;
    wire N__38891;
    wire N__38888;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38874;
    wire N__38873;
    wire N__38870;
    wire N__38867;
    wire N__38862;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38846;
    wire N__38843;
    wire N__38840;
    wire N__38839;
    wire N__38834;
    wire N__38831;
    wire N__38830;
    wire N__38827;
    wire N__38824;
    wire N__38819;
    wire N__38818;
    wire N__38815;
    wire N__38812;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38800;
    wire N__38797;
    wire N__38794;
    wire N__38793;
    wire N__38788;
    wire N__38785;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38770;
    wire N__38767;
    wire N__38764;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38746;
    wire N__38743;
    wire N__38740;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38722;
    wire N__38717;
    wire N__38714;
    wire N__38711;
    wire N__38710;
    wire N__38707;
    wire N__38704;
    wire N__38699;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38672;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38651;
    wire N__38650;
    wire N__38647;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38620;
    wire N__38617;
    wire N__38614;
    wire N__38609;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38573;
    wire N__38572;
    wire N__38571;
    wire N__38570;
    wire N__38567;
    wire N__38562;
    wire N__38559;
    wire N__38552;
    wire N__38549;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38537;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38525;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38513;
    wire N__38512;
    wire N__38509;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38492;
    wire N__38489;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38477;
    wire N__38474;
    wire N__38473;
    wire N__38472;
    wire N__38469;
    wire N__38464;
    wire N__38459;
    wire N__38456;
    wire N__38455;
    wire N__38452;
    wire N__38449;
    wire N__38444;
    wire N__38441;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38418;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38402;
    wire N__38399;
    wire N__38396;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38384;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38357;
    wire N__38354;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38342;
    wire N__38339;
    wire N__38336;
    wire N__38333;
    wire N__38330;
    wire N__38327;
    wire N__38324;
    wire N__38321;
    wire N__38318;
    wire N__38315;
    wire N__38312;
    wire N__38309;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38295;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38279;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38267;
    wire N__38264;
    wire N__38263;
    wire N__38260;
    wire N__38259;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38242;
    wire N__38237;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38222;
    wire N__38219;
    wire N__38216;
    wire N__38213;
    wire N__38210;
    wire N__38209;
    wire N__38204;
    wire N__38203;
    wire N__38200;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38180;
    wire N__38179;
    wire N__38178;
    wire N__38177;
    wire N__38176;
    wire N__38175;
    wire N__38162;
    wire N__38159;
    wire N__38156;
    wire N__38155;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38132;
    wire N__38131;
    wire N__38126;
    wire N__38123;
    wire N__38122;
    wire N__38119;
    wire N__38118;
    wire N__38115;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38093;
    wire N__38090;
    wire N__38087;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38075;
    wire N__38074;
    wire N__38069;
    wire N__38066;
    wire N__38065;
    wire N__38060;
    wire N__38057;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38036;
    wire N__38033;
    wire N__38030;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38018;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38006;
    wire N__38003;
    wire N__38002;
    wire N__37999;
    wire N__37996;
    wire N__37991;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37979;
    wire N__37976;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37962;
    wire N__37957;
    wire N__37954;
    wire N__37949;
    wire N__37946;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37934;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37921;
    wire N__37920;
    wire N__37917;
    wire N__37914;
    wire N__37911;
    wire N__37904;
    wire N__37903;
    wire N__37900;
    wire N__37897;
    wire N__37892;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37872;
    wire N__37865;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37835;
    wire N__37834;
    wire N__37833;
    wire N__37830;
    wire N__37825;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37808;
    wire N__37807;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37778;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37766;
    wire N__37763;
    wire N__37762;
    wire N__37759;
    wire N__37758;
    wire N__37755;
    wire N__37752;
    wire N__37749;
    wire N__37742;
    wire N__37741;
    wire N__37738;
    wire N__37735;
    wire N__37730;
    wire N__37727;
    wire N__37726;
    wire N__37725;
    wire N__37724;
    wire N__37723;
    wire N__37722;
    wire N__37721;
    wire N__37720;
    wire N__37717;
    wire N__37702;
    wire N__37701;
    wire N__37700;
    wire N__37699;
    wire N__37698;
    wire N__37697;
    wire N__37696;
    wire N__37695;
    wire N__37694;
    wire N__37693;
    wire N__37688;
    wire N__37673;
    wire N__37668;
    wire N__37661;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37634;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37622;
    wire N__37621;
    wire N__37620;
    wire N__37619;
    wire N__37618;
    wire N__37617;
    wire N__37616;
    wire N__37609;
    wire N__37606;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37592;
    wire N__37591;
    wire N__37590;
    wire N__37589;
    wire N__37588;
    wire N__37587;
    wire N__37586;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37562;
    wire N__37557;
    wire N__37544;
    wire N__37541;
    wire N__37540;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37530;
    wire N__37527;
    wire N__37524;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37502;
    wire N__37499;
    wire N__37498;
    wire N__37497;
    wire N__37494;
    wire N__37493;
    wire N__37492;
    wire N__37489;
    wire N__37488;
    wire N__37485;
    wire N__37482;
    wire N__37479;
    wire N__37474;
    wire N__37469;
    wire N__37466;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37450;
    wire N__37449;
    wire N__37446;
    wire N__37441;
    wire N__37436;
    wire N__37435;
    wire N__37432;
    wire N__37429;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37411;
    wire N__37408;
    wire N__37405;
    wire N__37400;
    wire N__37399;
    wire N__37396;
    wire N__37393;
    wire N__37388;
    wire N__37387;
    wire N__37384;
    wire N__37381;
    wire N__37376;
    wire N__37375;
    wire N__37372;
    wire N__37369;
    wire N__37364;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37352;
    wire N__37351;
    wire N__37348;
    wire N__37345;
    wire N__37340;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37332;
    wire N__37329;
    wire N__37324;
    wire N__37321;
    wire N__37318;
    wire N__37313;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37301;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37291;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37274;
    wire N__37271;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37259;
    wire N__37258;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37245;
    wire N__37240;
    wire N__37237;
    wire N__37232;
    wire N__37229;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37217;
    wire N__37216;
    wire N__37213;
    wire N__37210;
    wire N__37207;
    wire N__37204;
    wire N__37199;
    wire N__37196;
    wire N__37195;
    wire N__37192;
    wire N__37189;
    wire N__37186;
    wire N__37181;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37171;
    wire N__37170;
    wire N__37167;
    wire N__37164;
    wire N__37161;
    wire N__37154;
    wire N__37153;
    wire N__37150;
    wire N__37147;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37120;
    wire N__37117;
    wire N__37114;
    wire N__37113;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37091;
    wire N__37088;
    wire N__37087;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37079;
    wire N__37078;
    wire N__37075;
    wire N__37070;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37056;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37033;
    wire N__37030;
    wire N__37029;
    wire N__37026;
    wire N__37023;
    wire N__37022;
    wire N__37021;
    wire N__37020;
    wire N__37019;
    wire N__37018;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__37000;
    wire N__36995;
    wire N__36992;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36970;
    wire N__36969;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36956;
    wire N__36947;
    wire N__36944;
    wire N__36943;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36926;
    wire N__36923;
    wire N__36922;
    wire N__36919;
    wire N__36918;
    wire N__36917;
    wire N__36914;
    wire N__36911;
    wire N__36906;
    wire N__36899;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36872;
    wire N__36871;
    wire N__36868;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36858;
    wire N__36855;
    wire N__36852;
    wire N__36849;
    wire N__36842;
    wire N__36841;
    wire N__36838;
    wire N__36837;
    wire N__36836;
    wire N__36833;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36815;
    wire N__36814;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36794;
    wire N__36789;
    wire N__36786;
    wire N__36783;
    wire N__36776;
    wire N__36775;
    wire N__36774;
    wire N__36771;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36751;
    wire N__36748;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36728;
    wire N__36725;
    wire N__36724;
    wire N__36719;
    wire N__36716;
    wire N__36715;
    wire N__36714;
    wire N__36711;
    wire N__36706;
    wire N__36703;
    wire N__36698;
    wire N__36697;
    wire N__36696;
    wire N__36693;
    wire N__36692;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36674;
    wire N__36673;
    wire N__36672;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36631;
    wire N__36630;
    wire N__36627;
    wire N__36624;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36614;
    wire N__36611;
    wire N__36606;
    wire N__36603;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36589;
    wire N__36588;
    wire N__36585;
    wire N__36580;
    wire N__36577;
    wire N__36572;
    wire N__36569;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36553;
    wire N__36550;
    wire N__36549;
    wire N__36548;
    wire N__36547;
    wire N__36544;
    wire N__36543;
    wire N__36542;
    wire N__36541;
    wire N__36540;
    wire N__36539;
    wire N__36534;
    wire N__36531;
    wire N__36530;
    wire N__36529;
    wire N__36526;
    wire N__36525;
    wire N__36524;
    wire N__36521;
    wire N__36520;
    wire N__36519;
    wire N__36518;
    wire N__36517;
    wire N__36516;
    wire N__36515;
    wire N__36514;
    wire N__36513;
    wire N__36512;
    wire N__36511;
    wire N__36510;
    wire N__36509;
    wire N__36508;
    wire N__36507;
    wire N__36506;
    wire N__36503;
    wire N__36502;
    wire N__36493;
    wire N__36488;
    wire N__36485;
    wire N__36480;
    wire N__36477;
    wire N__36474;
    wire N__36471;
    wire N__36466;
    wire N__36459;
    wire N__36454;
    wire N__36443;
    wire N__36434;
    wire N__36431;
    wire N__36426;
    wire N__36421;
    wire N__36398;
    wire N__36397;
    wire N__36396;
    wire N__36393;
    wire N__36390;
    wire N__36389;
    wire N__36386;
    wire N__36385;
    wire N__36378;
    wire N__36377;
    wire N__36376;
    wire N__36371;
    wire N__36370;
    wire N__36367;
    wire N__36364;
    wire N__36363;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36348;
    wire N__36343;
    wire N__36340;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36322;
    wire N__36321;
    wire N__36318;
    wire N__36315;
    wire N__36314;
    wire N__36311;
    wire N__36310;
    wire N__36309;
    wire N__36308;
    wire N__36307;
    wire N__36304;
    wire N__36301;
    wire N__36298;
    wire N__36293;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36269;
    wire N__36266;
    wire N__36265;
    wire N__36264;
    wire N__36261;
    wire N__36256;
    wire N__36251;
    wire N__36250;
    wire N__36249;
    wire N__36244;
    wire N__36241;
    wire N__36236;
    wire N__36233;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36203;
    wire N__36200;
    wire N__36197;
    wire N__36194;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36182;
    wire N__36179;
    wire N__36178;
    wire N__36177;
    wire N__36176;
    wire N__36173;
    wire N__36172;
    wire N__36171;
    wire N__36168;
    wire N__36167;
    wire N__36164;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36156;
    wire N__36155;
    wire N__36154;
    wire N__36153;
    wire N__36152;
    wire N__36149;
    wire N__36146;
    wire N__36145;
    wire N__36144;
    wire N__36141;
    wire N__36138;
    wire N__36135;
    wire N__36130;
    wire N__36129;
    wire N__36128;
    wire N__36127;
    wire N__36126;
    wire N__36125;
    wire N__36124;
    wire N__36121;
    wire N__36114;
    wire N__36107;
    wire N__36100;
    wire N__36091;
    wire N__36088;
    wire N__36081;
    wire N__36076;
    wire N__36059;
    wire N__36056;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36044;
    wire N__36041;
    wire N__36040;
    wire N__36037;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36010;
    wire N__36009;
    wire N__36006;
    wire N__36001;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35971;
    wire N__35968;
    wire N__35965;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35920;
    wire N__35915;
    wire N__35914;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35878;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35867;
    wire N__35864;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35850;
    wire N__35845;
    wire N__35842;
    wire N__35839;
    wire N__35834;
    wire N__35833;
    wire N__35832;
    wire N__35831;
    wire N__35830;
    wire N__35829;
    wire N__35828;
    wire N__35827;
    wire N__35826;
    wire N__35825;
    wire N__35822;
    wire N__35821;
    wire N__35820;
    wire N__35819;
    wire N__35818;
    wire N__35815;
    wire N__35814;
    wire N__35813;
    wire N__35812;
    wire N__35811;
    wire N__35810;
    wire N__35801;
    wire N__35796;
    wire N__35791;
    wire N__35788;
    wire N__35779;
    wire N__35778;
    wire N__35767;
    wire N__35764;
    wire N__35763;
    wire N__35762;
    wire N__35761;
    wire N__35760;
    wire N__35759;
    wire N__35758;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35741;
    wire N__35740;
    wire N__35739;
    wire N__35738;
    wire N__35737;
    wire N__35736;
    wire N__35731;
    wire N__35718;
    wire N__35715;
    wire N__35712;
    wire N__35707;
    wire N__35694;
    wire N__35691;
    wire N__35678;
    wire N__35677;
    wire N__35676;
    wire N__35675;
    wire N__35674;
    wire N__35673;
    wire N__35672;
    wire N__35671;
    wire N__35666;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35654;
    wire N__35653;
    wire N__35652;
    wire N__35651;
    wire N__35650;
    wire N__35649;
    wire N__35648;
    wire N__35647;
    wire N__35646;
    wire N__35645;
    wire N__35644;
    wire N__35643;
    wire N__35642;
    wire N__35639;
    wire N__35636;
    wire N__35635;
    wire N__35634;
    wire N__35633;
    wire N__35632;
    wire N__35631;
    wire N__35630;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35610;
    wire N__35599;
    wire N__35590;
    wire N__35589;
    wire N__35588;
    wire N__35587;
    wire N__35586;
    wire N__35575;
    wire N__35570;
    wire N__35565;
    wire N__35562;
    wire N__35557;
    wire N__35552;
    wire N__35543;
    wire N__35538;
    wire N__35535;
    wire N__35528;
    wire N__35519;
    wire N__35518;
    wire N__35517;
    wire N__35516;
    wire N__35515;
    wire N__35514;
    wire N__35513;
    wire N__35512;
    wire N__35511;
    wire N__35510;
    wire N__35509;
    wire N__35508;
    wire N__35507;
    wire N__35506;
    wire N__35505;
    wire N__35504;
    wire N__35501;
    wire N__35498;
    wire N__35495;
    wire N__35494;
    wire N__35493;
    wire N__35492;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35476;
    wire N__35475;
    wire N__35472;
    wire N__35469;
    wire N__35466;
    wire N__35463;
    wire N__35462;
    wire N__35459;
    wire N__35446;
    wire N__35445;
    wire N__35444;
    wire N__35443;
    wire N__35440;
    wire N__35439;
    wire N__35436;
    wire N__35433;
    wire N__35432;
    wire N__35431;
    wire N__35426;
    wire N__35419;
    wire N__35410;
    wire N__35405;
    wire N__35400;
    wire N__35397;
    wire N__35388;
    wire N__35377;
    wire N__35372;
    wire N__35365;
    wire N__35360;
    wire N__35355;
    wire N__35352;
    wire N__35349;
    wire N__35346;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35329;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35307;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35286;
    wire N__35283;
    wire N__35276;
    wire N__35273;
    wire N__35272;
    wire N__35269;
    wire N__35266;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35251;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35221;
    wire N__35218;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35207;
    wire N__35206;
    wire N__35203;
    wire N__35198;
    wire N__35193;
    wire N__35188;
    wire N__35185;
    wire N__35180;
    wire N__35177;
    wire N__35174;
    wire N__35171;
    wire N__35170;
    wire N__35167;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35129;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35111;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35100;
    wire N__35099;
    wire N__35096;
    wire N__35093;
    wire N__35090;
    wire N__35087;
    wire N__35080;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35047;
    wire N__35044;
    wire N__35043;
    wire N__35042;
    wire N__35039;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35006;
    wire N__35003;
    wire N__34994;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34964;
    wire N__34963;
    wire N__34962;
    wire N__34961;
    wire N__34960;
    wire N__34959;
    wire N__34956;
    wire N__34955;
    wire N__34954;
    wire N__34953;
    wire N__34950;
    wire N__34949;
    wire N__34948;
    wire N__34947;
    wire N__34944;
    wire N__34943;
    wire N__34942;
    wire N__34939;
    wire N__34938;
    wire N__34937;
    wire N__34934;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34916;
    wire N__34915;
    wire N__34914;
    wire N__34913;
    wire N__34912;
    wire N__34909;
    wire N__34906;
    wire N__34905;
    wire N__34902;
    wire N__34901;
    wire N__34900;
    wire N__34899;
    wire N__34898;
    wire N__34897;
    wire N__34894;
    wire N__34891;
    wire N__34890;
    wire N__34887;
    wire N__34886;
    wire N__34885;
    wire N__34884;
    wire N__34883;
    wire N__34882;
    wire N__34881;
    wire N__34880;
    wire N__34879;
    wire N__34878;
    wire N__34877;
    wire N__34876;
    wire N__34875;
    wire N__34874;
    wire N__34873;
    wire N__34872;
    wire N__34869;
    wire N__34868;
    wire N__34867;
    wire N__34866;
    wire N__34865;
    wire N__34864;
    wire N__34851;
    wire N__34848;
    wire N__34839;
    wire N__34834;
    wire N__34833;
    wire N__34826;
    wire N__34823;
    wire N__34806;
    wire N__34801;
    wire N__34798;
    wire N__34787;
    wire N__34782;
    wire N__34771;
    wire N__34766;
    wire N__34763;
    wire N__34760;
    wire N__34757;
    wire N__34746;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34726;
    wire N__34711;
    wire N__34708;
    wire N__34703;
    wire N__34698;
    wire N__34691;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34645;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34631;
    wire N__34630;
    wire N__34627;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34611;
    wire N__34608;
    wire N__34601;
    wire N__34598;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34588;
    wire N__34585;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34567;
    wire N__34566;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34552;
    wire N__34549;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34528;
    wire N__34527;
    wire N__34524;
    wire N__34521;
    wire N__34518;
    wire N__34517;
    wire N__34512;
    wire N__34507;
    wire N__34504;
    wire N__34501;
    wire N__34498;
    wire N__34495;
    wire N__34490;
    wire N__34487;
    wire N__34486;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34478;
    wire N__34475;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34454;
    wire N__34453;
    wire N__34450;
    wire N__34447;
    wire N__34444;
    wire N__34441;
    wire N__34438;
    wire N__34437;
    wire N__34432;
    wire N__34429;
    wire N__34424;
    wire N__34421;
    wire N__34418;
    wire N__34415;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34397;
    wire N__34394;
    wire N__34391;
    wire N__34390;
    wire N__34387;
    wire N__34386;
    wire N__34385;
    wire N__34382;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34359;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34342;
    wire N__34341;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34331;
    wire N__34328;
    wire N__34325;
    wire N__34324;
    wire N__34321;
    wire N__34316;
    wire N__34313;
    wire N__34310;
    wire N__34307;
    wire N__34304;
    wire N__34295;
    wire N__34292;
    wire N__34289;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34229;
    wire N__34228;
    wire N__34227;
    wire N__34224;
    wire N__34223;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34202;
    wire N__34197;
    wire N__34194;
    wire N__34193;
    wire N__34188;
    wire N__34185;
    wire N__34182;
    wire N__34179;
    wire N__34172;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34145;
    wire N__34142;
    wire N__34139;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34121;
    wire N__34118;
    wire N__34115;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34100;
    wire N__34097;
    wire N__34094;
    wire N__34091;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34033;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34013;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33995;
    wire N__33992;
    wire N__33989;
    wire N__33986;
    wire N__33983;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33887;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33825;
    wire N__33822;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33799;
    wire N__33798;
    wire N__33795;
    wire N__33790;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33778;
    wire N__33777;
    wire N__33774;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33755;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33745;
    wire N__33742;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33691;
    wire N__33690;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33653;
    wire N__33650;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33614;
    wire N__33613;
    wire N__33612;
    wire N__33609;
    wire N__33604;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33551;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33516;
    wire N__33511;
    wire N__33508;
    wire N__33503;
    wire N__33500;
    wire N__33497;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33452;
    wire N__33451;
    wire N__33446;
    wire N__33443;
    wire N__33440;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33428;
    wire N__33427;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33341;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33331;
    wire N__33330;
    wire N__33327;
    wire N__33322;
    wire N__33317;
    wire N__33314;
    wire N__33311;
    wire N__33308;
    wire N__33305;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33293;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33268;
    wire N__33265;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33248;
    wire N__33245;
    wire N__33242;
    wire N__33239;
    wire N__33236;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33122;
    wire N__33119;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33059;
    wire N__33056;
    wire N__33053;
    wire N__33050;
    wire N__33047;
    wire N__33044;
    wire N__33041;
    wire N__33038;
    wire N__33035;
    wire N__33032;
    wire N__33029;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32984;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32933;
    wire N__32930;
    wire N__32927;
    wire N__32924;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32864;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32843;
    wire N__32840;
    wire N__32837;
    wire N__32834;
    wire N__32831;
    wire N__32828;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32792;
    wire N__32789;
    wire N__32786;
    wire N__32783;
    wire N__32780;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32660;
    wire N__32657;
    wire N__32654;
    wire N__32651;
    wire N__32648;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32621;
    wire N__32618;
    wire N__32617;
    wire N__32614;
    wire N__32613;
    wire N__32612;
    wire N__32609;
    wire N__32608;
    wire N__32605;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32582;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32557;
    wire N__32556;
    wire N__32553;
    wire N__32550;
    wire N__32549;
    wire N__32546;
    wire N__32543;
    wire N__32540;
    wire N__32537;
    wire N__32534;
    wire N__32533;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32510;
    wire N__32509;
    wire N__32508;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32491;
    wire N__32488;
    wire N__32483;
    wire N__32480;
    wire N__32477;
    wire N__32472;
    wire N__32465;
    wire N__32462;
    wire N__32461;
    wire N__32458;
    wire N__32455;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32443;
    wire N__32440;
    wire N__32437;
    wire N__32434;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32408;
    wire N__32407;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32380;
    wire N__32375;
    wire N__32372;
    wire N__32369;
    wire N__32366;
    wire N__32363;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32351;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32338;
    wire N__32337;
    wire N__32336;
    wire N__32333;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32316;
    wire N__32311;
    wire N__32308;
    wire N__32305;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32288;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32251;
    wire N__32248;
    wire N__32247;
    wire N__32246;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32225;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32180;
    wire N__32179;
    wire N__32178;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32056;
    wire N__32055;
    wire N__32054;
    wire N__32051;
    wire N__32050;
    wire N__32043;
    wire N__32038;
    wire N__32035;
    wire N__32030;
    wire N__32029;
    wire N__32026;
    wire N__32025;
    wire N__32024;
    wire N__32023;
    wire N__32016;
    wire N__32011;
    wire N__32008;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31958;
    wire N__31957;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31942;
    wire N__31937;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31915;
    wire N__31910;
    wire N__31907;
    wire N__31904;
    wire N__31901;
    wire N__31898;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31883;
    wire N__31880;
    wire N__31877;
    wire N__31874;
    wire N__31871;
    wire N__31868;
    wire N__31865;
    wire N__31864;
    wire N__31863;
    wire N__31860;
    wire N__31859;
    wire N__31858;
    wire N__31857;
    wire N__31856;
    wire N__31855;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31847;
    wire N__31844;
    wire N__31839;
    wire N__31836;
    wire N__31835;
    wire N__31830;
    wire N__31827;
    wire N__31820;
    wire N__31819;
    wire N__31818;
    wire N__31817;
    wire N__31816;
    wire N__31813;
    wire N__31810;
    wire N__31809;
    wire N__31808;
    wire N__31805;
    wire N__31804;
    wire N__31803;
    wire N__31802;
    wire N__31801;
    wire N__31800;
    wire N__31799;
    wire N__31796;
    wire N__31793;
    wire N__31788;
    wire N__31779;
    wire N__31778;
    wire N__31777;
    wire N__31776;
    wire N__31775;
    wire N__31774;
    wire N__31773;
    wire N__31772;
    wire N__31771;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31747;
    wire N__31742;
    wire N__31735;
    wire N__31732;
    wire N__31723;
    wire N__31714;
    wire N__31691;
    wire N__31688;
    wire N__31687;
    wire N__31684;
    wire N__31683;
    wire N__31680;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31658;
    wire N__31657;
    wire N__31654;
    wire N__31651;
    wire N__31650;
    wire N__31649;
    wire N__31646;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31638;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31621;
    wire N__31614;
    wire N__31609;
    wire N__31608;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31584;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31570;
    wire N__31567;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31528;
    wire N__31527;
    wire N__31526;
    wire N__31523;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31501;
    wire N__31498;
    wire N__31493;
    wire N__31488;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31472;
    wire N__31471;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31463;
    wire N__31462;
    wire N__31459;
    wire N__31458;
    wire N__31457;
    wire N__31456;
    wire N__31453;
    wire N__31448;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31434;
    wire N__31431;
    wire N__31428;
    wire N__31423;
    wire N__31420;
    wire N__31409;
    wire N__31408;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31293;
    wire N__31288;
    wire N__31285;
    wire N__31280;
    wire N__31277;
    wire N__31274;
    wire N__31271;
    wire N__31268;
    wire N__31267;
    wire N__31264;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31253;
    wire N__31250;
    wire N__31245;
    wire N__31242;
    wire N__31241;
    wire N__31234;
    wire N__31231;
    wire N__31226;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31216;
    wire N__31213;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31196;
    wire N__31193;
    wire N__31190;
    wire N__31187;
    wire N__31186;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31141;
    wire N__31138;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31121;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31100;
    wire N__31097;
    wire N__31096;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31067;
    wire N__31060;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31043;
    wire N__31040;
    wire N__31037;
    wire N__31034;
    wire N__31033;
    wire N__31030;
    wire N__31027;
    wire N__31022;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30995;
    wire N__30994;
    wire N__30991;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30975;
    wire N__30968;
    wire N__30967;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30947;
    wire N__30944;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30928;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30908;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30900;
    wire N__30897;
    wire N__30894;
    wire N__30893;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30880;
    wire N__30877;
    wire N__30872;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30854;
    wire N__30851;
    wire N__30848;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30826;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30809;
    wire N__30808;
    wire N__30805;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30791;
    wire N__30790;
    wire N__30787;
    wire N__30782;
    wire N__30777;
    wire N__30770;
    wire N__30769;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30739;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30703;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30686;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30671;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30643;
    wire N__30640;
    wire N__30637;
    wire N__30634;
    wire N__30631;
    wire N__30630;
    wire N__30627;
    wire N__30626;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30611;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30595;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30579;
    wire N__30572;
    wire N__30569;
    wire N__30566;
    wire N__30563;
    wire N__30560;
    wire N__30559;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30536;
    wire N__30533;
    wire N__30530;
    wire N__30529;
    wire N__30528;
    wire N__30525;
    wire N__30524;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30490;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30463;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30443;
    wire N__30440;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30421;
    wire N__30418;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30399;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30369;
    wire N__30368;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30353;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30335;
    wire N__30334;
    wire N__30331;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30287;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30277;
    wire N__30272;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30250;
    wire N__30249;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30223;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30202;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30187;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30168;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30152;
    wire N__30149;
    wire N__30148;
    wire N__30143;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30128;
    wire N__30125;
    wire N__30124;
    wire N__30123;
    wire N__30118;
    wire N__30115;
    wire N__30112;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30083;
    wire N__30080;
    wire N__30079;
    wire N__30078;
    wire N__30077;
    wire N__30076;
    wire N__30075;
    wire N__30074;
    wire N__30073;
    wire N__30072;
    wire N__30071;
    wire N__30070;
    wire N__30069;
    wire N__30060;
    wire N__30059;
    wire N__30058;
    wire N__30057;
    wire N__30056;
    wire N__30055;
    wire N__30054;
    wire N__30053;
    wire N__30052;
    wire N__30051;
    wire N__30050;
    wire N__30049;
    wire N__30048;
    wire N__30047;
    wire N__30046;
    wire N__30045;
    wire N__30044;
    wire N__30043;
    wire N__30042;
    wire N__30033;
    wire N__30024;
    wire N__30021;
    wire N__30016;
    wire N__30007;
    wire N__29998;
    wire N__29989;
    wire N__29980;
    wire N__29975;
    wire N__29960;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29950;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29936;
    wire N__29933;
    wire N__29932;
    wire N__29931;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29910;
    wire N__29907;
    wire N__29900;
    wire N__29899;
    wire N__29894;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29856;
    wire N__29851;
    wire N__29846;
    wire N__29843;
    wire N__29842;
    wire N__29839;
    wire N__29836;
    wire N__29833;
    wire N__29830;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29815;
    wire N__29810;
    wire N__29807;
    wire N__29806;
    wire N__29801;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29786;
    wire N__29783;
    wire N__29782;
    wire N__29781;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29765;
    wire N__29762;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29750;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29735;
    wire N__29732;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29720;
    wire N__29719;
    wire N__29716;
    wire N__29713;
    wire N__29710;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29698;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29683;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29664;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29648;
    wire N__29645;
    wire N__29644;
    wire N__29639;
    wire N__29638;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29614;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29555;
    wire N__29552;
    wire N__29551;
    wire N__29546;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29531;
    wire N__29528;
    wire N__29527;
    wire N__29526;
    wire N__29521;
    wire N__29518;
    wire N__29515;
    wire N__29510;
    wire N__29507;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29495;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29480;
    wire N__29477;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29465;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29455;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29436;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29413;
    wire N__29412;
    wire N__29407;
    wire N__29404;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29368;
    wire N__29367;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29351;
    wire N__29348;
    wire N__29347;
    wire N__29344;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29320;
    wire N__29317;
    wire N__29314;
    wire N__29311;
    wire N__29310;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29287;
    wire N__29284;
    wire N__29281;
    wire N__29280;
    wire N__29275;
    wire N__29272;
    wire N__29269;
    wire N__29264;
    wire N__29261;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29249;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29219;
    wire N__29216;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29136;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29117;
    wire N__29108;
    wire N__29105;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29097;
    wire N__29094;
    wire N__29091;
    wire N__29088;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29066;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29055;
    wire N__29054;
    wire N__29051;
    wire N__29048;
    wire N__29043;
    wire N__29040;
    wire N__29033;
    wire N__29032;
    wire N__29031;
    wire N__29030;
    wire N__29021;
    wire N__29020;
    wire N__29019;
    wire N__29018;
    wire N__29017;
    wire N__29016;
    wire N__29015;
    wire N__29014;
    wire N__29013;
    wire N__29012;
    wire N__29011;
    wire N__29010;
    wire N__29009;
    wire N__29008;
    wire N__29007;
    wire N__29006;
    wire N__29005;
    wire N__29004;
    wire N__29003;
    wire N__29002;
    wire N__29001;
    wire N__29000;
    wire N__28999;
    wire N__28996;
    wire N__28987;
    wire N__28978;
    wire N__28977;
    wire N__28976;
    wire N__28975;
    wire N__28974;
    wire N__28969;
    wire N__28960;
    wire N__28951;
    wire N__28942;
    wire N__28935;
    wire N__28926;
    wire N__28921;
    wire N__28918;
    wire N__28913;
    wire N__28910;
    wire N__28901;
    wire N__28898;
    wire N__28895;
    wire N__28894;
    wire N__28891;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28867;
    wire N__28864;
    wire N__28859;
    wire N__28858;
    wire N__28857;
    wire N__28856;
    wire N__28853;
    wire N__28852;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28838;
    wire N__28835;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28814;
    wire N__28813;
    wire N__28810;
    wire N__28809;
    wire N__28808;
    wire N__28805;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28797;
    wire N__28794;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28762;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28733;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28725;
    wire N__28720;
    wire N__28717;
    wire N__28714;
    wire N__28709;
    wire N__28706;
    wire N__28705;
    wire N__28702;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28692;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28663;
    wire N__28662;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28641;
    wire N__28640;
    wire N__28637;
    wire N__28632;
    wire N__28629;
    wire N__28622;
    wire N__28619;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28597;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28589;
    wire N__28580;
    wire N__28579;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28559;
    wire N__28556;
    wire N__28555;
    wire N__28554;
    wire N__28553;
    wire N__28552;
    wire N__28549;
    wire N__28540;
    wire N__28537;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28520;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28493;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28445;
    wire N__28442;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28406;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28291;
    wire N__28290;
    wire N__28287;
    wire N__28282;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28270;
    wire N__28269;
    wire N__28266;
    wire N__28261;
    wire N__28256;
    wire N__28253;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28166;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28147;
    wire N__28144;
    wire N__28141;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28129;
    wire N__28128;
    wire N__28127;
    wire N__28120;
    wire N__28117;
    wire N__28112;
    wire N__28111;
    wire N__28110;
    wire N__28109;
    wire N__28106;
    wire N__28099;
    wire N__28094;
    wire N__28091;
    wire N__28090;
    wire N__28089;
    wire N__28088;
    wire N__28083;
    wire N__28078;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28045;
    wire N__28040;
    wire N__28037;
    wire N__28036;
    wire N__28033;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28019;
    wire N__28016;
    wire N__28015;
    wire N__28012;
    wire N__28011;
    wire N__28010;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__28000;
    wire N__27995;
    wire N__27986;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27952;
    wire N__27951;
    wire N__27948;
    wire N__27943;
    wire N__27938;
    wire N__27937;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27908;
    wire N__27907;
    wire N__27906;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27895;
    wire N__27892;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27868;
    wire N__27863;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27739;
    wire N__27736;
    wire N__27733;
    wire N__27728;
    wire N__27725;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27680;
    wire N__27679;
    wire N__27676;
    wire N__27673;
    wire N__27670;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27629;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27619;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27527;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27512;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27479;
    wire N__27478;
    wire N__27475;
    wire N__27472;
    wire N__27469;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27280;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27161;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27115;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27040;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27025;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26945;
    wire N__26942;
    wire N__26939;
    wire N__26936;
    wire N__26933;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26902;
    wire N__26901;
    wire N__26898;
    wire N__26893;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26798;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26782;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26753;
    wire N__26750;
    wire N__26747;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26723;
    wire N__26720;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26701;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26666;
    wire N__26665;
    wire N__26664;
    wire N__26663;
    wire N__26660;
    wire N__26657;
    wire N__26652;
    wire N__26651;
    wire N__26650;
    wire N__26647;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26627;
    wire N__26624;
    wire N__26623;
    wire N__26622;
    wire N__26619;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26603;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26592;
    wire N__26591;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26569;
    wire N__26564;
    wire N__26559;
    wire N__26556;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26446;
    wire N__26445;
    wire N__26444;
    wire N__26441;
    wire N__26434;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26398;
    wire N__26397;
    wire N__26396;
    wire N__26395;
    wire N__26394;
    wire N__26391;
    wire N__26390;
    wire N__26389;
    wire N__26386;
    wire N__26383;
    wire N__26382;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26374;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26341;
    wire N__26340;
    wire N__26339;
    wire N__26338;
    wire N__26335;
    wire N__26334;
    wire N__26333;
    wire N__26332;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26304;
    wire N__26299;
    wire N__26290;
    wire N__26283;
    wire N__26276;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26248;
    wire N__26245;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26225;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26213;
    wire N__26210;
    wire N__26209;
    wire N__26206;
    wire N__26205;
    wire N__26204;
    wire N__26201;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26180;
    wire N__26171;
    wire N__26168;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26147;
    wire N__26144;
    wire N__26143;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26125;
    wire N__26122;
    wire N__26121;
    wire N__26120;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26077;
    wire N__26076;
    wire N__26073;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26058;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26038;
    wire N__26037;
    wire N__26036;
    wire N__26035;
    wire N__26034;
    wire N__26033;
    wire N__26032;
    wire N__26031;
    wire N__26030;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26022;
    wire N__26019;
    wire N__26016;
    wire N__26015;
    wire N__26012;
    wire N__26011;
    wire N__26010;
    wire N__26009;
    wire N__26008;
    wire N__26005;
    wire N__26004;
    wire N__26003;
    wire N__26000;
    wire N__25999;
    wire N__25998;
    wire N__25997;
    wire N__25996;
    wire N__25987;
    wire N__25982;
    wire N__25981;
    wire N__25978;
    wire N__25961;
    wire N__25944;
    wire N__25941;
    wire N__25940;
    wire N__25939;
    wire N__25938;
    wire N__25937;
    wire N__25936;
    wire N__25935;
    wire N__25934;
    wire N__25933;
    wire N__25932;
    wire N__25931;
    wire N__25930;
    wire N__25929;
    wire N__25926;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25911;
    wire N__25906;
    wire N__25893;
    wire N__25884;
    wire N__25881;
    wire N__25876;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25850;
    wire N__25847;
    wire N__25846;
    wire N__25845;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25829;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25804;
    wire N__25801;
    wire N__25800;
    wire N__25799;
    wire N__25798;
    wire N__25797;
    wire N__25796;
    wire N__25793;
    wire N__25792;
    wire N__25791;
    wire N__25790;
    wire N__25789;
    wire N__25788;
    wire N__25787;
    wire N__25786;
    wire N__25785;
    wire N__25782;
    wire N__25777;
    wire N__25766;
    wire N__25761;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25733;
    wire N__25732;
    wire N__25731;
    wire N__25730;
    wire N__25729;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25721;
    wire N__25720;
    wire N__25719;
    wire N__25716;
    wire N__25715;
    wire N__25714;
    wire N__25711;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25689;
    wire N__25686;
    wire N__25673;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25642;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25607;
    wire N__25606;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25596;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25537;
    wire N__25536;
    wire N__25533;
    wire N__25528;
    wire N__25523;
    wire N__25520;
    wire N__25519;
    wire N__25516;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25468;
    wire N__25465;
    wire N__25464;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25450;
    wire N__25449;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25437;
    wire N__25432;
    wire N__25429;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25372;
    wire N__25369;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25248;
    wire N__25245;
    wire N__25244;
    wire N__25241;
    wire N__25240;
    wire N__25239;
    wire N__25236;
    wire N__25235;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25214;
    wire N__25211;
    wire N__25202;
    wire N__25201;
    wire N__25200;
    wire N__25199;
    wire N__25196;
    wire N__25195;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25185;
    wire N__25182;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25164;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25150;
    wire N__25147;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25130;
    wire N__25127;
    wire N__25126;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25118;
    wire N__25115;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25052;
    wire N__25051;
    wire N__25046;
    wire N__25043;
    wire N__25042;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24997;
    wire N__24996;
    wire N__24995;
    wire N__24994;
    wire N__24991;
    wire N__24982;
    wire N__24977;
    wire N__24976;
    wire N__24975;
    wire N__24972;
    wire N__24971;
    wire N__24970;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24938;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24927;
    wire N__24922;
    wire N__24919;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24892;
    wire N__24891;
    wire N__24888;
    wire N__24887;
    wire N__24884;
    wire N__24883;
    wire N__24882;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24868;
    wire N__24865;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24805;
    wire N__24804;
    wire N__24801;
    wire N__24796;
    wire N__24791;
    wire N__24788;
    wire N__24787;
    wire N__24786;
    wire N__24783;
    wire N__24778;
    wire N__24773;
    wire N__24772;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24757;
    wire N__24752;
    wire N__24751;
    wire N__24750;
    wire N__24749;
    wire N__24748;
    wire N__24745;
    wire N__24744;
    wire N__24743;
    wire N__24742;
    wire N__24741;
    wire N__24740;
    wire N__24739;
    wire N__24738;
    wire N__24737;
    wire N__24728;
    wire N__24727;
    wire N__24726;
    wire N__24715;
    wire N__24710;
    wire N__24705;
    wire N__24702;
    wire N__24701;
    wire N__24700;
    wire N__24699;
    wire N__24696;
    wire N__24693;
    wire N__24692;
    wire N__24691;
    wire N__24690;
    wire N__24689;
    wire N__24688;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24674;
    wire N__24671;
    wire N__24670;
    wire N__24669;
    wire N__24668;
    wire N__24651;
    wire N__24646;
    wire N__24643;
    wire N__24638;
    wire N__24631;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24547;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24526;
    wire N__24525;
    wire N__24524;
    wire N__24523;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24511;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24495;
    wire N__24492;
    wire N__24487;
    wire N__24482;
    wire N__24481;
    wire N__24480;
    wire N__24475;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24443;
    wire N__24440;
    wire N__24439;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24418;
    wire N__24413;
    wire N__24410;
    wire N__24409;
    wire N__24408;
    wire N__24405;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24325;
    wire N__24322;
    wire N__24319;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24158;
    wire N__24155;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24109;
    wire N__24106;
    wire N__24103;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24049;
    wire N__24046;
    wire N__24043;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23771;
    wire N__23768;
    wire N__23767;
    wire N__23766;
    wire N__23763;
    wire N__23758;
    wire N__23753;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23741;
    wire N__23740;
    wire N__23739;
    wire N__23736;
    wire N__23731;
    wire N__23726;
    wire N__23723;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23713;
    wire N__23712;
    wire N__23707;
    wire N__23704;
    wire N__23699;
    wire N__23696;
    wire N__23695;
    wire N__23692;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23675;
    wire N__23674;
    wire N__23671;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23654;
    wire N__23653;
    wire N__23652;
    wire N__23651;
    wire N__23650;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23536;
    wire N__23531;
    wire N__23528;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23509;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23480;
    wire N__23477;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23465;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23446;
    wire N__23443;
    wire N__23438;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23428;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23416;
    wire N__23413;
    wire N__23412;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23401;
    wire N__23398;
    wire N__23391;
    wire N__23388;
    wire N__23381;
    wire N__23378;
    wire N__23377;
    wire N__23376;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23345;
    wire N__23342;
    wire N__23341;
    wire N__23340;
    wire N__23337;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23251;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23213;
    wire N__23210;
    wire N__23209;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23179;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23056;
    wire N__23055;
    wire N__23054;
    wire N__23053;
    wire N__23050;
    wire N__23049;
    wire N__23046;
    wire N__23045;
    wire N__23042;
    wire N__23041;
    wire N__23040;
    wire N__23039;
    wire N__23038;
    wire N__23037;
    wire N__23036;
    wire N__23035;
    wire N__23018;
    wire N__23017;
    wire N__23014;
    wire N__23013;
    wire N__23010;
    wire N__23009;
    wire N__23006;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22998;
    wire N__22995;
    wire N__22994;
    wire N__22991;
    wire N__22974;
    wire N__22965;
    wire N__22958;
    wire N__22955;
    wire N__22954;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22937;
    wire N__22934;
    wire N__22933;
    wire N__22932;
    wire N__22929;
    wire N__22924;
    wire N__22919;
    wire N__22916;
    wire N__22915;
    wire N__22914;
    wire N__22911;
    wire N__22906;
    wire N__22901;
    wire N__22898;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22871;
    wire N__22868;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22834;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22810;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22793;
    wire N__22790;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22760;
    wire N__22757;
    wire N__22756;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22739;
    wire N__22736;
    wire N__22735;
    wire N__22734;
    wire N__22731;
    wire N__22726;
    wire N__22721;
    wire N__22718;
    wire N__22717;
    wire N__22716;
    wire N__22713;
    wire N__22708;
    wire N__22703;
    wire N__22700;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22673;
    wire N__22670;
    wire N__22669;
    wire N__22666;
    wire N__22663;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22636;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22612;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22588;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22564;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22547;
    wire N__22544;
    wire N__22543;
    wire N__22542;
    wire N__22539;
    wire N__22534;
    wire N__22529;
    wire N__22526;
    wire N__22525;
    wire N__22524;
    wire N__22521;
    wire N__22516;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22478;
    wire N__22475;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22441;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22417;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22393;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22376;
    wire N__22373;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22361;
    wire N__22358;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22339;
    wire N__22338;
    wire N__22335;
    wire N__22330;
    wire N__22325;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22317;
    wire N__22314;
    wire N__22309;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22243;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22219;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22195;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22185;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22121;
    wire N__22120;
    wire N__22115;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22100;
    wire N__22099;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22075;
    wire N__22070;
    wire N__22069;
    wire N__22066;
    wire N__22065;
    wire N__22062;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22040;
    wire N__22037;
    wire N__22036;
    wire N__22035;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22015;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21934;
    wire N__21931;
    wire N__21930;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21922;
    wire N__21917;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21899;
    wire N__21896;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21888;
    wire N__21887;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21869;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21857;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21833;
    wire N__21832;
    wire N__21831;
    wire N__21830;
    wire N__21827;
    wire N__21826;
    wire N__21825;
    wire N__21824;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21816;
    wire N__21811;
    wire N__21806;
    wire N__21801;
    wire N__21796;
    wire N__21793;
    wire N__21782;
    wire N__21781;
    wire N__21778;
    wire N__21777;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21765;
    wire N__21758;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21746;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21673;
    wire N__21672;
    wire N__21671;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21663;
    wire N__21662;
    wire N__21661;
    wire N__21656;
    wire N__21653;
    wire N__21652;
    wire N__21651;
    wire N__21646;
    wire N__21643;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21627;
    wire N__21624;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21605;
    wire N__21602;
    wire N__21593;
    wire N__21590;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21578;
    wire N__21577;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21530;
    wire N__21527;
    wire N__21526;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21493;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21464;
    wire N__21461;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21398;
    wire N__21395;
    wire N__21394;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21326;
    wire N__21323;
    wire N__21322;
    wire N__21317;
    wire N__21314;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21286;
    wire N__21281;
    wire N__21278;
    wire N__21275;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21255;
    wire N__21250;
    wire N__21247;
    wire N__21242;
    wire N__21239;
    wire N__21238;
    wire N__21235;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21220;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21193;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21175;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21150;
    wire N__21145;
    wire N__21142;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21127;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21049;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21034;
    wire N__21031;
    wire N__21028;
    wire N__21023;
    wire N__21020;
    wire N__21019;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20777;
    wire N__20774;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20741;
    wire N__20740;
    wire N__20739;
    wire N__20736;
    wire N__20731;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20653;
    wire N__20652;
    wire N__20649;
    wire N__20644;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20632;
    wire N__20629;
    wire N__20628;
    wire N__20625;
    wire N__20624;
    wire N__20621;
    wire N__20614;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20554;
    wire N__20553;
    wire N__20552;
    wire N__20549;
    wire N__20548;
    wire N__20547;
    wire N__20546;
    wire N__20541;
    wire N__20538;
    wire N__20535;
    wire N__20534;
    wire N__20531;
    wire N__20526;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20499;
    wire N__20494;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20377;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20320;
    wire N__20319;
    wire N__20316;
    wire N__20315;
    wire N__20312;
    wire N__20311;
    wire N__20310;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20294;
    wire N__20291;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20279;
    wire N__20276;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20245;
    wire N__20242;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20209;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20179;
    wire N__20176;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20134;
    wire N__20131;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20101;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20053;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20017;
    wire N__20014;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19978;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19945;
    wire N__19944;
    wire N__19941;
    wire N__19936;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19867;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19816;
    wire N__19813;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19782;
    wire N__19777;
    wire N__19774;
    wire N__19769;
    wire N__19768;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19742;
    wire N__19739;
    wire N__19738;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19711;
    wire N__19706;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19643;
    wire N__19642;
    wire N__19641;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19633;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19585;
    wire N__19584;
    wire N__19583;
    wire N__19582;
    wire N__19581;
    wire N__19580;
    wire N__19579;
    wire N__19578;
    wire N__19577;
    wire N__19568;
    wire N__19563;
    wire N__19554;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19501;
    wire N__19500;
    wire N__19499;
    wire N__19498;
    wire N__19497;
    wire N__19496;
    wire N__19495;
    wire N__19494;
    wire N__19493;
    wire N__19488;
    wire N__19483;
    wire N__19480;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19450;
    wire N__19445;
    wire N__19444;
    wire N__19443;
    wire N__19442;
    wire N__19441;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19433;
    wire N__19432;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19422;
    wire N__19419;
    wire N__19418;
    wire N__19417;
    wire N__19416;
    wire N__19415;
    wire N__19414;
    wire N__19413;
    wire N__19412;
    wire N__19411;
    wire N__19406;
    wire N__19403;
    wire N__19392;
    wire N__19387;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19369;
    wire N__19366;
    wire N__19365;
    wire N__19364;
    wire N__19363;
    wire N__19362;
    wire N__19361;
    wire N__19360;
    wire N__19359;
    wire N__19358;
    wire N__19357;
    wire N__19356;
    wire N__19355;
    wire N__19354;
    wire N__19353;
    wire N__19352;
    wire N__19351;
    wire N__19346;
    wire N__19341;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19313;
    wire N__19298;
    wire N__19293;
    wire N__19288;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19264;
    wire N__19259;
    wire N__19258;
    wire N__19257;
    wire N__19256;
    wire N__19255;
    wire N__19254;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19236;
    wire N__19235;
    wire N__19234;
    wire N__19227;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19160;
    wire N__19157;
    wire N__19156;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19146;
    wire N__19141;
    wire N__19136;
    wire N__19133;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19121;
    wire N__19118;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19106;
    wire N__19103;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19073;
    wire N__19072;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19048;
    wire N__19047;
    wire N__19046;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19029;
    wire N__19028;
    wire N__19023;
    wire N__19022;
    wire N__19019;
    wire N__19018;
    wire N__19015;
    wire N__19008;
    wire N__19007;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18989;
    wire N__18984;
    wire N__18979;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18934;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18911;
    wire N__18910;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18865;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18849;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18817;
    wire N__18814;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18797;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18776;
    wire N__18773;
    wire N__18772;
    wire N__18771;
    wire N__18768;
    wire N__18763;
    wire N__18758;
    wire N__18755;
    wire N__18754;
    wire N__18751;
    wire N__18748;
    wire N__18743;
    wire N__18742;
    wire N__18741;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18640;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18589;
    wire N__18588;
    wire N__18583;
    wire N__18580;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18376;
    wire N__18375;
    wire N__18374;
    wire N__18373;
    wire N__18372;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18350;
    wire N__18345;
    wire N__18336;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18265;
    wire N__18264;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18232;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17653;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire bfn_1_9_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire bfn_1_10_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire bfn_1_11_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire N_38_i_i;
    wire rgb_drv_RNOZ0;
    wire bfn_2_8_0_;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire bfn_2_9_0_;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire bfn_2_10_0_;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire bfn_2_11_0_;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire bfn_2_12_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire pwm_duty_input_5;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_3_9_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_3_10_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire bfn_3_11_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire pwm_duty_input_3;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.N_154 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.N_16 ;
    wire N_19_1;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire bfn_4_9_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_4_10_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire pwm_duty_input_4;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ;
    wire pwm_duty_input_9;
    wire pwm_duty_input_6;
    wire pwm_duty_input_7;
    wire pwm_duty_input_8;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.N_149 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_153 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire il_max_comp2_c;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_5_9_0_;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_5_10_0_;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.N_53 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ;
    wire il_max_comp2_D1;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.N_155 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ;
    wire elapsed_time_ns_1_RNI3VBED1_0_16_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9_cascade_ ;
    wire elapsed_time_ns_1_RNIP1MD11_0_12_cascade_;
    wire elapsed_time_ns_1_RNIP1MD11_0_12;
    wire elapsed_time_ns_1_RNINVLD11_0_10_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2_cascade_ ;
    wire elapsed_time_ns_1_RNIQ2MD11_0_13;
    wire elapsed_time_ns_1_RNI51CED1_0_18_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_ ;
    wire bfn_7_18_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire bfn_7_19_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire bfn_7_20_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire bfn_7_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire il_min_comp2_c;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_8_10_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_8_11_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire bfn_8_12_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_8_13_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_f0_i_1Z0Z_9 ;
    wire elapsed_time_ns_1_RNINVLD11_0_10;
    wire \phase_controller_inst1.stoper_hc.N_315 ;
    wire elapsed_time_ns_1_RNIO0MD11_0_11;
    wire elapsed_time_ns_1_RNIR4ND11_0_23;
    wire elapsed_time_ns_1_RNIS5ND11_0_24;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14 ;
    wire elapsed_time_ns_1_RNI1TBED1_0_14;
    wire elapsed_time_ns_1_RNI1TBED1_0_14_cascade_;
    wire elapsed_time_ns_1_RNIL13KD1_0_9;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ;
    wire bfn_8_19_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_8_20_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_8_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_8_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire s4_phy_c;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire bfn_9_13_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire bfn_9_14_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire bfn_9_15_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire elapsed_time_ns_1_RNI40CED1_0_17;
    wire elapsed_time_ns_1_RNI51CED1_0_18;
    wire elapsed_time_ns_1_RNI3VBED1_0_16;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3Z0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_328 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire elapsed_time_ns_1_RNI1BND11_0_29;
    wire elapsed_time_ns_1_RNIP2ND11_0_21;
    wire elapsed_time_ns_1_RNI1BND11_0_29_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_o5_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_o5_7Z0Z_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire elapsed_time_ns_1_RNIO1ND11_0_20;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire elapsed_time_ns_1_RNIQ3ND11_0_22;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire elapsed_time_ns_1_RNIT6ND11_0_25;
    wire elapsed_time_ns_1_RNIT6ND11_0_25_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_o5_6Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire elapsed_time_ns_1_RNIV8ND11_0_27;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire elapsed_time_ns_1_RNIU7ND11_0_26;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire elapsed_time_ns_1_RNI0AND11_0_28;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire elapsed_time_ns_1_RNIP3OD11_0_30;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.N_432_i_g ;
    wire \delay_measurement_inst.delay_hc_timer.N_432_i ;
    wire il_min_comp2_D1;
    wire s3_phy_c;
    wire il_min_comp1_c;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire il_min_comp1_D1;
    wire il_max_comp1_c;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_10_13_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_10_14_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire bfn_10_15_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire il_max_comp1_D1;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire elapsed_time_ns_1_RNI62CED1_0_19;
    wire elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a5_1_1_9 ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.N_325_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2 ;
    wire elapsed_time_ns_1_RNIS4MD11_0_15;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_307_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0 ;
    wire \phase_controller_inst1.stoper_hc.N_45_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire il_max_comp2_D2;
    wire T12_c;
    wire state_ns_i_a3_1;
    wire delay_hc_input_c_g;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_stoper_state12_1_0_i ;
    wire bfn_11_13_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire bfn_11_14_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire bfn_11_15_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire elapsed_time_ns_1_RNID6DJ11_0_7;
    wire elapsed_time_ns_1_RNID6DJ11_0_7_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ;
    wire elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_i_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire elapsed_time_ns_1_RNIA3DJ11_0_4;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire elapsed_time_ns_1_RNIB4DJ11_0_5;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire elapsed_time_ns_1_RNIE7DJ11_0_8;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire elapsed_time_ns_1_RNIQ4OD11_0_31;
    wire elapsed_time_ns_1_RNIDP2KD1_0_1;
    wire \phase_controller_inst1.stoper_hc.target_time_7_f0_0_1Z0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.N_325 ;
    wire \phase_controller_inst1.stoper_hc.N_327 ;
    wire \phase_controller_inst1.stoper_hc.target_time_7_f0_0_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa_0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_433_i ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire elapsed_time_ns_1_RNI81DJ11_0_2;
    wire elapsed_time_ns_1_RNI81DJ11_0_2_cascade_;
    wire elapsed_time_ns_1_RNIQURR91_0_3;
    wire \phase_controller_inst1.stoper_hc.N_283 ;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_ ;
    wire \phase_controller_inst1.N_56 ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst2.start_timer_hc_RNOZ0Z_0_cascade_ ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.start_timer_tr_0_sqmuxa_cascade_ ;
    wire bfn_11_21_0_;
    wire \current_shift_inst.control_input_1_cry_0 ;
    wire \current_shift_inst.control_inputZ0Z_2 ;
    wire \current_shift_inst.control_input_1_cry_1 ;
    wire \current_shift_inst.control_inputZ0Z_3 ;
    wire \current_shift_inst.control_input_1_cry_2 ;
    wire \current_shift_inst.control_inputZ0Z_4 ;
    wire \current_shift_inst.control_input_1_cry_3 ;
    wire \current_shift_inst.control_input_1_cry_4 ;
    wire \current_shift_inst.control_input_1_cry_5 ;
    wire \current_shift_inst.control_inputZ0Z_7 ;
    wire \current_shift_inst.control_input_1_cry_6 ;
    wire \current_shift_inst.control_input_1_cry_7 ;
    wire bfn_11_22_0_;
    wire \current_shift_inst.control_input_1_cry_8 ;
    wire \current_shift_inst.control_inputZ0Z_10 ;
    wire \current_shift_inst.control_input_1_cry_9 ;
    wire \current_shift_inst.control_input_1_cry_10 ;
    wire \current_shift_inst.control_input_1_axb_10 ;
    wire \current_shift_inst.control_inputZ0Z_9 ;
    wire start_stop_c;
    wire phase_controller_inst1_state_4;
    wire il_min_comp2_D2;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire T23_c;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ;
    wire \current_shift_inst.PI_CTRL.N_74_16_cascade_ ;
    wire \current_shift_inst.control_inputZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_12_11_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire bfn_12_12_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.control_inputZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.control_inputZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_inputZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire \current_shift_inst.control_inputZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHEZ0 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_12_15_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_12_16_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_17 ;
    wire bfn_12_17_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire bfn_12_18_0_;
    wire \current_shift_inst.un38_control_input_cry_0_c_THRU_CO ;
    wire \current_shift_inst.un38_control_input_cry_0 ;
    wire \current_shift_inst.un38_control_input_cry_1 ;
    wire \current_shift_inst.un38_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2 ;
    wire \current_shift_inst.un38_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3 ;
    wire \current_shift_inst.un38_control_input_cry_4 ;
    wire \current_shift_inst.un38_control_input_cry_5 ;
    wire \current_shift_inst.un38_control_input_cry_6 ;
    wire \current_shift_inst.un38_control_input_cry_7_c_RNOZ0 ;
    wire bfn_12_19_0_;
    wire \current_shift_inst.un38_control_input_cry_7 ;
    wire \current_shift_inst.un38_control_input_cry_8 ;
    wire \current_shift_inst.un38_control_input_cry_9 ;
    wire \current_shift_inst.un38_control_input_cry_10 ;
    wire \current_shift_inst.un38_control_input_cry_11 ;
    wire \current_shift_inst.un38_control_input_cry_12 ;
    wire \current_shift_inst.un38_control_input_cry_13 ;
    wire \current_shift_inst.un38_control_input_cry_14 ;
    wire bfn_12_20_0_;
    wire \current_shift_inst.un38_control_input_cry_15 ;
    wire \current_shift_inst.un38_control_input_cry_16 ;
    wire \current_shift_inst.un38_control_input_cry_17 ;
    wire \current_shift_inst.un38_control_input_cry_18 ;
    wire \current_shift_inst.control_input_1_axb_0 ;
    wire \current_shift_inst.un38_control_input_cry_19 ;
    wire \current_shift_inst.control_input_1_axb_1 ;
    wire \current_shift_inst.un38_control_input_cry_20 ;
    wire \current_shift_inst.control_input_1_axb_2 ;
    wire \current_shift_inst.un38_control_input_cry_21 ;
    wire \current_shift_inst.un38_control_input_cry_22 ;
    wire \current_shift_inst.control_input_1_axb_3 ;
    wire bfn_12_21_0_;
    wire \current_shift_inst.control_input_1_axb_4 ;
    wire \current_shift_inst.un38_control_input_cry_23 ;
    wire \current_shift_inst.control_input_1_axb_5 ;
    wire \current_shift_inst.un38_control_input_cry_24 ;
    wire \current_shift_inst.control_input_1_axb_6 ;
    wire \current_shift_inst.un38_control_input_cry_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.control_input_1_axb_7 ;
    wire \current_shift_inst.un38_control_input_cry_26 ;
    wire \current_shift_inst.control_input_1_axb_8 ;
    wire \current_shift_inst.un38_control_input_cry_27 ;
    wire \current_shift_inst.control_input_1_axb_9 ;
    wire \current_shift_inst.un38_control_input_cry_28 ;
    wire \current_shift_inst.un38_control_input_cry_29 ;
    wire \current_shift_inst.un38_control_input_cry_29_THRU_CO ;
    wire \current_shift_inst.un38_control_input_axb_30 ;
    wire \phase_controller_inst2.time_passed_RNI9M3O ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire T01_c;
    wire s1_phy_c;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire T45_c;
    wire \current_shift_inst.timer_s1.N_166_i ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \pll_inst.red_c_i ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_62 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.N_74_21 ;
    wire \current_shift_inst.PI_CTRL.N_72 ;
    wire \current_shift_inst.PI_CTRL.N_75 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ;
    wire bfn_13_11_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ;
    wire bfn_13_12_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ;
    wire bfn_13_13_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ;
    wire bfn_13_14_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_31 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.N_45 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.un38_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_1_c_RNOZ0 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire il_max_comp1_D2;
    wire state_3;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire il_min_comp1_D2;
    wire bfn_13_19_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire bfn_13_20_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire bfn_13_21_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire bfn_13_22_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire bfn_13_24_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_13_25_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_13_26_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_13_27_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_167_i ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ;
    wire \delay_measurement_inst.delay_tr_timer.N_358_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ;
    wire elapsed_time_ns_1_RNIFJ2591_0_7_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_382_i ;
    wire elapsed_time_ns_1_RNIIU2KD1_0_6;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6 ;
    wire \phase_controller_inst1.stoper_tr.N_235_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa_0 ;
    wire \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst2.stoper_hc.un1_stoper_state12_1_0_i ;
    wire \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.N_45 ;
    wire \phase_controller_inst1.stoper_tr.N_219 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.un38_control_input_cry_0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_12 ;
    wire bfn_15_7_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integrator_i_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_2 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire bfn_15_8_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire bfn_15_9_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_23 ;
    wire bfn_15_10_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_25 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_28 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_0_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_30 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_30 ;
    wire bfn_15_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6 ;
    wire \delay_measurement_inst.delay_tr_timer.N_363_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ;
    wire elapsed_time_ns_1_RNI3JIF91_0_29;
    wire elapsed_time_ns_1_RNIRBJF91_0_30;
    wire elapsed_time_ns_1_RNIRAIF91_0_21;
    wire elapsed_time_ns_1_RNI3JIF91_0_29_cascade_;
    wire elapsed_time_ns_1_RNIQ9IF91_0_20;
    wire elapsed_time_ns_1_RNISBIF91_0_22;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_o5_7Z0Z_15_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_381 ;
    wire \delay_measurement_inst.delay_tr_timer.N_359_1 ;
    wire \delay_measurement_inst.delay_tr_timer.N_381_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ;
    wire elapsed_time_ns_1_RNISAHF91_0_13_cascade_;
    wire elapsed_time_ns_1_RNIUCHF91_0_15_cascade_;
    wire \phase_controller_inst1.stoper_tr.N_251_cascade_ ;
    wire elapsed_time_ns_1_RNIDH2591_0_5_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3Z0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.N_241_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_ ;
    wire elapsed_time_ns_1_RNIPFL2M1_0_1;
    wire elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_7_f0_0_1Z0Z_1 ;
    wire elapsed_time_ns_1_RNISCJF91_0_31_cascade_;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire bfn_15_17_0_;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire bfn_15_18_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire bfn_15_19_0_;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_15_20_0_;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire delay_tr_input_c_g;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.N_74_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0 ;
    wire \current_shift_inst.PI_CTRL.N_103 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_380 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ;
    wire \delay_measurement_inst.delay_tr_timer.N_341 ;
    wire \delay_measurement_inst.delay_tr_timer.N_367 ;
    wire \delay_measurement_inst.delay_tr_timer.N_367_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_378 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.N_349 ;
    wire elapsed_time_ns_1_RNIVEIF91_0_25;
    wire elapsed_time_ns_1_RNIVEIF91_0_25_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_o5_6Z0Z_15 ;
    wire elapsed_time_ns_1_RNI2IIF91_0_28;
    wire \delay_measurement_inst.delay_tr_timer.N_345 ;
    wire \delay_measurement_inst.delay_tr_timer.N_348 ;
    wire \delay_measurement_inst.delay_tr_timer.N_347 ;
    wire \delay_measurement_inst.delay_tr_timer.N_347_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_365 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ;
    wire elapsed_time_ns_1_RNI0GIF91_0_26;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6 ;
    wire elapsed_time_ns_1_RNITCIF91_0_23;
    wire elapsed_time_ns_1_RNITCIF91_0_23_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_0_15 ;
    wire elapsed_time_ns_1_RNI1HIF91_0_27;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ;
    wire elapsed_time_ns_1_RNIUDIF91_0_24;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_434_i ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.N_55 ;
    wire \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ;
    wire elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_;
    wire elapsed_time_ns_1_RNI1OL2M1_0_9;
    wire \phase_controller_inst1.stoper_tr.N_244 ;
    wire \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_0_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_249_cascade_ ;
    wire elapsed_time_ns_1_RNIFJ2591_0_7;
    wire elapsed_time_ns_1_RNIGK2591_0_8;
    wire elapsed_time_ns_1_RNIUKL2M1_0_6;
    wire \phase_controller_inst1.stoper_tr.N_250 ;
    wire \phase_controller_inst1.stoper_tr.target_time_7_f0_i_1Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9 ;
    wire elapsed_time_ns_1_RNIAE2591_0_2;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_0_2 ;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2 ;
    wire elapsed_time_ns_1_RNIRHL2M1_0_3;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2_cascade_ ;
    wire elapsed_time_ns_1_RNIUCHF91_0_15;
    wire \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9 ;
    wire elapsed_time_ns_1_RNIDH2591_0_5;
    wire \phase_controller_inst1.stoper_tr.N_249 ;
    wire elapsed_time_ns_1_RNICG2591_0_4;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un38_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.N_166_i_g ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.control_inputZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_c_RNOZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire bfn_17_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire bfn_17_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire bfn_17_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_17_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.delay_tr_timer.N_434_i_g ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire bfn_17_14_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_17_15_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_17_16_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.un1_stoper_state12_1_0_i ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire bfn_17_17_0_;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_17_18_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire bfn_17_19_0_;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire bfn_17_20_0_;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.N_1310_i ;
    wire \phase_controller_inst2.stoper_tr.N_45_cascade_ ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_18_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_18_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_18_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_18_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_435_i ;
    wire elapsed_time_ns_1_RNIR9HF91_0_12;
    wire elapsed_time_ns_1_RNIDE4DM1_0_14;
    wire elapsed_time_ns_1_RNIP7HF91_0_10;
    wire elapsed_time_ns_1_RNIQ8HF91_0_11;
    wire elapsed_time_ns_1_RNIFG4DM1_0_16;
    wire \phase_controller_inst1.stoper_tr.N_241 ;
    wire elapsed_time_ns_1_RNISAHF91_0_13;
    wire elapsed_time_ns_1_RNIIJ4DM1_0_19;
    wire elapsed_time_ns_1_RNIHI4DM1_0_18;
    wire elapsed_time_ns_1_RNIGH4DM1_0_17;
    wire elapsed_time_ns_1_RNISCJF91_0_31;
    wire \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa_0 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_18_13_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_18_14_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_18_15_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_18_16_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_18_17_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_17 ;
    wire bfn_18_18_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire red_c_g;
    wire \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire bfn_18_19_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84ADZ0 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_18_20_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_18_21_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire \phase_controller_inst2.stoper_tr.un1_stoper_state12_1_0_i ;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__20453),
            .RESETB(N__28073),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__40612),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__40608),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__19364,N__19357,N__19362,N__19356,N__19363,N__19355,N__19365,N__19352,N__19358,N__19351,N__19359,N__19353,N__19360,N__19354,N__19361}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__40615,N__40611,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__40609,N__40614,N__40610,N__40613}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__40469),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__40462),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .ADDSUBBOT(),
            .A({dangling_wire_74,N__19411,N__19416,N__19412,N__19417,N__19413,N__19782,N__19692,N__19737,N__19767,N__18231,N__19540,N__18813,N__19102,N__19117,N__19132}),
            .C({dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90}),
            .B({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,N__40468,N__40465,dangling_wire_98,dangling_wire_99,dangling_wire_100,N__40463,N__40467,N__40464,N__40466}),
            .OHOLDTOP(),
            .O({dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__45222),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__45224),
            .DIN(N__45223),
            .DOUT(N__45222),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__45224),
            .PADOUT(N__45223),
            .PADIN(N__45222),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T01_obuf_iopad (
            .OE(N__45213),
            .DIN(N__45212),
            .DOUT(N__45211),
            .PACKAGEPIN(T01));
    defparam T01_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T01_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T01_obuf_preio (
            .PADOEN(N__45213),
            .PADOUT(N__45212),
            .PADIN(N__45211),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27986),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__45204),
            .DIN(N__45203),
            .DOUT(N__45202),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__45204),
            .PADOUT(N__45203),
            .PADIN(N__45202),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__45195),
            .DIN(N__45194),
            .DOUT(N__45193),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__45195),
            .PADOUT(N__45194),
            .PADIN(N__45193),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__45186),
            .DIN(N__45185),
            .DOUT(N__45184),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__45186),
            .PADOUT(N__45185),
            .PADIN(N__45184),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26549),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__45177),
            .DIN(N__45176),
            .DOUT(N__45175),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__45177),
            .PADOUT(N__45176),
            .PADIN(N__45175),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20345),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__45168),
            .DIN(N__45167),
            .DOUT(N__45166),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__45168),
            .PADOUT(N__45167),
            .PADIN(N__45166),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__45159),
            .DIN(N__45158),
            .DOUT(N__45157),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__45159),
            .PADOUT(N__45158),
            .PADIN(N__45157),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29384),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__45150),
            .DIN(N__45149),
            .DOUT(N__45148),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__45150),
            .PADOUT(N__45149),
            .PADIN(N__45148),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25076),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__45141),
            .DIN(N__45140),
            .DOUT(N__45139),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__45141),
            .PADOUT(N__45140),
            .PADIN(N__45139),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__45132),
            .DIN(N__45131),
            .DOUT(N__45130),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__45132),
            .PADOUT(N__45131),
            .PADIN(N__45130),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27962),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__45123),
            .DIN(N__45122),
            .DOUT(N__45121),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__45123),
            .PADOUT(N__45122),
            .PADIN(N__45121),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23114),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__45114),
            .DIN(N__45113),
            .DOUT(N__45112),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__45114),
            .PADOUT(N__45113),
            .PADIN(N__45112),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__45105),
            .DIN(N__45104),
            .DOUT(N__45103),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__45105),
            .PADOUT(N__45104),
            .PADIN(N__45103),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23906),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T45_obuf_iopad (
            .OE(N__45096),
            .DIN(N__45095),
            .DOUT(N__45094),
            .PACKAGEPIN(T45));
    defparam T45_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T45_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T45_obuf_preio (
            .PADOEN(N__45096),
            .PADOUT(N__45095),
            .PADIN(N__45094),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27854),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__45087),
            .DIN(N__45086),
            .DOUT(N__45085),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__45087),
            .PADOUT(N__45086),
            .PADIN(N__45085),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__45078),
            .DIN(N__45077),
            .DOUT(N__45076),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__45078),
            .PADOUT(N__45077),
            .PADIN(N__45076),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__10663 (
            .O(N__45059),
            .I(N__45055));
    InMux I__10662 (
            .O(N__45058),
            .I(N__45052));
    LocalMux I__10661 (
            .O(N__45055),
            .I(N__45049));
    LocalMux I__10660 (
            .O(N__45052),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__10659 (
            .O(N__45049),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__10658 (
            .O(N__45044),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__10657 (
            .O(N__45041),
            .I(N__45037));
    InMux I__10656 (
            .O(N__45040),
            .I(N__45034));
    LocalMux I__10655 (
            .O(N__45037),
            .I(N__45031));
    LocalMux I__10654 (
            .O(N__45034),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv12 I__10653 (
            .O(N__45031),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__10652 (
            .O(N__45026),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__10651 (
            .O(N__45023),
            .I(N__45019));
    InMux I__10650 (
            .O(N__45022),
            .I(N__45016));
    LocalMux I__10649 (
            .O(N__45019),
            .I(N__45013));
    LocalMux I__10648 (
            .O(N__45016),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv12 I__10647 (
            .O(N__45013),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__10646 (
            .O(N__45008),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__10645 (
            .O(N__45005),
            .I(N__45001));
    InMux I__10644 (
            .O(N__45004),
            .I(N__44998));
    LocalMux I__10643 (
            .O(N__45001),
            .I(N__44995));
    LocalMux I__10642 (
            .O(N__44998),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__10641 (
            .O(N__44995),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__10640 (
            .O(N__44990),
            .I(bfn_18_21_0_));
    InMux I__10639 (
            .O(N__44987),
            .I(N__44983));
    InMux I__10638 (
            .O(N__44986),
            .I(N__44980));
    LocalMux I__10637 (
            .O(N__44983),
            .I(N__44977));
    LocalMux I__10636 (
            .O(N__44980),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__10635 (
            .O(N__44977),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__10634 (
            .O(N__44972),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__10633 (
            .O(N__44969),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__10632 (
            .O(N__44966),
            .I(N__44962));
    InMux I__10631 (
            .O(N__44965),
            .I(N__44959));
    LocalMux I__10630 (
            .O(N__44962),
            .I(N__44956));
    LocalMux I__10629 (
            .O(N__44959),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__10628 (
            .O(N__44956),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    ClkMux I__10627 (
            .O(N__44951),
            .I(N__44591));
    ClkMux I__10626 (
            .O(N__44950),
            .I(N__44591));
    ClkMux I__10625 (
            .O(N__44949),
            .I(N__44591));
    ClkMux I__10624 (
            .O(N__44948),
            .I(N__44591));
    ClkMux I__10623 (
            .O(N__44947),
            .I(N__44591));
    ClkMux I__10622 (
            .O(N__44946),
            .I(N__44591));
    ClkMux I__10621 (
            .O(N__44945),
            .I(N__44591));
    ClkMux I__10620 (
            .O(N__44944),
            .I(N__44591));
    ClkMux I__10619 (
            .O(N__44943),
            .I(N__44591));
    ClkMux I__10618 (
            .O(N__44942),
            .I(N__44591));
    ClkMux I__10617 (
            .O(N__44941),
            .I(N__44591));
    ClkMux I__10616 (
            .O(N__44940),
            .I(N__44591));
    ClkMux I__10615 (
            .O(N__44939),
            .I(N__44591));
    ClkMux I__10614 (
            .O(N__44938),
            .I(N__44591));
    ClkMux I__10613 (
            .O(N__44937),
            .I(N__44591));
    ClkMux I__10612 (
            .O(N__44936),
            .I(N__44591));
    ClkMux I__10611 (
            .O(N__44935),
            .I(N__44591));
    ClkMux I__10610 (
            .O(N__44934),
            .I(N__44591));
    ClkMux I__10609 (
            .O(N__44933),
            .I(N__44591));
    ClkMux I__10608 (
            .O(N__44932),
            .I(N__44591));
    ClkMux I__10607 (
            .O(N__44931),
            .I(N__44591));
    ClkMux I__10606 (
            .O(N__44930),
            .I(N__44591));
    ClkMux I__10605 (
            .O(N__44929),
            .I(N__44591));
    ClkMux I__10604 (
            .O(N__44928),
            .I(N__44591));
    ClkMux I__10603 (
            .O(N__44927),
            .I(N__44591));
    ClkMux I__10602 (
            .O(N__44926),
            .I(N__44591));
    ClkMux I__10601 (
            .O(N__44925),
            .I(N__44591));
    ClkMux I__10600 (
            .O(N__44924),
            .I(N__44591));
    ClkMux I__10599 (
            .O(N__44923),
            .I(N__44591));
    ClkMux I__10598 (
            .O(N__44922),
            .I(N__44591));
    ClkMux I__10597 (
            .O(N__44921),
            .I(N__44591));
    ClkMux I__10596 (
            .O(N__44920),
            .I(N__44591));
    ClkMux I__10595 (
            .O(N__44919),
            .I(N__44591));
    ClkMux I__10594 (
            .O(N__44918),
            .I(N__44591));
    ClkMux I__10593 (
            .O(N__44917),
            .I(N__44591));
    ClkMux I__10592 (
            .O(N__44916),
            .I(N__44591));
    ClkMux I__10591 (
            .O(N__44915),
            .I(N__44591));
    ClkMux I__10590 (
            .O(N__44914),
            .I(N__44591));
    ClkMux I__10589 (
            .O(N__44913),
            .I(N__44591));
    ClkMux I__10588 (
            .O(N__44912),
            .I(N__44591));
    ClkMux I__10587 (
            .O(N__44911),
            .I(N__44591));
    ClkMux I__10586 (
            .O(N__44910),
            .I(N__44591));
    ClkMux I__10585 (
            .O(N__44909),
            .I(N__44591));
    ClkMux I__10584 (
            .O(N__44908),
            .I(N__44591));
    ClkMux I__10583 (
            .O(N__44907),
            .I(N__44591));
    ClkMux I__10582 (
            .O(N__44906),
            .I(N__44591));
    ClkMux I__10581 (
            .O(N__44905),
            .I(N__44591));
    ClkMux I__10580 (
            .O(N__44904),
            .I(N__44591));
    ClkMux I__10579 (
            .O(N__44903),
            .I(N__44591));
    ClkMux I__10578 (
            .O(N__44902),
            .I(N__44591));
    ClkMux I__10577 (
            .O(N__44901),
            .I(N__44591));
    ClkMux I__10576 (
            .O(N__44900),
            .I(N__44591));
    ClkMux I__10575 (
            .O(N__44899),
            .I(N__44591));
    ClkMux I__10574 (
            .O(N__44898),
            .I(N__44591));
    ClkMux I__10573 (
            .O(N__44897),
            .I(N__44591));
    ClkMux I__10572 (
            .O(N__44896),
            .I(N__44591));
    ClkMux I__10571 (
            .O(N__44895),
            .I(N__44591));
    ClkMux I__10570 (
            .O(N__44894),
            .I(N__44591));
    ClkMux I__10569 (
            .O(N__44893),
            .I(N__44591));
    ClkMux I__10568 (
            .O(N__44892),
            .I(N__44591));
    ClkMux I__10567 (
            .O(N__44891),
            .I(N__44591));
    ClkMux I__10566 (
            .O(N__44890),
            .I(N__44591));
    ClkMux I__10565 (
            .O(N__44889),
            .I(N__44591));
    ClkMux I__10564 (
            .O(N__44888),
            .I(N__44591));
    ClkMux I__10563 (
            .O(N__44887),
            .I(N__44591));
    ClkMux I__10562 (
            .O(N__44886),
            .I(N__44591));
    ClkMux I__10561 (
            .O(N__44885),
            .I(N__44591));
    ClkMux I__10560 (
            .O(N__44884),
            .I(N__44591));
    ClkMux I__10559 (
            .O(N__44883),
            .I(N__44591));
    ClkMux I__10558 (
            .O(N__44882),
            .I(N__44591));
    ClkMux I__10557 (
            .O(N__44881),
            .I(N__44591));
    ClkMux I__10556 (
            .O(N__44880),
            .I(N__44591));
    ClkMux I__10555 (
            .O(N__44879),
            .I(N__44591));
    ClkMux I__10554 (
            .O(N__44878),
            .I(N__44591));
    ClkMux I__10553 (
            .O(N__44877),
            .I(N__44591));
    ClkMux I__10552 (
            .O(N__44876),
            .I(N__44591));
    ClkMux I__10551 (
            .O(N__44875),
            .I(N__44591));
    ClkMux I__10550 (
            .O(N__44874),
            .I(N__44591));
    ClkMux I__10549 (
            .O(N__44873),
            .I(N__44591));
    ClkMux I__10548 (
            .O(N__44872),
            .I(N__44591));
    ClkMux I__10547 (
            .O(N__44871),
            .I(N__44591));
    ClkMux I__10546 (
            .O(N__44870),
            .I(N__44591));
    ClkMux I__10545 (
            .O(N__44869),
            .I(N__44591));
    ClkMux I__10544 (
            .O(N__44868),
            .I(N__44591));
    ClkMux I__10543 (
            .O(N__44867),
            .I(N__44591));
    ClkMux I__10542 (
            .O(N__44866),
            .I(N__44591));
    ClkMux I__10541 (
            .O(N__44865),
            .I(N__44591));
    ClkMux I__10540 (
            .O(N__44864),
            .I(N__44591));
    ClkMux I__10539 (
            .O(N__44863),
            .I(N__44591));
    ClkMux I__10538 (
            .O(N__44862),
            .I(N__44591));
    ClkMux I__10537 (
            .O(N__44861),
            .I(N__44591));
    ClkMux I__10536 (
            .O(N__44860),
            .I(N__44591));
    ClkMux I__10535 (
            .O(N__44859),
            .I(N__44591));
    ClkMux I__10534 (
            .O(N__44858),
            .I(N__44591));
    ClkMux I__10533 (
            .O(N__44857),
            .I(N__44591));
    ClkMux I__10532 (
            .O(N__44856),
            .I(N__44591));
    ClkMux I__10531 (
            .O(N__44855),
            .I(N__44591));
    ClkMux I__10530 (
            .O(N__44854),
            .I(N__44591));
    ClkMux I__10529 (
            .O(N__44853),
            .I(N__44591));
    ClkMux I__10528 (
            .O(N__44852),
            .I(N__44591));
    ClkMux I__10527 (
            .O(N__44851),
            .I(N__44591));
    ClkMux I__10526 (
            .O(N__44850),
            .I(N__44591));
    ClkMux I__10525 (
            .O(N__44849),
            .I(N__44591));
    ClkMux I__10524 (
            .O(N__44848),
            .I(N__44591));
    ClkMux I__10523 (
            .O(N__44847),
            .I(N__44591));
    ClkMux I__10522 (
            .O(N__44846),
            .I(N__44591));
    ClkMux I__10521 (
            .O(N__44845),
            .I(N__44591));
    ClkMux I__10520 (
            .O(N__44844),
            .I(N__44591));
    ClkMux I__10519 (
            .O(N__44843),
            .I(N__44591));
    ClkMux I__10518 (
            .O(N__44842),
            .I(N__44591));
    ClkMux I__10517 (
            .O(N__44841),
            .I(N__44591));
    ClkMux I__10516 (
            .O(N__44840),
            .I(N__44591));
    ClkMux I__10515 (
            .O(N__44839),
            .I(N__44591));
    ClkMux I__10514 (
            .O(N__44838),
            .I(N__44591));
    ClkMux I__10513 (
            .O(N__44837),
            .I(N__44591));
    ClkMux I__10512 (
            .O(N__44836),
            .I(N__44591));
    ClkMux I__10511 (
            .O(N__44835),
            .I(N__44591));
    ClkMux I__10510 (
            .O(N__44834),
            .I(N__44591));
    ClkMux I__10509 (
            .O(N__44833),
            .I(N__44591));
    ClkMux I__10508 (
            .O(N__44832),
            .I(N__44591));
    GlobalMux I__10507 (
            .O(N__44591),
            .I(clk_100mhz_0));
    SRMux I__10506 (
            .O(N__44588),
            .I(N__44584));
    SRMux I__10505 (
            .O(N__44587),
            .I(N__44581));
    LocalMux I__10504 (
            .O(N__44584),
            .I(N__44578));
    LocalMux I__10503 (
            .O(N__44581),
            .I(N__44573));
    Span4Mux_v I__10502 (
            .O(N__44578),
            .I(N__44570));
    SRMux I__10501 (
            .O(N__44577),
            .I(N__44567));
    SRMux I__10500 (
            .O(N__44576),
            .I(N__44564));
    Span4Mux_h I__10499 (
            .O(N__44573),
            .I(N__44561));
    Span4Mux_h I__10498 (
            .O(N__44570),
            .I(N__44556));
    LocalMux I__10497 (
            .O(N__44567),
            .I(N__44556));
    LocalMux I__10496 (
            .O(N__44564),
            .I(N__44553));
    Odrv4 I__10495 (
            .O(N__44561),
            .I(\phase_controller_inst2.stoper_tr.un1_stoper_state12_1_0_i ));
    Odrv4 I__10494 (
            .O(N__44556),
            .I(\phase_controller_inst2.stoper_tr.un1_stoper_state12_1_0_i ));
    Odrv4 I__10493 (
            .O(N__44553),
            .I(\phase_controller_inst2.stoper_tr.un1_stoper_state12_1_0_i ));
    InMux I__10492 (
            .O(N__44546),
            .I(N__44542));
    InMux I__10491 (
            .O(N__44545),
            .I(N__44539));
    LocalMux I__10490 (
            .O(N__44542),
            .I(N__44536));
    LocalMux I__10489 (
            .O(N__44539),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__10488 (
            .O(N__44536),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__10487 (
            .O(N__44531),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__10486 (
            .O(N__44528),
            .I(N__44524));
    InMux I__10485 (
            .O(N__44527),
            .I(N__44521));
    LocalMux I__10484 (
            .O(N__44524),
            .I(N__44518));
    LocalMux I__10483 (
            .O(N__44521),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__10482 (
            .O(N__44518),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__10481 (
            .O(N__44513),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__10480 (
            .O(N__44510),
            .I(N__44506));
    InMux I__10479 (
            .O(N__44509),
            .I(N__44503));
    LocalMux I__10478 (
            .O(N__44506),
            .I(N__44500));
    LocalMux I__10477 (
            .O(N__44503),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv12 I__10476 (
            .O(N__44500),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__10475 (
            .O(N__44495),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__10474 (
            .O(N__44492),
            .I(N__44488));
    InMux I__10473 (
            .O(N__44491),
            .I(N__44485));
    LocalMux I__10472 (
            .O(N__44488),
            .I(N__44482));
    LocalMux I__10471 (
            .O(N__44485),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv12 I__10470 (
            .O(N__44482),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__10469 (
            .O(N__44477),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__10468 (
            .O(N__44474),
            .I(N__44470));
    InMux I__10467 (
            .O(N__44473),
            .I(N__44467));
    LocalMux I__10466 (
            .O(N__44470),
            .I(N__44464));
    LocalMux I__10465 (
            .O(N__44467),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__10464 (
            .O(N__44464),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__10463 (
            .O(N__44459),
            .I(bfn_18_20_0_));
    InMux I__10462 (
            .O(N__44456),
            .I(N__44452));
    InMux I__10461 (
            .O(N__44455),
            .I(N__44449));
    LocalMux I__10460 (
            .O(N__44452),
            .I(N__44446));
    LocalMux I__10459 (
            .O(N__44449),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__10458 (
            .O(N__44446),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__10457 (
            .O(N__44441),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__10456 (
            .O(N__44438),
            .I(N__44434));
    InMux I__10455 (
            .O(N__44437),
            .I(N__44431));
    LocalMux I__10454 (
            .O(N__44434),
            .I(N__44428));
    LocalMux I__10453 (
            .O(N__44431),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__10452 (
            .O(N__44428),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__10451 (
            .O(N__44423),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__10450 (
            .O(N__44420),
            .I(N__44416));
    InMux I__10449 (
            .O(N__44419),
            .I(N__44413));
    LocalMux I__10448 (
            .O(N__44416),
            .I(N__44410));
    LocalMux I__10447 (
            .O(N__44413),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__10446 (
            .O(N__44410),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__10445 (
            .O(N__44405),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__10444 (
            .O(N__44402),
            .I(N__44398));
    InMux I__10443 (
            .O(N__44401),
            .I(N__44395));
    LocalMux I__10442 (
            .O(N__44398),
            .I(N__44392));
    LocalMux I__10441 (
            .O(N__44395),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__10440 (
            .O(N__44392),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__10439 (
            .O(N__44387),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__10438 (
            .O(N__44384),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__10437 (
            .O(N__44381),
            .I(N__44371));
    InMux I__10436 (
            .O(N__44380),
            .I(N__44371));
    InMux I__10435 (
            .O(N__44379),
            .I(N__44371));
    InMux I__10434 (
            .O(N__44378),
            .I(N__44368));
    LocalMux I__10433 (
            .O(N__44371),
            .I(N__44364));
    LocalMux I__10432 (
            .O(N__44368),
            .I(N__44361));
    CascadeMux I__10431 (
            .O(N__44367),
            .I(N__44358));
    Span4Mux_h I__10430 (
            .O(N__44364),
            .I(N__44354));
    Span4Mux_v I__10429 (
            .O(N__44361),
            .I(N__44351));
    InMux I__10428 (
            .O(N__44358),
            .I(N__44346));
    InMux I__10427 (
            .O(N__44357),
            .I(N__44346));
    Odrv4 I__10426 (
            .O(N__44354),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__10425 (
            .O(N__44351),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__10424 (
            .O(N__44346),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__10423 (
            .O(N__44339),
            .I(N__44328));
    CascadeMux I__10422 (
            .O(N__44338),
            .I(N__44323));
    InMux I__10421 (
            .O(N__44337),
            .I(N__44308));
    InMux I__10420 (
            .O(N__44336),
            .I(N__44305));
    InMux I__10419 (
            .O(N__44335),
            .I(N__44302));
    InMux I__10418 (
            .O(N__44334),
            .I(N__44299));
    InMux I__10417 (
            .O(N__44333),
            .I(N__44296));
    InMux I__10416 (
            .O(N__44332),
            .I(N__44293));
    InMux I__10415 (
            .O(N__44331),
            .I(N__44290));
    InMux I__10414 (
            .O(N__44328),
            .I(N__44285));
    InMux I__10413 (
            .O(N__44327),
            .I(N__44285));
    InMux I__10412 (
            .O(N__44326),
            .I(N__44282));
    InMux I__10411 (
            .O(N__44323),
            .I(N__44275));
    InMux I__10410 (
            .O(N__44322),
            .I(N__44275));
    InMux I__10409 (
            .O(N__44321),
            .I(N__44275));
    InMux I__10408 (
            .O(N__44320),
            .I(N__44272));
    InMux I__10407 (
            .O(N__44319),
            .I(N__44267));
    InMux I__10406 (
            .O(N__44318),
            .I(N__44267));
    InMux I__10405 (
            .O(N__44317),
            .I(N__44262));
    InMux I__10404 (
            .O(N__44316),
            .I(N__44262));
    InMux I__10403 (
            .O(N__44315),
            .I(N__44259));
    InMux I__10402 (
            .O(N__44314),
            .I(N__44254));
    InMux I__10401 (
            .O(N__44313),
            .I(N__44254));
    InMux I__10400 (
            .O(N__44312),
            .I(N__44249));
    InMux I__10399 (
            .O(N__44311),
            .I(N__44249));
    LocalMux I__10398 (
            .O(N__44308),
            .I(N__44246));
    LocalMux I__10397 (
            .O(N__44305),
            .I(N__44243));
    LocalMux I__10396 (
            .O(N__44302),
            .I(N__44240));
    LocalMux I__10395 (
            .O(N__44299),
            .I(N__44235));
    LocalMux I__10394 (
            .O(N__44296),
            .I(N__44211));
    LocalMux I__10393 (
            .O(N__44293),
            .I(N__44205));
    LocalMux I__10392 (
            .O(N__44290),
            .I(N__44202));
    LocalMux I__10391 (
            .O(N__44285),
            .I(N__44196));
    LocalMux I__10390 (
            .O(N__44282),
            .I(N__44193));
    LocalMux I__10389 (
            .O(N__44275),
            .I(N__44190));
    LocalMux I__10388 (
            .O(N__44272),
            .I(N__44165));
    LocalMux I__10387 (
            .O(N__44267),
            .I(N__44154));
    LocalMux I__10386 (
            .O(N__44262),
            .I(N__44147));
    LocalMux I__10385 (
            .O(N__44259),
            .I(N__44140));
    LocalMux I__10384 (
            .O(N__44254),
            .I(N__44132));
    LocalMux I__10383 (
            .O(N__44249),
            .I(N__44126));
    Glb2LocalMux I__10382 (
            .O(N__44246),
            .I(N__43874));
    Glb2LocalMux I__10381 (
            .O(N__44243),
            .I(N__43874));
    Glb2LocalMux I__10380 (
            .O(N__44240),
            .I(N__43874));
    SRMux I__10379 (
            .O(N__44239),
            .I(N__43874));
    SRMux I__10378 (
            .O(N__44238),
            .I(N__43874));
    Glb2LocalMux I__10377 (
            .O(N__44235),
            .I(N__43874));
    SRMux I__10376 (
            .O(N__44234),
            .I(N__43874));
    SRMux I__10375 (
            .O(N__44233),
            .I(N__43874));
    SRMux I__10374 (
            .O(N__44232),
            .I(N__43874));
    SRMux I__10373 (
            .O(N__44231),
            .I(N__43874));
    SRMux I__10372 (
            .O(N__44230),
            .I(N__43874));
    SRMux I__10371 (
            .O(N__44229),
            .I(N__43874));
    SRMux I__10370 (
            .O(N__44228),
            .I(N__43874));
    SRMux I__10369 (
            .O(N__44227),
            .I(N__43874));
    SRMux I__10368 (
            .O(N__44226),
            .I(N__43874));
    SRMux I__10367 (
            .O(N__44225),
            .I(N__43874));
    SRMux I__10366 (
            .O(N__44224),
            .I(N__43874));
    SRMux I__10365 (
            .O(N__44223),
            .I(N__43874));
    SRMux I__10364 (
            .O(N__44222),
            .I(N__43874));
    SRMux I__10363 (
            .O(N__44221),
            .I(N__43874));
    SRMux I__10362 (
            .O(N__44220),
            .I(N__43874));
    SRMux I__10361 (
            .O(N__44219),
            .I(N__43874));
    SRMux I__10360 (
            .O(N__44218),
            .I(N__43874));
    SRMux I__10359 (
            .O(N__44217),
            .I(N__43874));
    SRMux I__10358 (
            .O(N__44216),
            .I(N__43874));
    SRMux I__10357 (
            .O(N__44215),
            .I(N__43874));
    SRMux I__10356 (
            .O(N__44214),
            .I(N__43874));
    Glb2LocalMux I__10355 (
            .O(N__44211),
            .I(N__43874));
    SRMux I__10354 (
            .O(N__44210),
            .I(N__43874));
    SRMux I__10353 (
            .O(N__44209),
            .I(N__43874));
    SRMux I__10352 (
            .O(N__44208),
            .I(N__43874));
    Glb2LocalMux I__10351 (
            .O(N__44205),
            .I(N__43874));
    Glb2LocalMux I__10350 (
            .O(N__44202),
            .I(N__43874));
    SRMux I__10349 (
            .O(N__44201),
            .I(N__43874));
    SRMux I__10348 (
            .O(N__44200),
            .I(N__43874));
    SRMux I__10347 (
            .O(N__44199),
            .I(N__43874));
    Glb2LocalMux I__10346 (
            .O(N__44196),
            .I(N__43874));
    Glb2LocalMux I__10345 (
            .O(N__44193),
            .I(N__43874));
    Glb2LocalMux I__10344 (
            .O(N__44190),
            .I(N__43874));
    SRMux I__10343 (
            .O(N__44189),
            .I(N__43874));
    SRMux I__10342 (
            .O(N__44188),
            .I(N__43874));
    SRMux I__10341 (
            .O(N__44187),
            .I(N__43874));
    SRMux I__10340 (
            .O(N__44186),
            .I(N__43874));
    SRMux I__10339 (
            .O(N__44185),
            .I(N__43874));
    SRMux I__10338 (
            .O(N__44184),
            .I(N__43874));
    SRMux I__10337 (
            .O(N__44183),
            .I(N__43874));
    SRMux I__10336 (
            .O(N__44182),
            .I(N__43874));
    SRMux I__10335 (
            .O(N__44181),
            .I(N__43874));
    SRMux I__10334 (
            .O(N__44180),
            .I(N__43874));
    SRMux I__10333 (
            .O(N__44179),
            .I(N__43874));
    SRMux I__10332 (
            .O(N__44178),
            .I(N__43874));
    SRMux I__10331 (
            .O(N__44177),
            .I(N__43874));
    SRMux I__10330 (
            .O(N__44176),
            .I(N__43874));
    SRMux I__10329 (
            .O(N__44175),
            .I(N__43874));
    SRMux I__10328 (
            .O(N__44174),
            .I(N__43874));
    SRMux I__10327 (
            .O(N__44173),
            .I(N__43874));
    SRMux I__10326 (
            .O(N__44172),
            .I(N__43874));
    SRMux I__10325 (
            .O(N__44171),
            .I(N__43874));
    SRMux I__10324 (
            .O(N__44170),
            .I(N__43874));
    SRMux I__10323 (
            .O(N__44169),
            .I(N__43874));
    SRMux I__10322 (
            .O(N__44168),
            .I(N__43874));
    Glb2LocalMux I__10321 (
            .O(N__44165),
            .I(N__43874));
    SRMux I__10320 (
            .O(N__44164),
            .I(N__43874));
    SRMux I__10319 (
            .O(N__44163),
            .I(N__43874));
    SRMux I__10318 (
            .O(N__44162),
            .I(N__43874));
    SRMux I__10317 (
            .O(N__44161),
            .I(N__43874));
    SRMux I__10316 (
            .O(N__44160),
            .I(N__43874));
    SRMux I__10315 (
            .O(N__44159),
            .I(N__43874));
    SRMux I__10314 (
            .O(N__44158),
            .I(N__43874));
    SRMux I__10313 (
            .O(N__44157),
            .I(N__43874));
    Glb2LocalMux I__10312 (
            .O(N__44154),
            .I(N__43874));
    SRMux I__10311 (
            .O(N__44153),
            .I(N__43874));
    SRMux I__10310 (
            .O(N__44152),
            .I(N__43874));
    SRMux I__10309 (
            .O(N__44151),
            .I(N__43874));
    SRMux I__10308 (
            .O(N__44150),
            .I(N__43874));
    Glb2LocalMux I__10307 (
            .O(N__44147),
            .I(N__43874));
    SRMux I__10306 (
            .O(N__44146),
            .I(N__43874));
    SRMux I__10305 (
            .O(N__44145),
            .I(N__43874));
    SRMux I__10304 (
            .O(N__44144),
            .I(N__43874));
    SRMux I__10303 (
            .O(N__44143),
            .I(N__43874));
    Glb2LocalMux I__10302 (
            .O(N__44140),
            .I(N__43874));
    SRMux I__10301 (
            .O(N__44139),
            .I(N__43874));
    SRMux I__10300 (
            .O(N__44138),
            .I(N__43874));
    SRMux I__10299 (
            .O(N__44137),
            .I(N__43874));
    SRMux I__10298 (
            .O(N__44136),
            .I(N__43874));
    SRMux I__10297 (
            .O(N__44135),
            .I(N__43874));
    Glb2LocalMux I__10296 (
            .O(N__44132),
            .I(N__43874));
    SRMux I__10295 (
            .O(N__44131),
            .I(N__43874));
    SRMux I__10294 (
            .O(N__44130),
            .I(N__43874));
    SRMux I__10293 (
            .O(N__44129),
            .I(N__43874));
    Glb2LocalMux I__10292 (
            .O(N__44126),
            .I(N__43874));
    SRMux I__10291 (
            .O(N__44125),
            .I(N__43874));
    SRMux I__10290 (
            .O(N__44124),
            .I(N__43874));
    SRMux I__10289 (
            .O(N__44123),
            .I(N__43874));
    SRMux I__10288 (
            .O(N__44122),
            .I(N__43874));
    SRMux I__10287 (
            .O(N__44121),
            .I(N__43874));
    SRMux I__10286 (
            .O(N__44120),
            .I(N__43874));
    SRMux I__10285 (
            .O(N__44119),
            .I(N__43874));
    SRMux I__10284 (
            .O(N__44118),
            .I(N__43874));
    SRMux I__10283 (
            .O(N__44117),
            .I(N__43874));
    SRMux I__10282 (
            .O(N__44116),
            .I(N__43874));
    SRMux I__10281 (
            .O(N__44115),
            .I(N__43874));
    SRMux I__10280 (
            .O(N__44114),
            .I(N__43874));
    SRMux I__10279 (
            .O(N__44113),
            .I(N__43874));
    SRMux I__10278 (
            .O(N__44112),
            .I(N__43874));
    SRMux I__10277 (
            .O(N__44111),
            .I(N__43874));
    SRMux I__10276 (
            .O(N__44110),
            .I(N__43874));
    SRMux I__10275 (
            .O(N__44109),
            .I(N__43874));
    SRMux I__10274 (
            .O(N__44108),
            .I(N__43874));
    SRMux I__10273 (
            .O(N__44107),
            .I(N__43874));
    SRMux I__10272 (
            .O(N__44106),
            .I(N__43874));
    SRMux I__10271 (
            .O(N__44105),
            .I(N__43874));
    SRMux I__10270 (
            .O(N__44104),
            .I(N__43874));
    SRMux I__10269 (
            .O(N__44103),
            .I(N__43874));
    GlobalMux I__10268 (
            .O(N__43874),
            .I(N__43871));
    gio2CtrlBuf I__10267 (
            .O(N__43871),
            .I(red_c_g));
    InMux I__10266 (
            .O(N__43868),
            .I(N__43865));
    LocalMux I__10265 (
            .O(N__43865),
            .I(N__43861));
    CascadeMux I__10264 (
            .O(N__43864),
            .I(N__43857));
    Span4Mux_h I__10263 (
            .O(N__43861),
            .I(N__43852));
    InMux I__10262 (
            .O(N__43860),
            .I(N__43843));
    InMux I__10261 (
            .O(N__43857),
            .I(N__43843));
    InMux I__10260 (
            .O(N__43856),
            .I(N__43843));
    InMux I__10259 (
            .O(N__43855),
            .I(N__43843));
    Odrv4 I__10258 (
            .O(N__43852),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__10257 (
            .O(N__43843),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__10256 (
            .O(N__43838),
            .I(N__43834));
    CascadeMux I__10255 (
            .O(N__43837),
            .I(N__43829));
    LocalMux I__10254 (
            .O(N__43834),
            .I(N__43823));
    CascadeMux I__10253 (
            .O(N__43833),
            .I(N__43820));
    CascadeMux I__10252 (
            .O(N__43832),
            .I(N__43816));
    InMux I__10251 (
            .O(N__43829),
            .I(N__43809));
    InMux I__10250 (
            .O(N__43828),
            .I(N__43809));
    InMux I__10249 (
            .O(N__43827),
            .I(N__43809));
    InMux I__10248 (
            .O(N__43826),
            .I(N__43806));
    Span4Mux_v I__10247 (
            .O(N__43823),
            .I(N__43803));
    InMux I__10246 (
            .O(N__43820),
            .I(N__43796));
    InMux I__10245 (
            .O(N__43819),
            .I(N__43796));
    InMux I__10244 (
            .O(N__43816),
            .I(N__43796));
    LocalMux I__10243 (
            .O(N__43809),
            .I(N__43793));
    LocalMux I__10242 (
            .O(N__43806),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__10241 (
            .O(N__43803),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__10240 (
            .O(N__43796),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__10239 (
            .O(N__43793),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    InMux I__10238 (
            .O(N__43784),
            .I(N__43781));
    LocalMux I__10237 (
            .O(N__43781),
            .I(N__43774));
    InMux I__10236 (
            .O(N__43780),
            .I(N__43765));
    InMux I__10235 (
            .O(N__43779),
            .I(N__43765));
    InMux I__10234 (
            .O(N__43778),
            .I(N__43765));
    InMux I__10233 (
            .O(N__43777),
            .I(N__43765));
    Span4Mux_v I__10232 (
            .O(N__43774),
            .I(N__43760));
    LocalMux I__10231 (
            .O(N__43765),
            .I(N__43760));
    Span4Mux_h I__10230 (
            .O(N__43760),
            .I(N__43756));
    InMux I__10229 (
            .O(N__43759),
            .I(N__43753));
    Span4Mux_h I__10228 (
            .O(N__43756),
            .I(N__43750));
    LocalMux I__10227 (
            .O(N__43753),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__10226 (
            .O(N__43750),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    CEMux I__10225 (
            .O(N__43745),
            .I(N__43740));
    CEMux I__10224 (
            .O(N__43744),
            .I(N__43737));
    CEMux I__10223 (
            .O(N__43743),
            .I(N__43732));
    LocalMux I__10222 (
            .O(N__43740),
            .I(N__43729));
    LocalMux I__10221 (
            .O(N__43737),
            .I(N__43726));
    CEMux I__10220 (
            .O(N__43736),
            .I(N__43723));
    CEMux I__10219 (
            .O(N__43735),
            .I(N__43720));
    LocalMux I__10218 (
            .O(N__43732),
            .I(N__43717));
    Span4Mux_v I__10217 (
            .O(N__43729),
            .I(N__43714));
    Span4Mux_v I__10216 (
            .O(N__43726),
            .I(N__43711));
    LocalMux I__10215 (
            .O(N__43723),
            .I(N__43708));
    LocalMux I__10214 (
            .O(N__43720),
            .I(N__43705));
    Span4Mux_h I__10213 (
            .O(N__43717),
            .I(N__43702));
    Span4Mux_v I__10212 (
            .O(N__43714),
            .I(N__43699));
    Span4Mux_v I__10211 (
            .O(N__43711),
            .I(N__43694));
    Span4Mux_h I__10210 (
            .O(N__43708),
            .I(N__43694));
    Span4Mux_v I__10209 (
            .O(N__43705),
            .I(N__43691));
    Odrv4 I__10208 (
            .O(N__43702),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0 ));
    Odrv4 I__10207 (
            .O(N__43699),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0 ));
    Odrv4 I__10206 (
            .O(N__43694),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0 ));
    Odrv4 I__10205 (
            .O(N__43691),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0 ));
    InMux I__10204 (
            .O(N__43682),
            .I(N__43678));
    InMux I__10203 (
            .O(N__43681),
            .I(N__43675));
    LocalMux I__10202 (
            .O(N__43678),
            .I(N__43672));
    LocalMux I__10201 (
            .O(N__43675),
            .I(N__43668));
    Span4Mux_v I__10200 (
            .O(N__43672),
            .I(N__43665));
    InMux I__10199 (
            .O(N__43671),
            .I(N__43662));
    Span4Mux_h I__10198 (
            .O(N__43668),
            .I(N__43659));
    Span4Mux_h I__10197 (
            .O(N__43665),
            .I(N__43656));
    LocalMux I__10196 (
            .O(N__43662),
            .I(N__43651));
    Span4Mux_v I__10195 (
            .O(N__43659),
            .I(N__43651));
    Odrv4 I__10194 (
            .O(N__43656),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__10193 (
            .O(N__43651),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__10192 (
            .O(N__43646),
            .I(N__43643));
    InMux I__10191 (
            .O(N__43643),
            .I(N__43640));
    LocalMux I__10190 (
            .O(N__43640),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    InMux I__10189 (
            .O(N__43637),
            .I(N__43633));
    InMux I__10188 (
            .O(N__43636),
            .I(N__43630));
    LocalMux I__10187 (
            .O(N__43633),
            .I(N__43627));
    LocalMux I__10186 (
            .O(N__43630),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__10185 (
            .O(N__43627),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__10184 (
            .O(N__43622),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ));
    CascadeMux I__10183 (
            .O(N__43619),
            .I(N__43616));
    InMux I__10182 (
            .O(N__43616),
            .I(N__43613));
    LocalMux I__10181 (
            .O(N__43613),
            .I(N__43610));
    Odrv4 I__10180 (
            .O(N__43610),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84ADZ0 ));
    InMux I__10179 (
            .O(N__43607),
            .I(N__43603));
    InMux I__10178 (
            .O(N__43606),
            .I(N__43600));
    LocalMux I__10177 (
            .O(N__43603),
            .I(N__43597));
    LocalMux I__10176 (
            .O(N__43600),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__10175 (
            .O(N__43597),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__10174 (
            .O(N__43592),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__10173 (
            .O(N__43589),
            .I(N__43585));
    InMux I__10172 (
            .O(N__43588),
            .I(N__43582));
    LocalMux I__10171 (
            .O(N__43585),
            .I(N__43579));
    LocalMux I__10170 (
            .O(N__43582),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__10169 (
            .O(N__43579),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__10168 (
            .O(N__43574),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__10167 (
            .O(N__43571),
            .I(N__43568));
    LocalMux I__10166 (
            .O(N__43568),
            .I(N__43565));
    Span4Mux_v I__10165 (
            .O(N__43565),
            .I(N__43562));
    Odrv4 I__10164 (
            .O(N__43562),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__10163 (
            .O(N__43559),
            .I(N__43556));
    InMux I__10162 (
            .O(N__43556),
            .I(N__43553));
    LocalMux I__10161 (
            .O(N__43553),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__10160 (
            .O(N__43550),
            .I(N__43547));
    LocalMux I__10159 (
            .O(N__43547),
            .I(N__43544));
    Span4Mux_v I__10158 (
            .O(N__43544),
            .I(N__43541));
    Odrv4 I__10157 (
            .O(N__43541),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__10156 (
            .O(N__43538),
            .I(N__43535));
    InMux I__10155 (
            .O(N__43535),
            .I(N__43532));
    LocalMux I__10154 (
            .O(N__43532),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__10153 (
            .O(N__43529),
            .I(N__43526));
    LocalMux I__10152 (
            .O(N__43526),
            .I(N__43523));
    Odrv12 I__10151 (
            .O(N__43523),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__10150 (
            .O(N__43520),
            .I(N__43517));
    InMux I__10149 (
            .O(N__43517),
            .I(N__43514));
    LocalMux I__10148 (
            .O(N__43514),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__10147 (
            .O(N__43511),
            .I(N__43508));
    LocalMux I__10146 (
            .O(N__43508),
            .I(N__43505));
    Span4Mux_v I__10145 (
            .O(N__43505),
            .I(N__43502));
    Odrv4 I__10144 (
            .O(N__43502),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__10143 (
            .O(N__43499),
            .I(N__43496));
    InMux I__10142 (
            .O(N__43496),
            .I(N__43493));
    LocalMux I__10141 (
            .O(N__43493),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__10140 (
            .O(N__43490),
            .I(N__43487));
    InMux I__10139 (
            .O(N__43487),
            .I(N__43484));
    LocalMux I__10138 (
            .O(N__43484),
            .I(N__43481));
    Span4Mux_h I__10137 (
            .O(N__43481),
            .I(N__43478));
    Odrv4 I__10136 (
            .O(N__43478),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    InMux I__10135 (
            .O(N__43475),
            .I(N__43472));
    LocalMux I__10134 (
            .O(N__43472),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ));
    InMux I__10133 (
            .O(N__43469),
            .I(N__43466));
    LocalMux I__10132 (
            .O(N__43466),
            .I(N__43463));
    Span4Mux_h I__10131 (
            .O(N__43463),
            .I(N__43460));
    Odrv4 I__10130 (
            .O(N__43460),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__10129 (
            .O(N__43457),
            .I(N__43454));
    InMux I__10128 (
            .O(N__43454),
            .I(N__43451));
    LocalMux I__10127 (
            .O(N__43451),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ));
    InMux I__10126 (
            .O(N__43448),
            .I(N__43445));
    LocalMux I__10125 (
            .O(N__43445),
            .I(N__43442));
    Odrv12 I__10124 (
            .O(N__43442),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__10123 (
            .O(N__43439),
            .I(N__43436));
    InMux I__10122 (
            .O(N__43436),
            .I(N__43433));
    LocalMux I__10121 (
            .O(N__43433),
            .I(N__43430));
    Odrv4 I__10120 (
            .O(N__43430),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ));
    InMux I__10119 (
            .O(N__43427),
            .I(N__43424));
    LocalMux I__10118 (
            .O(N__43424),
            .I(N__43421));
    Span4Mux_v I__10117 (
            .O(N__43421),
            .I(N__43418));
    Odrv4 I__10116 (
            .O(N__43418),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__10115 (
            .O(N__43415),
            .I(N__43412));
    InMux I__10114 (
            .O(N__43412),
            .I(N__43409));
    LocalMux I__10113 (
            .O(N__43409),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ));
    CascadeMux I__10112 (
            .O(N__43406),
            .I(N__43403));
    InMux I__10111 (
            .O(N__43403),
            .I(N__43400));
    LocalMux I__10110 (
            .O(N__43400),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__10109 (
            .O(N__43397),
            .I(N__43394));
    InMux I__10108 (
            .O(N__43394),
            .I(N__43391));
    LocalMux I__10107 (
            .O(N__43391),
            .I(N__43388));
    Odrv4 I__10106 (
            .O(N__43388),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    InMux I__10105 (
            .O(N__43385),
            .I(N__43382));
    LocalMux I__10104 (
            .O(N__43382),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__10103 (
            .O(N__43379),
            .I(N__43376));
    LocalMux I__10102 (
            .O(N__43376),
            .I(N__43373));
    Span4Mux_h I__10101 (
            .O(N__43373),
            .I(N__43370));
    Odrv4 I__10100 (
            .O(N__43370),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__10099 (
            .O(N__43367),
            .I(N__43364));
    InMux I__10098 (
            .O(N__43364),
            .I(N__43361));
    LocalMux I__10097 (
            .O(N__43361),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__10096 (
            .O(N__43358),
            .I(N__43355));
    LocalMux I__10095 (
            .O(N__43355),
            .I(N__43352));
    Span4Mux_h I__10094 (
            .O(N__43352),
            .I(N__43349));
    Odrv4 I__10093 (
            .O(N__43349),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__10092 (
            .O(N__43346),
            .I(N__43343));
    InMux I__10091 (
            .O(N__43343),
            .I(N__43340));
    LocalMux I__10090 (
            .O(N__43340),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    InMux I__10089 (
            .O(N__43337),
            .I(N__43334));
    LocalMux I__10088 (
            .O(N__43334),
            .I(N__43331));
    Span4Mux_v I__10087 (
            .O(N__43331),
            .I(N__43328));
    Odrv4 I__10086 (
            .O(N__43328),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__10085 (
            .O(N__43325),
            .I(N__43322));
    InMux I__10084 (
            .O(N__43322),
            .I(N__43319));
    LocalMux I__10083 (
            .O(N__43319),
            .I(N__43316));
    Odrv4 I__10082 (
            .O(N__43316),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__10081 (
            .O(N__43313),
            .I(N__43310));
    LocalMux I__10080 (
            .O(N__43310),
            .I(N__43307));
    Span4Mux_h I__10079 (
            .O(N__43307),
            .I(N__43304));
    Span4Mux_h I__10078 (
            .O(N__43304),
            .I(N__43301));
    Odrv4 I__10077 (
            .O(N__43301),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__10076 (
            .O(N__43298),
            .I(N__43295));
    InMux I__10075 (
            .O(N__43295),
            .I(N__43292));
    LocalMux I__10074 (
            .O(N__43292),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__10073 (
            .O(N__43289),
            .I(N__43286));
    LocalMux I__10072 (
            .O(N__43286),
            .I(N__43283));
    Odrv12 I__10071 (
            .O(N__43283),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__10070 (
            .O(N__43280),
            .I(N__43277));
    InMux I__10069 (
            .O(N__43277),
            .I(N__43274));
    LocalMux I__10068 (
            .O(N__43274),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__10067 (
            .O(N__43271),
            .I(N__43268));
    InMux I__10066 (
            .O(N__43268),
            .I(N__43265));
    LocalMux I__10065 (
            .O(N__43265),
            .I(N__43262));
    Odrv12 I__10064 (
            .O(N__43262),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    InMux I__10063 (
            .O(N__43259),
            .I(N__43256));
    LocalMux I__10062 (
            .O(N__43256),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__10061 (
            .O(N__43253),
            .I(N__43249));
    InMux I__10060 (
            .O(N__43252),
            .I(N__43246));
    LocalMux I__10059 (
            .O(N__43249),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__10058 (
            .O(N__43246),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__10057 (
            .O(N__43241),
            .I(N__43238));
    LocalMux I__10056 (
            .O(N__43238),
            .I(N__43235));
    Odrv4 I__10055 (
            .O(N__43235),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__10054 (
            .O(N__43232),
            .I(N__43229));
    InMux I__10053 (
            .O(N__43229),
            .I(N__43226));
    LocalMux I__10052 (
            .O(N__43226),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    InMux I__10051 (
            .O(N__43223),
            .I(N__43220));
    LocalMux I__10050 (
            .O(N__43220),
            .I(N__43217));
    Odrv4 I__10049 (
            .O(N__43217),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__10048 (
            .O(N__43214),
            .I(N__43210));
    InMux I__10047 (
            .O(N__43213),
            .I(N__43207));
    LocalMux I__10046 (
            .O(N__43210),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__10045 (
            .O(N__43207),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__10044 (
            .O(N__43202),
            .I(N__43199));
    InMux I__10043 (
            .O(N__43199),
            .I(N__43196));
    LocalMux I__10042 (
            .O(N__43196),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__10041 (
            .O(N__43193),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__10040 (
            .O(N__43190),
            .I(N__43185));
    InMux I__10039 (
            .O(N__43189),
            .I(N__43182));
    CascadeMux I__10038 (
            .O(N__43188),
            .I(N__43175));
    LocalMux I__10037 (
            .O(N__43185),
            .I(N__43171));
    LocalMux I__10036 (
            .O(N__43182),
            .I(N__43168));
    InMux I__10035 (
            .O(N__43181),
            .I(N__43155));
    InMux I__10034 (
            .O(N__43180),
            .I(N__43155));
    InMux I__10033 (
            .O(N__43179),
            .I(N__43155));
    InMux I__10032 (
            .O(N__43178),
            .I(N__43155));
    InMux I__10031 (
            .O(N__43175),
            .I(N__43155));
    InMux I__10030 (
            .O(N__43174),
            .I(N__43155));
    Odrv4 I__10029 (
            .O(N__43171),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv12 I__10028 (
            .O(N__43168),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__10027 (
            .O(N__43155),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    InMux I__10026 (
            .O(N__43148),
            .I(N__43145));
    LocalMux I__10025 (
            .O(N__43145),
            .I(N__43140));
    CascadeMux I__10024 (
            .O(N__43144),
            .I(N__43136));
    CascadeMux I__10023 (
            .O(N__43143),
            .I(N__43133));
    Span4Mux_v I__10022 (
            .O(N__43140),
            .I(N__43128));
    InMux I__10021 (
            .O(N__43139),
            .I(N__43119));
    InMux I__10020 (
            .O(N__43136),
            .I(N__43119));
    InMux I__10019 (
            .O(N__43133),
            .I(N__43119));
    InMux I__10018 (
            .O(N__43132),
            .I(N__43119));
    InMux I__10017 (
            .O(N__43131),
            .I(N__43116));
    Sp12to4 I__10016 (
            .O(N__43128),
            .I(N__43111));
    LocalMux I__10015 (
            .O(N__43119),
            .I(N__43111));
    LocalMux I__10014 (
            .O(N__43116),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__10013 (
            .O(N__43111),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__10012 (
            .O(N__43106),
            .I(N__43103));
    LocalMux I__10011 (
            .O(N__43103),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0 ));
    CascadeMux I__10010 (
            .O(N__43100),
            .I(N__43097));
    InMux I__10009 (
            .O(N__43097),
            .I(N__43094));
    LocalMux I__10008 (
            .O(N__43094),
            .I(N__43091));
    Span4Mux_v I__10007 (
            .O(N__43091),
            .I(N__43088));
    Odrv4 I__10006 (
            .O(N__43088),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    InMux I__10005 (
            .O(N__43085),
            .I(N__43082));
    LocalMux I__10004 (
            .O(N__43082),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    InMux I__10003 (
            .O(N__43079),
            .I(N__43076));
    LocalMux I__10002 (
            .O(N__43076),
            .I(N__43073));
    Odrv4 I__10001 (
            .O(N__43073),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__10000 (
            .O(N__43070),
            .I(N__43067));
    InMux I__9999 (
            .O(N__43067),
            .I(N__43064));
    LocalMux I__9998 (
            .O(N__43064),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    InMux I__9997 (
            .O(N__43061),
            .I(N__43058));
    LocalMux I__9996 (
            .O(N__43058),
            .I(N__43055));
    Span4Mux_v I__9995 (
            .O(N__43055),
            .I(N__43052));
    Odrv4 I__9994 (
            .O(N__43052),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__9993 (
            .O(N__43049),
            .I(N__43046));
    InMux I__9992 (
            .O(N__43046),
            .I(N__43043));
    LocalMux I__9991 (
            .O(N__43043),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__9990 (
            .O(N__43040),
            .I(N__43037));
    LocalMux I__9989 (
            .O(N__43037),
            .I(N__43034));
    Odrv12 I__9988 (
            .O(N__43034),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    InMux I__9987 (
            .O(N__43031),
            .I(N__43027));
    InMux I__9986 (
            .O(N__43030),
            .I(N__43024));
    LocalMux I__9985 (
            .O(N__43027),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__9984 (
            .O(N__43024),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__9983 (
            .O(N__43019),
            .I(N__43016));
    LocalMux I__9982 (
            .O(N__43016),
            .I(N__43013));
    Odrv4 I__9981 (
            .O(N__43013),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__9980 (
            .O(N__43010),
            .I(N__43007));
    InMux I__9979 (
            .O(N__43007),
            .I(N__43004));
    LocalMux I__9978 (
            .O(N__43004),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__9977 (
            .O(N__43001),
            .I(N__42998));
    LocalMux I__9976 (
            .O(N__42998),
            .I(N__42995));
    Odrv4 I__9975 (
            .O(N__42995),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__9974 (
            .O(N__42992),
            .I(N__42988));
    InMux I__9973 (
            .O(N__42991),
            .I(N__42985));
    LocalMux I__9972 (
            .O(N__42988),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__9971 (
            .O(N__42985),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    CascadeMux I__9970 (
            .O(N__42980),
            .I(N__42977));
    InMux I__9969 (
            .O(N__42977),
            .I(N__42974));
    LocalMux I__9968 (
            .O(N__42974),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__9967 (
            .O(N__42971),
            .I(N__42968));
    LocalMux I__9966 (
            .O(N__42968),
            .I(N__42965));
    Span4Mux_v I__9965 (
            .O(N__42965),
            .I(N__42962));
    Odrv4 I__9964 (
            .O(N__42962),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    InMux I__9963 (
            .O(N__42959),
            .I(N__42955));
    InMux I__9962 (
            .O(N__42958),
            .I(N__42952));
    LocalMux I__9961 (
            .O(N__42955),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__9960 (
            .O(N__42952),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    CascadeMux I__9959 (
            .O(N__42947),
            .I(N__42944));
    InMux I__9958 (
            .O(N__42944),
            .I(N__42941));
    LocalMux I__9957 (
            .O(N__42941),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__9956 (
            .O(N__42938),
            .I(N__42935));
    InMux I__9955 (
            .O(N__42935),
            .I(N__42932));
    LocalMux I__9954 (
            .O(N__42932),
            .I(N__42929));
    Odrv4 I__9953 (
            .O(N__42929),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__9952 (
            .O(N__42926),
            .I(N__42922));
    InMux I__9951 (
            .O(N__42925),
            .I(N__42919));
    LocalMux I__9950 (
            .O(N__42922),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__9949 (
            .O(N__42919),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__9948 (
            .O(N__42914),
            .I(N__42911));
    LocalMux I__9947 (
            .O(N__42911),
            .I(N__42908));
    Odrv4 I__9946 (
            .O(N__42908),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__9945 (
            .O(N__42905),
            .I(N__42902));
    LocalMux I__9944 (
            .O(N__42902),
            .I(N__42899));
    Odrv4 I__9943 (
            .O(N__42899),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__9942 (
            .O(N__42896),
            .I(N__42892));
    InMux I__9941 (
            .O(N__42895),
            .I(N__42889));
    LocalMux I__9940 (
            .O(N__42892),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__9939 (
            .O(N__42889),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__9938 (
            .O(N__42884),
            .I(N__42881));
    InMux I__9937 (
            .O(N__42881),
            .I(N__42878));
    LocalMux I__9936 (
            .O(N__42878),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__9935 (
            .O(N__42875),
            .I(N__42872));
    InMux I__9934 (
            .O(N__42872),
            .I(N__42869));
    LocalMux I__9933 (
            .O(N__42869),
            .I(N__42866));
    Span4Mux_h I__9932 (
            .O(N__42866),
            .I(N__42863));
    Odrv4 I__9931 (
            .O(N__42863),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__9930 (
            .O(N__42860),
            .I(N__42856));
    InMux I__9929 (
            .O(N__42859),
            .I(N__42853));
    LocalMux I__9928 (
            .O(N__42856),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__9927 (
            .O(N__42853),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__9926 (
            .O(N__42848),
            .I(N__42845));
    LocalMux I__9925 (
            .O(N__42845),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__9924 (
            .O(N__42842),
            .I(N__42838));
    InMux I__9923 (
            .O(N__42841),
            .I(N__42835));
    LocalMux I__9922 (
            .O(N__42838),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__9921 (
            .O(N__42835),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__9920 (
            .O(N__42830),
            .I(N__42827));
    LocalMux I__9919 (
            .O(N__42827),
            .I(N__42824));
    Odrv4 I__9918 (
            .O(N__42824),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__9917 (
            .O(N__42821),
            .I(N__42818));
    InMux I__9916 (
            .O(N__42818),
            .I(N__42815));
    LocalMux I__9915 (
            .O(N__42815),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    CascadeMux I__9914 (
            .O(N__42812),
            .I(N__42809));
    InMux I__9913 (
            .O(N__42809),
            .I(N__42806));
    LocalMux I__9912 (
            .O(N__42806),
            .I(N__42803));
    Odrv12 I__9911 (
            .O(N__42803),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__9910 (
            .O(N__42800),
            .I(N__42796));
    InMux I__9909 (
            .O(N__42799),
            .I(N__42793));
    LocalMux I__9908 (
            .O(N__42796),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__9907 (
            .O(N__42793),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__9906 (
            .O(N__42788),
            .I(N__42785));
    LocalMux I__9905 (
            .O(N__42785),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    CascadeMux I__9904 (
            .O(N__42782),
            .I(N__42779));
    InMux I__9903 (
            .O(N__42779),
            .I(N__42776));
    LocalMux I__9902 (
            .O(N__42776),
            .I(N__42773));
    Span4Mux_h I__9901 (
            .O(N__42773),
            .I(N__42770));
    Span4Mux_v I__9900 (
            .O(N__42770),
            .I(N__42767));
    Odrv4 I__9899 (
            .O(N__42767),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__9898 (
            .O(N__42764),
            .I(N__42761));
    InMux I__9897 (
            .O(N__42761),
            .I(N__42757));
    InMux I__9896 (
            .O(N__42760),
            .I(N__42754));
    LocalMux I__9895 (
            .O(N__42757),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__9894 (
            .O(N__42754),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__9893 (
            .O(N__42749),
            .I(N__42746));
    LocalMux I__9892 (
            .O(N__42746),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__9891 (
            .O(N__42743),
            .I(N__42740));
    LocalMux I__9890 (
            .O(N__42740),
            .I(N__42737));
    Span4Mux_h I__9889 (
            .O(N__42737),
            .I(N__42734));
    Span4Mux_v I__9888 (
            .O(N__42734),
            .I(N__42731));
    Odrv4 I__9887 (
            .O(N__42731),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__9886 (
            .O(N__42728),
            .I(N__42724));
    InMux I__9885 (
            .O(N__42727),
            .I(N__42721));
    LocalMux I__9884 (
            .O(N__42724),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__9883 (
            .O(N__42721),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    CascadeMux I__9882 (
            .O(N__42716),
            .I(N__42713));
    InMux I__9881 (
            .O(N__42713),
            .I(N__42710));
    LocalMux I__9880 (
            .O(N__42710),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__9879 (
            .O(N__42707),
            .I(N__42704));
    LocalMux I__9878 (
            .O(N__42704),
            .I(N__42701));
    Span4Mux_v I__9877 (
            .O(N__42701),
            .I(N__42698));
    Odrv4 I__9876 (
            .O(N__42698),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__9875 (
            .O(N__42695),
            .I(N__42691));
    InMux I__9874 (
            .O(N__42694),
            .I(N__42688));
    LocalMux I__9873 (
            .O(N__42691),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__9872 (
            .O(N__42688),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    CascadeMux I__9871 (
            .O(N__42683),
            .I(N__42680));
    InMux I__9870 (
            .O(N__42680),
            .I(N__42677));
    LocalMux I__9869 (
            .O(N__42677),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__9868 (
            .O(N__42674),
            .I(N__42671));
    LocalMux I__9867 (
            .O(N__42671),
            .I(N__42668));
    Span4Mux_h I__9866 (
            .O(N__42668),
            .I(N__42665));
    Odrv4 I__9865 (
            .O(N__42665),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    InMux I__9864 (
            .O(N__42662),
            .I(N__42658));
    InMux I__9863 (
            .O(N__42661),
            .I(N__42655));
    LocalMux I__9862 (
            .O(N__42658),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__9861 (
            .O(N__42655),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__9860 (
            .O(N__42650),
            .I(N__42647));
    InMux I__9859 (
            .O(N__42647),
            .I(N__42644));
    LocalMux I__9858 (
            .O(N__42644),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__9857 (
            .O(N__42641),
            .I(N__42638));
    LocalMux I__9856 (
            .O(N__42638),
            .I(N__42635));
    Span4Mux_v I__9855 (
            .O(N__42635),
            .I(N__42632));
    Odrv4 I__9854 (
            .O(N__42632),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__9853 (
            .O(N__42629),
            .I(N__42625));
    InMux I__9852 (
            .O(N__42628),
            .I(N__42622));
    LocalMux I__9851 (
            .O(N__42625),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__9850 (
            .O(N__42622),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__9849 (
            .O(N__42617),
            .I(N__42614));
    InMux I__9848 (
            .O(N__42614),
            .I(N__42611));
    LocalMux I__9847 (
            .O(N__42611),
            .I(N__42608));
    Odrv4 I__9846 (
            .O(N__42608),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__9845 (
            .O(N__42605),
            .I(N__42601));
    InMux I__9844 (
            .O(N__42604),
            .I(N__42598));
    LocalMux I__9843 (
            .O(N__42601),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__9842 (
            .O(N__42598),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__9841 (
            .O(N__42593),
            .I(N__42590));
    LocalMux I__9840 (
            .O(N__42590),
            .I(N__42587));
    Span4Mux_h I__9839 (
            .O(N__42587),
            .I(N__42584));
    Odrv4 I__9838 (
            .O(N__42584),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__9837 (
            .O(N__42581),
            .I(N__42578));
    InMux I__9836 (
            .O(N__42578),
            .I(N__42575));
    LocalMux I__9835 (
            .O(N__42575),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__9834 (
            .O(N__42572),
            .I(N__42569));
    LocalMux I__9833 (
            .O(N__42569),
            .I(N__42566));
    Span4Mux_v I__9832 (
            .O(N__42566),
            .I(N__42563));
    Odrv4 I__9831 (
            .O(N__42563),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__9830 (
            .O(N__42560),
            .I(N__42556));
    InMux I__9829 (
            .O(N__42559),
            .I(N__42553));
    LocalMux I__9828 (
            .O(N__42556),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__9827 (
            .O(N__42553),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__9826 (
            .O(N__42548),
            .I(N__42545));
    InMux I__9825 (
            .O(N__42545),
            .I(N__42542));
    LocalMux I__9824 (
            .O(N__42542),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__9823 (
            .O(N__42539),
            .I(N__42536));
    InMux I__9822 (
            .O(N__42536),
            .I(N__42531));
    CascadeMux I__9821 (
            .O(N__42535),
            .I(N__42528));
    InMux I__9820 (
            .O(N__42534),
            .I(N__42525));
    LocalMux I__9819 (
            .O(N__42531),
            .I(N__42522));
    InMux I__9818 (
            .O(N__42528),
            .I(N__42518));
    LocalMux I__9817 (
            .O(N__42525),
            .I(N__42515));
    Span4Mux_h I__9816 (
            .O(N__42522),
            .I(N__42512));
    InMux I__9815 (
            .O(N__42521),
            .I(N__42509));
    LocalMux I__9814 (
            .O(N__42518),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    Odrv12 I__9813 (
            .O(N__42515),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    Odrv4 I__9812 (
            .O(N__42512),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    LocalMux I__9811 (
            .O(N__42509),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    InMux I__9810 (
            .O(N__42500),
            .I(N__42495));
    InMux I__9809 (
            .O(N__42499),
            .I(N__42489));
    InMux I__9808 (
            .O(N__42498),
            .I(N__42489));
    LocalMux I__9807 (
            .O(N__42495),
            .I(N__42485));
    InMux I__9806 (
            .O(N__42494),
            .I(N__42482));
    LocalMux I__9805 (
            .O(N__42489),
            .I(N__42479));
    InMux I__9804 (
            .O(N__42488),
            .I(N__42476));
    Span4Mux_v I__9803 (
            .O(N__42485),
            .I(N__42473));
    LocalMux I__9802 (
            .O(N__42482),
            .I(N__42470));
    Span4Mux_h I__9801 (
            .O(N__42479),
            .I(N__42467));
    LocalMux I__9800 (
            .O(N__42476),
            .I(elapsed_time_ns_1_RNIFG4DM1_0_16));
    Odrv4 I__9799 (
            .O(N__42473),
            .I(elapsed_time_ns_1_RNIFG4DM1_0_16));
    Odrv12 I__9798 (
            .O(N__42470),
            .I(elapsed_time_ns_1_RNIFG4DM1_0_16));
    Odrv4 I__9797 (
            .O(N__42467),
            .I(elapsed_time_ns_1_RNIFG4DM1_0_16));
    InMux I__9796 (
            .O(N__42458),
            .I(N__42441));
    InMux I__9795 (
            .O(N__42457),
            .I(N__42441));
    InMux I__9794 (
            .O(N__42456),
            .I(N__42441));
    InMux I__9793 (
            .O(N__42455),
            .I(N__42441));
    InMux I__9792 (
            .O(N__42454),
            .I(N__42430));
    InMux I__9791 (
            .O(N__42453),
            .I(N__42430));
    InMux I__9790 (
            .O(N__42452),
            .I(N__42430));
    InMux I__9789 (
            .O(N__42451),
            .I(N__42430));
    InMux I__9788 (
            .O(N__42450),
            .I(N__42430));
    LocalMux I__9787 (
            .O(N__42441),
            .I(N__42424));
    LocalMux I__9786 (
            .O(N__42430),
            .I(N__42424));
    InMux I__9785 (
            .O(N__42429),
            .I(N__42421));
    Span4Mux_v I__9784 (
            .O(N__42424),
            .I(N__42418));
    LocalMux I__9783 (
            .O(N__42421),
            .I(\phase_controller_inst1.stoper_tr.N_241 ));
    Odrv4 I__9782 (
            .O(N__42418),
            .I(\phase_controller_inst1.stoper_tr.N_241 ));
    CascadeMux I__9781 (
            .O(N__42413),
            .I(N__42409));
    InMux I__9780 (
            .O(N__42412),
            .I(N__42406));
    InMux I__9779 (
            .O(N__42409),
            .I(N__42403));
    LocalMux I__9778 (
            .O(N__42406),
            .I(N__42400));
    LocalMux I__9777 (
            .O(N__42403),
            .I(N__42397));
    Span4Mux_h I__9776 (
            .O(N__42400),
            .I(N__42393));
    Span4Mux_v I__9775 (
            .O(N__42397),
            .I(N__42390));
    InMux I__9774 (
            .O(N__42396),
            .I(N__42387));
    Odrv4 I__9773 (
            .O(N__42393),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    Odrv4 I__9772 (
            .O(N__42390),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    LocalMux I__9771 (
            .O(N__42387),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    InMux I__9770 (
            .O(N__42380),
            .I(N__42376));
    InMux I__9769 (
            .O(N__42379),
            .I(N__42373));
    LocalMux I__9768 (
            .O(N__42376),
            .I(N__42366));
    LocalMux I__9767 (
            .O(N__42373),
            .I(N__42366));
    CascadeMux I__9766 (
            .O(N__42372),
            .I(N__42362));
    InMux I__9765 (
            .O(N__42371),
            .I(N__42359));
    Span4Mux_v I__9764 (
            .O(N__42366),
            .I(N__42356));
    InMux I__9763 (
            .O(N__42365),
            .I(N__42351));
    InMux I__9762 (
            .O(N__42362),
            .I(N__42351));
    LocalMux I__9761 (
            .O(N__42359),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19));
    Odrv4 I__9760 (
            .O(N__42356),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19));
    LocalMux I__9759 (
            .O(N__42351),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19));
    InMux I__9758 (
            .O(N__42344),
            .I(N__42340));
    InMux I__9757 (
            .O(N__42343),
            .I(N__42337));
    LocalMux I__9756 (
            .O(N__42340),
            .I(N__42334));
    LocalMux I__9755 (
            .O(N__42337),
            .I(N__42331));
    Span4Mux_h I__9754 (
            .O(N__42334),
            .I(N__42325));
    Span4Mux_v I__9753 (
            .O(N__42331),
            .I(N__42325));
    InMux I__9752 (
            .O(N__42330),
            .I(N__42320));
    Span4Mux_h I__9751 (
            .O(N__42325),
            .I(N__42317));
    InMux I__9750 (
            .O(N__42324),
            .I(N__42312));
    InMux I__9749 (
            .O(N__42323),
            .I(N__42312));
    LocalMux I__9748 (
            .O(N__42320),
            .I(elapsed_time_ns_1_RNIHI4DM1_0_18));
    Odrv4 I__9747 (
            .O(N__42317),
            .I(elapsed_time_ns_1_RNIHI4DM1_0_18));
    LocalMux I__9746 (
            .O(N__42312),
            .I(elapsed_time_ns_1_RNIHI4DM1_0_18));
    InMux I__9745 (
            .O(N__42305),
            .I(N__42300));
    InMux I__9744 (
            .O(N__42304),
            .I(N__42297));
    InMux I__9743 (
            .O(N__42303),
            .I(N__42294));
    LocalMux I__9742 (
            .O(N__42300),
            .I(N__42291));
    LocalMux I__9741 (
            .O(N__42297),
            .I(N__42286));
    LocalMux I__9740 (
            .O(N__42294),
            .I(N__42281));
    Span4Mux_h I__9739 (
            .O(N__42291),
            .I(N__42281));
    InMux I__9738 (
            .O(N__42290),
            .I(N__42276));
    InMux I__9737 (
            .O(N__42289),
            .I(N__42276));
    Odrv4 I__9736 (
            .O(N__42286),
            .I(elapsed_time_ns_1_RNIGH4DM1_0_17));
    Odrv4 I__9735 (
            .O(N__42281),
            .I(elapsed_time_ns_1_RNIGH4DM1_0_17));
    LocalMux I__9734 (
            .O(N__42276),
            .I(elapsed_time_ns_1_RNIGH4DM1_0_17));
    CascadeMux I__9733 (
            .O(N__42269),
            .I(N__42261));
    CascadeMux I__9732 (
            .O(N__42268),
            .I(N__42257));
    CascadeMux I__9731 (
            .O(N__42267),
            .I(N__42253));
    InMux I__9730 (
            .O(N__42266),
            .I(N__42233));
    InMux I__9729 (
            .O(N__42265),
            .I(N__42233));
    InMux I__9728 (
            .O(N__42264),
            .I(N__42233));
    InMux I__9727 (
            .O(N__42261),
            .I(N__42233));
    InMux I__9726 (
            .O(N__42260),
            .I(N__42233));
    InMux I__9725 (
            .O(N__42257),
            .I(N__42228));
    InMux I__9724 (
            .O(N__42256),
            .I(N__42228));
    InMux I__9723 (
            .O(N__42253),
            .I(N__42222));
    InMux I__9722 (
            .O(N__42252),
            .I(N__42222));
    InMux I__9721 (
            .O(N__42251),
            .I(N__42215));
    InMux I__9720 (
            .O(N__42250),
            .I(N__42215));
    InMux I__9719 (
            .O(N__42249),
            .I(N__42215));
    InMux I__9718 (
            .O(N__42248),
            .I(N__42204));
    InMux I__9717 (
            .O(N__42247),
            .I(N__42204));
    InMux I__9716 (
            .O(N__42246),
            .I(N__42204));
    InMux I__9715 (
            .O(N__42245),
            .I(N__42204));
    InMux I__9714 (
            .O(N__42244),
            .I(N__42204));
    LocalMux I__9713 (
            .O(N__42233),
            .I(N__42199));
    LocalMux I__9712 (
            .O(N__42228),
            .I(N__42199));
    CascadeMux I__9711 (
            .O(N__42227),
            .I(N__42191));
    LocalMux I__9710 (
            .O(N__42222),
            .I(N__42176));
    LocalMux I__9709 (
            .O(N__42215),
            .I(N__42171));
    LocalMux I__9708 (
            .O(N__42204),
            .I(N__42171));
    Span4Mux_h I__9707 (
            .O(N__42199),
            .I(N__42168));
    InMux I__9706 (
            .O(N__42198),
            .I(N__42158));
    InMux I__9705 (
            .O(N__42197),
            .I(N__42158));
    InMux I__9704 (
            .O(N__42196),
            .I(N__42158));
    InMux I__9703 (
            .O(N__42195),
            .I(N__42141));
    InMux I__9702 (
            .O(N__42194),
            .I(N__42141));
    InMux I__9701 (
            .O(N__42191),
            .I(N__42141));
    InMux I__9700 (
            .O(N__42190),
            .I(N__42141));
    InMux I__9699 (
            .O(N__42189),
            .I(N__42141));
    InMux I__9698 (
            .O(N__42188),
            .I(N__42141));
    InMux I__9697 (
            .O(N__42187),
            .I(N__42141));
    InMux I__9696 (
            .O(N__42186),
            .I(N__42141));
    InMux I__9695 (
            .O(N__42185),
            .I(N__42126));
    InMux I__9694 (
            .O(N__42184),
            .I(N__42126));
    InMux I__9693 (
            .O(N__42183),
            .I(N__42126));
    InMux I__9692 (
            .O(N__42182),
            .I(N__42126));
    InMux I__9691 (
            .O(N__42181),
            .I(N__42126));
    InMux I__9690 (
            .O(N__42180),
            .I(N__42126));
    InMux I__9689 (
            .O(N__42179),
            .I(N__42126));
    Span4Mux_v I__9688 (
            .O(N__42176),
            .I(N__42123));
    Span4Mux_h I__9687 (
            .O(N__42171),
            .I(N__42120));
    Span4Mux_v I__9686 (
            .O(N__42168),
            .I(N__42117));
    InMux I__9685 (
            .O(N__42167),
            .I(N__42114));
    InMux I__9684 (
            .O(N__42166),
            .I(N__42109));
    InMux I__9683 (
            .O(N__42165),
            .I(N__42109));
    LocalMux I__9682 (
            .O(N__42158),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__9681 (
            .O(N__42141),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__9680 (
            .O(N__42126),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__9679 (
            .O(N__42123),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__9678 (
            .O(N__42120),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__9677 (
            .O(N__42117),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__9676 (
            .O(N__42114),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__9675 (
            .O(N__42109),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    CascadeMux I__9674 (
            .O(N__42092),
            .I(N__42082));
    CascadeMux I__9673 (
            .O(N__42091),
            .I(N__42079));
    CascadeMux I__9672 (
            .O(N__42090),
            .I(N__42076));
    CascadeMux I__9671 (
            .O(N__42089),
            .I(N__42063));
    InMux I__9670 (
            .O(N__42088),
            .I(N__42043));
    InMux I__9669 (
            .O(N__42087),
            .I(N__42043));
    InMux I__9668 (
            .O(N__42086),
            .I(N__42043));
    InMux I__9667 (
            .O(N__42085),
            .I(N__42043));
    InMux I__9666 (
            .O(N__42082),
            .I(N__42043));
    InMux I__9665 (
            .O(N__42079),
            .I(N__42043));
    InMux I__9664 (
            .O(N__42076),
            .I(N__42043));
    InMux I__9663 (
            .O(N__42075),
            .I(N__42043));
    CascadeMux I__9662 (
            .O(N__42074),
            .I(N__42039));
    InMux I__9661 (
            .O(N__42073),
            .I(N__42029));
    InMux I__9660 (
            .O(N__42072),
            .I(N__42029));
    InMux I__9659 (
            .O(N__42071),
            .I(N__42029));
    InMux I__9658 (
            .O(N__42070),
            .I(N__42029));
    InMux I__9657 (
            .O(N__42069),
            .I(N__42026));
    InMux I__9656 (
            .O(N__42068),
            .I(N__42010));
    InMux I__9655 (
            .O(N__42067),
            .I(N__42010));
    InMux I__9654 (
            .O(N__42066),
            .I(N__42010));
    InMux I__9653 (
            .O(N__42063),
            .I(N__42010));
    InMux I__9652 (
            .O(N__42062),
            .I(N__42010));
    InMux I__9651 (
            .O(N__42061),
            .I(N__42010));
    InMux I__9650 (
            .O(N__42060),
            .I(N__42010));
    LocalMux I__9649 (
            .O(N__42043),
            .I(N__42003));
    InMux I__9648 (
            .O(N__42042),
            .I(N__41996));
    InMux I__9647 (
            .O(N__42039),
            .I(N__41996));
    InMux I__9646 (
            .O(N__42038),
            .I(N__41996));
    LocalMux I__9645 (
            .O(N__42029),
            .I(N__41993));
    LocalMux I__9644 (
            .O(N__42026),
            .I(N__41990));
    InMux I__9643 (
            .O(N__42025),
            .I(N__41987));
    LocalMux I__9642 (
            .O(N__42010),
            .I(N__41984));
    InMux I__9641 (
            .O(N__42009),
            .I(N__41981));
    InMux I__9640 (
            .O(N__42008),
            .I(N__41978));
    InMux I__9639 (
            .O(N__42007),
            .I(N__41973));
    InMux I__9638 (
            .O(N__42006),
            .I(N__41973));
    Span4Mux_h I__9637 (
            .O(N__42003),
            .I(N__41970));
    LocalMux I__9636 (
            .O(N__41996),
            .I(N__41961));
    Span4Mux_v I__9635 (
            .O(N__41993),
            .I(N__41961));
    Span4Mux_h I__9634 (
            .O(N__41990),
            .I(N__41961));
    LocalMux I__9633 (
            .O(N__41987),
            .I(N__41961));
    Span4Mux_h I__9632 (
            .O(N__41984),
            .I(N__41952));
    LocalMux I__9631 (
            .O(N__41981),
            .I(N__41952));
    LocalMux I__9630 (
            .O(N__41978),
            .I(N__41952));
    LocalMux I__9629 (
            .O(N__41973),
            .I(N__41952));
    Odrv4 I__9628 (
            .O(N__41970),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_o5_0Z0Z_15 ));
    Odrv4 I__9627 (
            .O(N__41961),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_o5_0Z0Z_15 ));
    Odrv4 I__9626 (
            .O(N__41952),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_o5_0Z0Z_15 ));
    CEMux I__9625 (
            .O(N__41945),
            .I(N__41942));
    LocalMux I__9624 (
            .O(N__41942),
            .I(N__41938));
    CEMux I__9623 (
            .O(N__41941),
            .I(N__41935));
    Span4Mux_v I__9622 (
            .O(N__41938),
            .I(N__41931));
    LocalMux I__9621 (
            .O(N__41935),
            .I(N__41928));
    CEMux I__9620 (
            .O(N__41934),
            .I(N__41925));
    Span4Mux_h I__9619 (
            .O(N__41931),
            .I(N__41920));
    Span4Mux_v I__9618 (
            .O(N__41928),
            .I(N__41920));
    LocalMux I__9617 (
            .O(N__41925),
            .I(N__41917));
    Span4Mux_v I__9616 (
            .O(N__41920),
            .I(N__41914));
    Span4Mux_h I__9615 (
            .O(N__41917),
            .I(N__41911));
    Odrv4 I__9614 (
            .O(N__41914),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa_0 ));
    Odrv4 I__9613 (
            .O(N__41911),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa_0 ));
    InMux I__9612 (
            .O(N__41906),
            .I(N__41903));
    LocalMux I__9611 (
            .O(N__41903),
            .I(N__41900));
    Span4Mux_h I__9610 (
            .O(N__41900),
            .I(N__41897));
    Span4Mux_v I__9609 (
            .O(N__41897),
            .I(N__41894));
    Span4Mux_v I__9608 (
            .O(N__41894),
            .I(N__41891));
    Odrv4 I__9607 (
            .O(N__41891),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__9606 (
            .O(N__41888),
            .I(N__41885));
    LocalMux I__9605 (
            .O(N__41885),
            .I(N__41882));
    Span4Mux_v I__9604 (
            .O(N__41882),
            .I(N__41877));
    InMux I__9603 (
            .O(N__41881),
            .I(N__41874));
    InMux I__9602 (
            .O(N__41880),
            .I(N__41871));
    Sp12to4 I__9601 (
            .O(N__41877),
            .I(N__41866));
    LocalMux I__9600 (
            .O(N__41874),
            .I(N__41866));
    LocalMux I__9599 (
            .O(N__41871),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__9598 (
            .O(N__41866),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__9597 (
            .O(N__41861),
            .I(N__41858));
    InMux I__9596 (
            .O(N__41858),
            .I(N__41855));
    LocalMux I__9595 (
            .O(N__41855),
            .I(N__41852));
    Odrv4 I__9594 (
            .O(N__41852),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__9593 (
            .O(N__41849),
            .I(N__41845));
    InMux I__9592 (
            .O(N__41848),
            .I(N__41842));
    LocalMux I__9591 (
            .O(N__41845),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__9590 (
            .O(N__41842),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__9589 (
            .O(N__41837),
            .I(N__41834));
    LocalMux I__9588 (
            .O(N__41834),
            .I(N__41831));
    Span4Mux_h I__9587 (
            .O(N__41831),
            .I(N__41828));
    Odrv4 I__9586 (
            .O(N__41828),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__9585 (
            .O(N__41825),
            .I(N__41822));
    InMux I__9584 (
            .O(N__41822),
            .I(N__41819));
    LocalMux I__9583 (
            .O(N__41819),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__9582 (
            .O(N__41816),
            .I(N__41778));
    InMux I__9581 (
            .O(N__41815),
            .I(N__41778));
    InMux I__9580 (
            .O(N__41814),
            .I(N__41778));
    InMux I__9579 (
            .O(N__41813),
            .I(N__41778));
    InMux I__9578 (
            .O(N__41812),
            .I(N__41769));
    InMux I__9577 (
            .O(N__41811),
            .I(N__41769));
    InMux I__9576 (
            .O(N__41810),
            .I(N__41769));
    InMux I__9575 (
            .O(N__41809),
            .I(N__41769));
    InMux I__9574 (
            .O(N__41808),
            .I(N__41764));
    InMux I__9573 (
            .O(N__41807),
            .I(N__41764));
    InMux I__9572 (
            .O(N__41806),
            .I(N__41755));
    InMux I__9571 (
            .O(N__41805),
            .I(N__41755));
    InMux I__9570 (
            .O(N__41804),
            .I(N__41755));
    InMux I__9569 (
            .O(N__41803),
            .I(N__41755));
    InMux I__9568 (
            .O(N__41802),
            .I(N__41746));
    InMux I__9567 (
            .O(N__41801),
            .I(N__41746));
    InMux I__9566 (
            .O(N__41800),
            .I(N__41746));
    InMux I__9565 (
            .O(N__41799),
            .I(N__41746));
    InMux I__9564 (
            .O(N__41798),
            .I(N__41737));
    InMux I__9563 (
            .O(N__41797),
            .I(N__41737));
    InMux I__9562 (
            .O(N__41796),
            .I(N__41737));
    InMux I__9561 (
            .O(N__41795),
            .I(N__41737));
    InMux I__9560 (
            .O(N__41794),
            .I(N__41728));
    InMux I__9559 (
            .O(N__41793),
            .I(N__41728));
    InMux I__9558 (
            .O(N__41792),
            .I(N__41728));
    InMux I__9557 (
            .O(N__41791),
            .I(N__41728));
    InMux I__9556 (
            .O(N__41790),
            .I(N__41719));
    InMux I__9555 (
            .O(N__41789),
            .I(N__41719));
    InMux I__9554 (
            .O(N__41788),
            .I(N__41719));
    InMux I__9553 (
            .O(N__41787),
            .I(N__41719));
    LocalMux I__9552 (
            .O(N__41778),
            .I(N__41714));
    LocalMux I__9551 (
            .O(N__41769),
            .I(N__41714));
    LocalMux I__9550 (
            .O(N__41764),
            .I(N__41711));
    LocalMux I__9549 (
            .O(N__41755),
            .I(N__41704));
    LocalMux I__9548 (
            .O(N__41746),
            .I(N__41704));
    LocalMux I__9547 (
            .O(N__41737),
            .I(N__41704));
    LocalMux I__9546 (
            .O(N__41728),
            .I(N__41699));
    LocalMux I__9545 (
            .O(N__41719),
            .I(N__41699));
    Span4Mux_h I__9544 (
            .O(N__41714),
            .I(N__41696));
    Span4Mux_h I__9543 (
            .O(N__41711),
            .I(N__41693));
    Span4Mux_v I__9542 (
            .O(N__41704),
            .I(N__41686));
    Span4Mux_v I__9541 (
            .O(N__41699),
            .I(N__41686));
    Span4Mux_v I__9540 (
            .O(N__41696),
            .I(N__41686));
    Odrv4 I__9539 (
            .O(N__41693),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__9538 (
            .O(N__41686),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__9537 (
            .O(N__41681),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CascadeMux I__9536 (
            .O(N__41678),
            .I(N__41675));
    InMux I__9535 (
            .O(N__41675),
            .I(N__41672));
    LocalMux I__9534 (
            .O(N__41672),
            .I(N__41668));
    InMux I__9533 (
            .O(N__41671),
            .I(N__41665));
    Span4Mux_h I__9532 (
            .O(N__41668),
            .I(N__41662));
    LocalMux I__9531 (
            .O(N__41665),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv4 I__9530 (
            .O(N__41662),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CEMux I__9529 (
            .O(N__41657),
            .I(N__41652));
    CEMux I__9528 (
            .O(N__41656),
            .I(N__41649));
    CEMux I__9527 (
            .O(N__41655),
            .I(N__41646));
    LocalMux I__9526 (
            .O(N__41652),
            .I(N__41642));
    LocalMux I__9525 (
            .O(N__41649),
            .I(N__41639));
    LocalMux I__9524 (
            .O(N__41646),
            .I(N__41636));
    CEMux I__9523 (
            .O(N__41645),
            .I(N__41633));
    Span4Mux_v I__9522 (
            .O(N__41642),
            .I(N__41630));
    Span4Mux_h I__9521 (
            .O(N__41639),
            .I(N__41627));
    Span4Mux_h I__9520 (
            .O(N__41636),
            .I(N__41624));
    LocalMux I__9519 (
            .O(N__41633),
            .I(N__41621));
    Span4Mux_v I__9518 (
            .O(N__41630),
            .I(N__41618));
    Span4Mux_v I__9517 (
            .O(N__41627),
            .I(N__41615));
    Span4Mux_h I__9516 (
            .O(N__41624),
            .I(N__41612));
    Span4Mux_h I__9515 (
            .O(N__41621),
            .I(N__41609));
    Odrv4 I__9514 (
            .O(N__41618),
            .I(\delay_measurement_inst.delay_tr_timer.N_435_i ));
    Odrv4 I__9513 (
            .O(N__41615),
            .I(\delay_measurement_inst.delay_tr_timer.N_435_i ));
    Odrv4 I__9512 (
            .O(N__41612),
            .I(\delay_measurement_inst.delay_tr_timer.N_435_i ));
    Odrv4 I__9511 (
            .O(N__41609),
            .I(\delay_measurement_inst.delay_tr_timer.N_435_i ));
    CascadeMux I__9510 (
            .O(N__41600),
            .I(N__41597));
    InMux I__9509 (
            .O(N__41597),
            .I(N__41593));
    InMux I__9508 (
            .O(N__41596),
            .I(N__41589));
    LocalMux I__9507 (
            .O(N__41593),
            .I(N__41586));
    InMux I__9506 (
            .O(N__41592),
            .I(N__41582));
    LocalMux I__9505 (
            .O(N__41589),
            .I(N__41577));
    Span4Mux_h I__9504 (
            .O(N__41586),
            .I(N__41577));
    InMux I__9503 (
            .O(N__41585),
            .I(N__41574));
    LocalMux I__9502 (
            .O(N__41582),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    Odrv4 I__9501 (
            .O(N__41577),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    LocalMux I__9500 (
            .O(N__41574),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    InMux I__9499 (
            .O(N__41567),
            .I(N__41563));
    InMux I__9498 (
            .O(N__41566),
            .I(N__41560));
    LocalMux I__9497 (
            .O(N__41563),
            .I(N__41557));
    LocalMux I__9496 (
            .O(N__41560),
            .I(N__41554));
    Span4Mux_h I__9495 (
            .O(N__41557),
            .I(N__41548));
    Span4Mux_h I__9494 (
            .O(N__41554),
            .I(N__41545));
    InMux I__9493 (
            .O(N__41553),
            .I(N__41540));
    InMux I__9492 (
            .O(N__41552),
            .I(N__41540));
    InMux I__9491 (
            .O(N__41551),
            .I(N__41537));
    Odrv4 I__9490 (
            .O(N__41548),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    Odrv4 I__9489 (
            .O(N__41545),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    LocalMux I__9488 (
            .O(N__41540),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    LocalMux I__9487 (
            .O(N__41537),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    CascadeMux I__9486 (
            .O(N__41528),
            .I(N__41524));
    InMux I__9485 (
            .O(N__41527),
            .I(N__41521));
    InMux I__9484 (
            .O(N__41524),
            .I(N__41518));
    LocalMux I__9483 (
            .O(N__41521),
            .I(N__41512));
    LocalMux I__9482 (
            .O(N__41518),
            .I(N__41512));
    InMux I__9481 (
            .O(N__41517),
            .I(N__41508));
    Span4Mux_v I__9480 (
            .O(N__41512),
            .I(N__41505));
    InMux I__9479 (
            .O(N__41511),
            .I(N__41502));
    LocalMux I__9478 (
            .O(N__41508),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    Odrv4 I__9477 (
            .O(N__41505),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    LocalMux I__9476 (
            .O(N__41502),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    CascadeMux I__9475 (
            .O(N__41495),
            .I(N__41492));
    InMux I__9474 (
            .O(N__41492),
            .I(N__41488));
    InMux I__9473 (
            .O(N__41491),
            .I(N__41484));
    LocalMux I__9472 (
            .O(N__41488),
            .I(N__41481));
    InMux I__9471 (
            .O(N__41487),
            .I(N__41478));
    LocalMux I__9470 (
            .O(N__41484),
            .I(N__41473));
    Span4Mux_h I__9469 (
            .O(N__41481),
            .I(N__41473));
    LocalMux I__9468 (
            .O(N__41478),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv4 I__9467 (
            .O(N__41473),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__9466 (
            .O(N__41468),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__9465 (
            .O(N__41465),
            .I(N__41458));
    InMux I__9464 (
            .O(N__41464),
            .I(N__41458));
    InMux I__9463 (
            .O(N__41463),
            .I(N__41455));
    LocalMux I__9462 (
            .O(N__41458),
            .I(N__41452));
    LocalMux I__9461 (
            .O(N__41455),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__9460 (
            .O(N__41452),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__9459 (
            .O(N__41447),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    CascadeMux I__9458 (
            .O(N__41444),
            .I(N__41440));
    CascadeMux I__9457 (
            .O(N__41443),
            .I(N__41437));
    InMux I__9456 (
            .O(N__41440),
            .I(N__41431));
    InMux I__9455 (
            .O(N__41437),
            .I(N__41431));
    InMux I__9454 (
            .O(N__41436),
            .I(N__41428));
    LocalMux I__9453 (
            .O(N__41431),
            .I(N__41425));
    LocalMux I__9452 (
            .O(N__41428),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__9451 (
            .O(N__41425),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__9450 (
            .O(N__41420),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__9449 (
            .O(N__41417),
            .I(N__41413));
    CascadeMux I__9448 (
            .O(N__41416),
            .I(N__41410));
    LocalMux I__9447 (
            .O(N__41413),
            .I(N__41406));
    InMux I__9446 (
            .O(N__41410),
            .I(N__41403));
    InMux I__9445 (
            .O(N__41409),
            .I(N__41400));
    Span4Mux_v I__9444 (
            .O(N__41406),
            .I(N__41395));
    LocalMux I__9443 (
            .O(N__41403),
            .I(N__41395));
    LocalMux I__9442 (
            .O(N__41400),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__9441 (
            .O(N__41395),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__9440 (
            .O(N__41390),
            .I(bfn_18_10_0_));
    CascadeMux I__9439 (
            .O(N__41387),
            .I(N__41384));
    InMux I__9438 (
            .O(N__41384),
            .I(N__41380));
    InMux I__9437 (
            .O(N__41383),
            .I(N__41376));
    LocalMux I__9436 (
            .O(N__41380),
            .I(N__41373));
    InMux I__9435 (
            .O(N__41379),
            .I(N__41370));
    LocalMux I__9434 (
            .O(N__41376),
            .I(N__41365));
    Span4Mux_v I__9433 (
            .O(N__41373),
            .I(N__41365));
    LocalMux I__9432 (
            .O(N__41370),
            .I(N__41362));
    Odrv4 I__9431 (
            .O(N__41365),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__9430 (
            .O(N__41362),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__9429 (
            .O(N__41357),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    CascadeMux I__9428 (
            .O(N__41354),
            .I(N__41350));
    CascadeMux I__9427 (
            .O(N__41353),
            .I(N__41347));
    InMux I__9426 (
            .O(N__41350),
            .I(N__41341));
    InMux I__9425 (
            .O(N__41347),
            .I(N__41341));
    InMux I__9424 (
            .O(N__41346),
            .I(N__41338));
    LocalMux I__9423 (
            .O(N__41341),
            .I(N__41335));
    LocalMux I__9422 (
            .O(N__41338),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv4 I__9421 (
            .O(N__41335),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__9420 (
            .O(N__41330),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__9419 (
            .O(N__41327),
            .I(N__41320));
    InMux I__9418 (
            .O(N__41326),
            .I(N__41320));
    InMux I__9417 (
            .O(N__41325),
            .I(N__41317));
    LocalMux I__9416 (
            .O(N__41320),
            .I(N__41314));
    LocalMux I__9415 (
            .O(N__41317),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__9414 (
            .O(N__41314),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__9413 (
            .O(N__41309),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__9412 (
            .O(N__41306),
            .I(N__41303));
    LocalMux I__9411 (
            .O(N__41303),
            .I(N__41299));
    InMux I__9410 (
            .O(N__41302),
            .I(N__41296));
    Span4Mux_h I__9409 (
            .O(N__41299),
            .I(N__41293));
    LocalMux I__9408 (
            .O(N__41296),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv4 I__9407 (
            .O(N__41293),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__9406 (
            .O(N__41288),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    CascadeMux I__9405 (
            .O(N__41285),
            .I(N__41282));
    InMux I__9404 (
            .O(N__41282),
            .I(N__41278));
    InMux I__9403 (
            .O(N__41281),
            .I(N__41274));
    LocalMux I__9402 (
            .O(N__41278),
            .I(N__41271));
    InMux I__9401 (
            .O(N__41277),
            .I(N__41268));
    LocalMux I__9400 (
            .O(N__41274),
            .I(N__41263));
    Span4Mux_h I__9399 (
            .O(N__41271),
            .I(N__41263));
    LocalMux I__9398 (
            .O(N__41268),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv4 I__9397 (
            .O(N__41263),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__9396 (
            .O(N__41258),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__9395 (
            .O(N__41255),
            .I(N__41248));
    InMux I__9394 (
            .O(N__41254),
            .I(N__41248));
    InMux I__9393 (
            .O(N__41253),
            .I(N__41245));
    LocalMux I__9392 (
            .O(N__41248),
            .I(N__41242));
    LocalMux I__9391 (
            .O(N__41245),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__9390 (
            .O(N__41242),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__9389 (
            .O(N__41237),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    CascadeMux I__9388 (
            .O(N__41234),
            .I(N__41230));
    CascadeMux I__9387 (
            .O(N__41233),
            .I(N__41227));
    InMux I__9386 (
            .O(N__41230),
            .I(N__41221));
    InMux I__9385 (
            .O(N__41227),
            .I(N__41221));
    InMux I__9384 (
            .O(N__41226),
            .I(N__41218));
    LocalMux I__9383 (
            .O(N__41221),
            .I(N__41215));
    LocalMux I__9382 (
            .O(N__41218),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv4 I__9381 (
            .O(N__41215),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__9380 (
            .O(N__41210),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__9379 (
            .O(N__41207),
            .I(N__41203));
    CascadeMux I__9378 (
            .O(N__41206),
            .I(N__41200));
    LocalMux I__9377 (
            .O(N__41203),
            .I(N__41196));
    InMux I__9376 (
            .O(N__41200),
            .I(N__41193));
    InMux I__9375 (
            .O(N__41199),
            .I(N__41190));
    Span4Mux_v I__9374 (
            .O(N__41196),
            .I(N__41185));
    LocalMux I__9373 (
            .O(N__41193),
            .I(N__41185));
    LocalMux I__9372 (
            .O(N__41190),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__9371 (
            .O(N__41185),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__9370 (
            .O(N__41180),
            .I(bfn_18_9_0_));
    CascadeMux I__9369 (
            .O(N__41177),
            .I(N__41174));
    InMux I__9368 (
            .O(N__41174),
            .I(N__41171));
    LocalMux I__9367 (
            .O(N__41171),
            .I(N__41166));
    InMux I__9366 (
            .O(N__41170),
            .I(N__41163));
    InMux I__9365 (
            .O(N__41169),
            .I(N__41160));
    Span4Mux_v I__9364 (
            .O(N__41166),
            .I(N__41157));
    LocalMux I__9363 (
            .O(N__41163),
            .I(N__41154));
    LocalMux I__9362 (
            .O(N__41160),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__9361 (
            .O(N__41157),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__9360 (
            .O(N__41154),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__9359 (
            .O(N__41147),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    CascadeMux I__9358 (
            .O(N__41144),
            .I(N__41140));
    CascadeMux I__9357 (
            .O(N__41143),
            .I(N__41137));
    InMux I__9356 (
            .O(N__41140),
            .I(N__41131));
    InMux I__9355 (
            .O(N__41137),
            .I(N__41131));
    InMux I__9354 (
            .O(N__41136),
            .I(N__41128));
    LocalMux I__9353 (
            .O(N__41131),
            .I(N__41125));
    LocalMux I__9352 (
            .O(N__41128),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv4 I__9351 (
            .O(N__41125),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__9350 (
            .O(N__41120),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__9349 (
            .O(N__41117),
            .I(N__41110));
    InMux I__9348 (
            .O(N__41116),
            .I(N__41110));
    InMux I__9347 (
            .O(N__41115),
            .I(N__41107));
    LocalMux I__9346 (
            .O(N__41110),
            .I(N__41104));
    LocalMux I__9345 (
            .O(N__41107),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv4 I__9344 (
            .O(N__41104),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__9343 (
            .O(N__41099),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    CascadeMux I__9342 (
            .O(N__41096),
            .I(N__41092));
    InMux I__9341 (
            .O(N__41095),
            .I(N__41089));
    InMux I__9340 (
            .O(N__41092),
            .I(N__41085));
    LocalMux I__9339 (
            .O(N__41089),
            .I(N__41082));
    InMux I__9338 (
            .O(N__41088),
            .I(N__41079));
    LocalMux I__9337 (
            .O(N__41085),
            .I(N__41074));
    Span4Mux_h I__9336 (
            .O(N__41082),
            .I(N__41074));
    LocalMux I__9335 (
            .O(N__41079),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv4 I__9334 (
            .O(N__41074),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__9333 (
            .O(N__41069),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    CascadeMux I__9332 (
            .O(N__41066),
            .I(N__41062));
    InMux I__9331 (
            .O(N__41065),
            .I(N__41059));
    InMux I__9330 (
            .O(N__41062),
            .I(N__41055));
    LocalMux I__9329 (
            .O(N__41059),
            .I(N__41052));
    InMux I__9328 (
            .O(N__41058),
            .I(N__41049));
    LocalMux I__9327 (
            .O(N__41055),
            .I(N__41044));
    Span4Mux_h I__9326 (
            .O(N__41052),
            .I(N__41044));
    LocalMux I__9325 (
            .O(N__41049),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv4 I__9324 (
            .O(N__41044),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__9323 (
            .O(N__41039),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    CascadeMux I__9322 (
            .O(N__41036),
            .I(N__41033));
    InMux I__9321 (
            .O(N__41033),
            .I(N__41029));
    InMux I__9320 (
            .O(N__41032),
            .I(N__41025));
    LocalMux I__9319 (
            .O(N__41029),
            .I(N__41022));
    InMux I__9318 (
            .O(N__41028),
            .I(N__41019));
    LocalMux I__9317 (
            .O(N__41025),
            .I(N__41014));
    Span4Mux_h I__9316 (
            .O(N__41022),
            .I(N__41014));
    LocalMux I__9315 (
            .O(N__41019),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv4 I__9314 (
            .O(N__41014),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__9313 (
            .O(N__41009),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__9312 (
            .O(N__41006),
            .I(N__40999));
    InMux I__9311 (
            .O(N__41005),
            .I(N__40999));
    InMux I__9310 (
            .O(N__41004),
            .I(N__40996));
    LocalMux I__9309 (
            .O(N__40999),
            .I(N__40993));
    LocalMux I__9308 (
            .O(N__40996),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__9307 (
            .O(N__40993),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__9306 (
            .O(N__40988),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__9305 (
            .O(N__40985),
            .I(N__40981));
    CascadeMux I__9304 (
            .O(N__40984),
            .I(N__40978));
    InMux I__9303 (
            .O(N__40981),
            .I(N__40972));
    InMux I__9302 (
            .O(N__40978),
            .I(N__40972));
    InMux I__9301 (
            .O(N__40977),
            .I(N__40969));
    LocalMux I__9300 (
            .O(N__40972),
            .I(N__40966));
    LocalMux I__9299 (
            .O(N__40969),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__9298 (
            .O(N__40966),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__9297 (
            .O(N__40961),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__9296 (
            .O(N__40958),
            .I(N__40954));
    CascadeMux I__9295 (
            .O(N__40957),
            .I(N__40951));
    LocalMux I__9294 (
            .O(N__40954),
            .I(N__40947));
    InMux I__9293 (
            .O(N__40951),
            .I(N__40944));
    InMux I__9292 (
            .O(N__40950),
            .I(N__40941));
    Span4Mux_v I__9291 (
            .O(N__40947),
            .I(N__40936));
    LocalMux I__9290 (
            .O(N__40944),
            .I(N__40936));
    LocalMux I__9289 (
            .O(N__40941),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__9288 (
            .O(N__40936),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__9287 (
            .O(N__40931),
            .I(bfn_18_8_0_));
    CascadeMux I__9286 (
            .O(N__40928),
            .I(N__40925));
    InMux I__9285 (
            .O(N__40925),
            .I(N__40921));
    InMux I__9284 (
            .O(N__40924),
            .I(N__40917));
    LocalMux I__9283 (
            .O(N__40921),
            .I(N__40914));
    InMux I__9282 (
            .O(N__40920),
            .I(N__40911));
    LocalMux I__9281 (
            .O(N__40917),
            .I(N__40906));
    Span4Mux_v I__9280 (
            .O(N__40914),
            .I(N__40906));
    LocalMux I__9279 (
            .O(N__40911),
            .I(N__40903));
    Odrv4 I__9278 (
            .O(N__40906),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv4 I__9277 (
            .O(N__40903),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__9276 (
            .O(N__40898),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    CascadeMux I__9275 (
            .O(N__40895),
            .I(N__40891));
    CascadeMux I__9274 (
            .O(N__40894),
            .I(N__40888));
    InMux I__9273 (
            .O(N__40891),
            .I(N__40882));
    InMux I__9272 (
            .O(N__40888),
            .I(N__40882));
    InMux I__9271 (
            .O(N__40887),
            .I(N__40879));
    LocalMux I__9270 (
            .O(N__40882),
            .I(N__40876));
    LocalMux I__9269 (
            .O(N__40879),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__9268 (
            .O(N__40876),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__9267 (
            .O(N__40871),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__9266 (
            .O(N__40868),
            .I(N__40861));
    InMux I__9265 (
            .O(N__40867),
            .I(N__40861));
    InMux I__9264 (
            .O(N__40866),
            .I(N__40858));
    LocalMux I__9263 (
            .O(N__40861),
            .I(N__40855));
    LocalMux I__9262 (
            .O(N__40858),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__9261 (
            .O(N__40855),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__9260 (
            .O(N__40850),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    CascadeMux I__9259 (
            .O(N__40847),
            .I(N__40843));
    InMux I__9258 (
            .O(N__40846),
            .I(N__40840));
    InMux I__9257 (
            .O(N__40843),
            .I(N__40836));
    LocalMux I__9256 (
            .O(N__40840),
            .I(N__40833));
    InMux I__9255 (
            .O(N__40839),
            .I(N__40830));
    LocalMux I__9254 (
            .O(N__40836),
            .I(N__40825));
    Span4Mux_h I__9253 (
            .O(N__40833),
            .I(N__40825));
    LocalMux I__9252 (
            .O(N__40830),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv4 I__9251 (
            .O(N__40825),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__9250 (
            .O(N__40820),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    CascadeMux I__9249 (
            .O(N__40817),
            .I(\phase_controller_inst2.stoper_tr.N_45_cascade_ ));
    InMux I__9248 (
            .O(N__40814),
            .I(N__40810));
    InMux I__9247 (
            .O(N__40813),
            .I(N__40807));
    LocalMux I__9246 (
            .O(N__40810),
            .I(N__40804));
    LocalMux I__9245 (
            .O(N__40807),
            .I(N__40801));
    Span4Mux_h I__9244 (
            .O(N__40804),
            .I(N__40797));
    Span4Mux_v I__9243 (
            .O(N__40801),
            .I(N__40794));
    InMux I__9242 (
            .O(N__40800),
            .I(N__40791));
    Span4Mux_h I__9241 (
            .O(N__40797),
            .I(N__40788));
    Span4Mux_h I__9240 (
            .O(N__40794),
            .I(N__40785));
    LocalMux I__9239 (
            .O(N__40791),
            .I(\phase_controller_inst2.tr_time_passed ));
    Odrv4 I__9238 (
            .O(N__40788),
            .I(\phase_controller_inst2.tr_time_passed ));
    Odrv4 I__9237 (
            .O(N__40785),
            .I(\phase_controller_inst2.tr_time_passed ));
    InMux I__9236 (
            .O(N__40778),
            .I(N__40774));
    InMux I__9235 (
            .O(N__40777),
            .I(N__40771));
    LocalMux I__9234 (
            .O(N__40774),
            .I(N__40766));
    LocalMux I__9233 (
            .O(N__40771),
            .I(N__40766));
    Span4Mux_v I__9232 (
            .O(N__40766),
            .I(N__40762));
    InMux I__9231 (
            .O(N__40765),
            .I(N__40759));
    Odrv4 I__9230 (
            .O(N__40762),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__9229 (
            .O(N__40759),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__9228 (
            .O(N__40754),
            .I(bfn_18_7_0_));
    CascadeMux I__9227 (
            .O(N__40751),
            .I(N__40747));
    InMux I__9226 (
            .O(N__40750),
            .I(N__40744));
    InMux I__9225 (
            .O(N__40747),
            .I(N__40741));
    LocalMux I__9224 (
            .O(N__40744),
            .I(N__40735));
    LocalMux I__9223 (
            .O(N__40741),
            .I(N__40735));
    InMux I__9222 (
            .O(N__40740),
            .I(N__40732));
    Span4Mux_v I__9221 (
            .O(N__40735),
            .I(N__40729));
    LocalMux I__9220 (
            .O(N__40732),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__9219 (
            .O(N__40729),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__9218 (
            .O(N__40724),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    CascadeMux I__9217 (
            .O(N__40721),
            .I(N__40717));
    CascadeMux I__9216 (
            .O(N__40720),
            .I(N__40714));
    InMux I__9215 (
            .O(N__40717),
            .I(N__40708));
    InMux I__9214 (
            .O(N__40714),
            .I(N__40708));
    InMux I__9213 (
            .O(N__40713),
            .I(N__40705));
    LocalMux I__9212 (
            .O(N__40708),
            .I(N__40702));
    LocalMux I__9211 (
            .O(N__40705),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__9210 (
            .O(N__40702),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__9209 (
            .O(N__40697),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__9208 (
            .O(N__40694),
            .I(N__40687));
    InMux I__9207 (
            .O(N__40693),
            .I(N__40687));
    InMux I__9206 (
            .O(N__40692),
            .I(N__40684));
    LocalMux I__9205 (
            .O(N__40687),
            .I(N__40681));
    LocalMux I__9204 (
            .O(N__40684),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__9203 (
            .O(N__40681),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__9202 (
            .O(N__40676),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    CascadeMux I__9201 (
            .O(N__40673),
            .I(N__40670));
    InMux I__9200 (
            .O(N__40670),
            .I(N__40667));
    LocalMux I__9199 (
            .O(N__40667),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__9198 (
            .O(N__40664),
            .I(N__40661));
    LocalMux I__9197 (
            .O(N__40661),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__9196 (
            .O(N__40658),
            .I(N__40655));
    InMux I__9195 (
            .O(N__40655),
            .I(N__40652));
    LocalMux I__9194 (
            .O(N__40652),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__9193 (
            .O(N__40649),
            .I(N__40646));
    LocalMux I__9192 (
            .O(N__40646),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    CascadeMux I__9191 (
            .O(N__40643),
            .I(N__40640));
    InMux I__9190 (
            .O(N__40640),
            .I(N__40637));
    LocalMux I__9189 (
            .O(N__40637),
            .I(N__40634));
    Span4Mux_h I__9188 (
            .O(N__40634),
            .I(N__40631));
    Odrv4 I__9187 (
            .O(N__40631),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__9186 (
            .O(N__40628),
            .I(N__40625));
    LocalMux I__9185 (
            .O(N__40625),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__9184 (
            .O(N__40622),
            .I(N__40603));
    CascadeMux I__9183 (
            .O(N__40621),
            .I(N__40599));
    CascadeMux I__9182 (
            .O(N__40620),
            .I(N__40595));
    CascadeMux I__9181 (
            .O(N__40619),
            .I(N__40591));
    CascadeMux I__9180 (
            .O(N__40618),
            .I(N__40587));
    CascadeMux I__9179 (
            .O(N__40617),
            .I(N__40583));
    CascadeMux I__9178 (
            .O(N__40616),
            .I(N__40579));
    InMux I__9177 (
            .O(N__40615),
            .I(N__40564));
    InMux I__9176 (
            .O(N__40614),
            .I(N__40564));
    InMux I__9175 (
            .O(N__40613),
            .I(N__40564));
    InMux I__9174 (
            .O(N__40612),
            .I(N__40561));
    InMux I__9173 (
            .O(N__40611),
            .I(N__40552));
    InMux I__9172 (
            .O(N__40610),
            .I(N__40552));
    InMux I__9171 (
            .O(N__40609),
            .I(N__40552));
    InMux I__9170 (
            .O(N__40608),
            .I(N__40552));
    CascadeMux I__9169 (
            .O(N__40607),
            .I(N__40548));
    InMux I__9168 (
            .O(N__40606),
            .I(N__40532));
    InMux I__9167 (
            .O(N__40603),
            .I(N__40532));
    InMux I__9166 (
            .O(N__40602),
            .I(N__40532));
    InMux I__9165 (
            .O(N__40599),
            .I(N__40532));
    InMux I__9164 (
            .O(N__40598),
            .I(N__40532));
    InMux I__9163 (
            .O(N__40595),
            .I(N__40532));
    InMux I__9162 (
            .O(N__40594),
            .I(N__40532));
    InMux I__9161 (
            .O(N__40591),
            .I(N__40515));
    InMux I__9160 (
            .O(N__40590),
            .I(N__40515));
    InMux I__9159 (
            .O(N__40587),
            .I(N__40515));
    InMux I__9158 (
            .O(N__40586),
            .I(N__40515));
    InMux I__9157 (
            .O(N__40583),
            .I(N__40515));
    InMux I__9156 (
            .O(N__40582),
            .I(N__40515));
    InMux I__9155 (
            .O(N__40579),
            .I(N__40515));
    InMux I__9154 (
            .O(N__40578),
            .I(N__40515));
    CascadeMux I__9153 (
            .O(N__40577),
            .I(N__40511));
    CascadeMux I__9152 (
            .O(N__40576),
            .I(N__40507));
    CascadeMux I__9151 (
            .O(N__40575),
            .I(N__40503));
    CascadeMux I__9150 (
            .O(N__40574),
            .I(N__40499));
    CascadeMux I__9149 (
            .O(N__40573),
            .I(N__40495));
    CascadeMux I__9148 (
            .O(N__40572),
            .I(N__40491));
    CascadeMux I__9147 (
            .O(N__40571),
            .I(N__40487));
    LocalMux I__9146 (
            .O(N__40564),
            .I(N__40482));
    LocalMux I__9145 (
            .O(N__40561),
            .I(N__40477));
    LocalMux I__9144 (
            .O(N__40552),
            .I(N__40477));
    InMux I__9143 (
            .O(N__40551),
            .I(N__40470));
    InMux I__9142 (
            .O(N__40548),
            .I(N__40470));
    InMux I__9141 (
            .O(N__40547),
            .I(N__40470));
    LocalMux I__9140 (
            .O(N__40532),
            .I(N__40458));
    LocalMux I__9139 (
            .O(N__40515),
            .I(N__40455));
    InMux I__9138 (
            .O(N__40514),
            .I(N__40438));
    InMux I__9137 (
            .O(N__40511),
            .I(N__40438));
    InMux I__9136 (
            .O(N__40510),
            .I(N__40438));
    InMux I__9135 (
            .O(N__40507),
            .I(N__40438));
    InMux I__9134 (
            .O(N__40506),
            .I(N__40438));
    InMux I__9133 (
            .O(N__40503),
            .I(N__40438));
    InMux I__9132 (
            .O(N__40502),
            .I(N__40438));
    InMux I__9131 (
            .O(N__40499),
            .I(N__40438));
    InMux I__9130 (
            .O(N__40498),
            .I(N__40423));
    InMux I__9129 (
            .O(N__40495),
            .I(N__40423));
    InMux I__9128 (
            .O(N__40494),
            .I(N__40423));
    InMux I__9127 (
            .O(N__40491),
            .I(N__40423));
    InMux I__9126 (
            .O(N__40490),
            .I(N__40423));
    InMux I__9125 (
            .O(N__40487),
            .I(N__40423));
    InMux I__9124 (
            .O(N__40486),
            .I(N__40423));
    InMux I__9123 (
            .O(N__40485),
            .I(N__40420));
    Span4Mux_v I__9122 (
            .O(N__40482),
            .I(N__40413));
    Span4Mux_v I__9121 (
            .O(N__40477),
            .I(N__40413));
    LocalMux I__9120 (
            .O(N__40470),
            .I(N__40413));
    InMux I__9119 (
            .O(N__40469),
            .I(N__40410));
    InMux I__9118 (
            .O(N__40468),
            .I(N__40403));
    InMux I__9117 (
            .O(N__40467),
            .I(N__40403));
    InMux I__9116 (
            .O(N__40466),
            .I(N__40403));
    InMux I__9115 (
            .O(N__40465),
            .I(N__40394));
    InMux I__9114 (
            .O(N__40464),
            .I(N__40394));
    InMux I__9113 (
            .O(N__40463),
            .I(N__40394));
    InMux I__9112 (
            .O(N__40462),
            .I(N__40394));
    InMux I__9111 (
            .O(N__40461),
            .I(N__40391));
    Span4Mux_v I__9110 (
            .O(N__40458),
            .I(N__40382));
    Span4Mux_h I__9109 (
            .O(N__40455),
            .I(N__40382));
    LocalMux I__9108 (
            .O(N__40438),
            .I(N__40382));
    LocalMux I__9107 (
            .O(N__40423),
            .I(N__40382));
    LocalMux I__9106 (
            .O(N__40420),
            .I(N__40379));
    Span4Mux_v I__9105 (
            .O(N__40413),
            .I(N__40373));
    LocalMux I__9104 (
            .O(N__40410),
            .I(N__40366));
    LocalMux I__9103 (
            .O(N__40403),
            .I(N__40366));
    LocalMux I__9102 (
            .O(N__40394),
            .I(N__40366));
    LocalMux I__9101 (
            .O(N__40391),
            .I(N__40363));
    Span4Mux_v I__9100 (
            .O(N__40382),
            .I(N__40360));
    Span4Mux_v I__9099 (
            .O(N__40379),
            .I(N__40357));
    InMux I__9098 (
            .O(N__40378),
            .I(N__40354));
    InMux I__9097 (
            .O(N__40377),
            .I(N__40351));
    InMux I__9096 (
            .O(N__40376),
            .I(N__40348));
    Span4Mux_v I__9095 (
            .O(N__40373),
            .I(N__40345));
    Span4Mux_v I__9094 (
            .O(N__40366),
            .I(N__40342));
    Sp12to4 I__9093 (
            .O(N__40363),
            .I(N__40339));
    Span4Mux_v I__9092 (
            .O(N__40360),
            .I(N__40336));
    Sp12to4 I__9091 (
            .O(N__40357),
            .I(N__40333));
    LocalMux I__9090 (
            .O(N__40354),
            .I(N__40326));
    LocalMux I__9089 (
            .O(N__40351),
            .I(N__40326));
    LocalMux I__9088 (
            .O(N__40348),
            .I(N__40326));
    Span4Mux_v I__9087 (
            .O(N__40345),
            .I(N__40323));
    Span4Mux_h I__9086 (
            .O(N__40342),
            .I(N__40320));
    Span12Mux_v I__9085 (
            .O(N__40339),
            .I(N__40313));
    Sp12to4 I__9084 (
            .O(N__40336),
            .I(N__40313));
    Span12Mux_s9_h I__9083 (
            .O(N__40333),
            .I(N__40313));
    IoSpan4Mux I__9082 (
            .O(N__40326),
            .I(N__40310));
    Span4Mux_v I__9081 (
            .O(N__40323),
            .I(N__40307));
    Sp12to4 I__9080 (
            .O(N__40320),
            .I(N__40302));
    Span12Mux_h I__9079 (
            .O(N__40313),
            .I(N__40302));
    Span4Mux_s3_v I__9078 (
            .O(N__40310),
            .I(N__40299));
    Odrv4 I__9077 (
            .O(N__40307),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__9076 (
            .O(N__40302),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__9075 (
            .O(N__40299),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__9074 (
            .O(N__40292),
            .I(N__40289));
    InMux I__9073 (
            .O(N__40289),
            .I(N__40286));
    LocalMux I__9072 (
            .O(N__40286),
            .I(N__40283));
    Odrv4 I__9071 (
            .O(N__40283),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    CascadeMux I__9070 (
            .O(N__40280),
            .I(N__40266));
    CascadeMux I__9069 (
            .O(N__40279),
            .I(N__40262));
    CascadeMux I__9068 (
            .O(N__40278),
            .I(N__40259));
    CascadeMux I__9067 (
            .O(N__40277),
            .I(N__40256));
    CascadeMux I__9066 (
            .O(N__40276),
            .I(N__40252));
    CascadeMux I__9065 (
            .O(N__40275),
            .I(N__40249));
    CascadeMux I__9064 (
            .O(N__40274),
            .I(N__40245));
    CascadeMux I__9063 (
            .O(N__40273),
            .I(N__40242));
    CascadeMux I__9062 (
            .O(N__40272),
            .I(N__40239));
    CascadeMux I__9061 (
            .O(N__40271),
            .I(N__40236));
    CascadeMux I__9060 (
            .O(N__40270),
            .I(N__40233));
    CascadeMux I__9059 (
            .O(N__40269),
            .I(N__40230));
    InMux I__9058 (
            .O(N__40266),
            .I(N__40207));
    InMux I__9057 (
            .O(N__40265),
            .I(N__40207));
    InMux I__9056 (
            .O(N__40262),
            .I(N__40207));
    InMux I__9055 (
            .O(N__40259),
            .I(N__40207));
    InMux I__9054 (
            .O(N__40256),
            .I(N__40207));
    InMux I__9053 (
            .O(N__40255),
            .I(N__40194));
    InMux I__9052 (
            .O(N__40252),
            .I(N__40194));
    InMux I__9051 (
            .O(N__40249),
            .I(N__40194));
    InMux I__9050 (
            .O(N__40248),
            .I(N__40194));
    InMux I__9049 (
            .O(N__40245),
            .I(N__40194));
    InMux I__9048 (
            .O(N__40242),
            .I(N__40194));
    InMux I__9047 (
            .O(N__40239),
            .I(N__40185));
    InMux I__9046 (
            .O(N__40236),
            .I(N__40185));
    InMux I__9045 (
            .O(N__40233),
            .I(N__40185));
    InMux I__9044 (
            .O(N__40230),
            .I(N__40185));
    CascadeMux I__9043 (
            .O(N__40229),
            .I(N__40178));
    CascadeMux I__9042 (
            .O(N__40228),
            .I(N__40175));
    CascadeMux I__9041 (
            .O(N__40227),
            .I(N__40172));
    CascadeMux I__9040 (
            .O(N__40226),
            .I(N__40169));
    CascadeMux I__9039 (
            .O(N__40225),
            .I(N__40165));
    CascadeMux I__9038 (
            .O(N__40224),
            .I(N__40161));
    CascadeMux I__9037 (
            .O(N__40223),
            .I(N__40157));
    CascadeMux I__9036 (
            .O(N__40222),
            .I(N__40153));
    CascadeMux I__9035 (
            .O(N__40221),
            .I(N__40150));
    CascadeMux I__9034 (
            .O(N__40220),
            .I(N__40147));
    CascadeMux I__9033 (
            .O(N__40219),
            .I(N__40144));
    InMux I__9032 (
            .O(N__40218),
            .I(N__40140));
    LocalMux I__9031 (
            .O(N__40207),
            .I(N__40133));
    LocalMux I__9030 (
            .O(N__40194),
            .I(N__40133));
    LocalMux I__9029 (
            .O(N__40185),
            .I(N__40133));
    InMux I__9028 (
            .O(N__40184),
            .I(N__40126));
    InMux I__9027 (
            .O(N__40183),
            .I(N__40126));
    InMux I__9026 (
            .O(N__40182),
            .I(N__40126));
    InMux I__9025 (
            .O(N__40181),
            .I(N__40111));
    InMux I__9024 (
            .O(N__40178),
            .I(N__40102));
    InMux I__9023 (
            .O(N__40175),
            .I(N__40102));
    InMux I__9022 (
            .O(N__40172),
            .I(N__40097));
    InMux I__9021 (
            .O(N__40169),
            .I(N__40097));
    InMux I__9020 (
            .O(N__40168),
            .I(N__40080));
    InMux I__9019 (
            .O(N__40165),
            .I(N__40080));
    InMux I__9018 (
            .O(N__40164),
            .I(N__40080));
    InMux I__9017 (
            .O(N__40161),
            .I(N__40080));
    InMux I__9016 (
            .O(N__40160),
            .I(N__40080));
    InMux I__9015 (
            .O(N__40157),
            .I(N__40080));
    InMux I__9014 (
            .O(N__40156),
            .I(N__40080));
    InMux I__9013 (
            .O(N__40153),
            .I(N__40080));
    InMux I__9012 (
            .O(N__40150),
            .I(N__40071));
    InMux I__9011 (
            .O(N__40147),
            .I(N__40071));
    InMux I__9010 (
            .O(N__40144),
            .I(N__40071));
    InMux I__9009 (
            .O(N__40143),
            .I(N__40071));
    LocalMux I__9008 (
            .O(N__40140),
            .I(N__40064));
    Span4Mux_v I__9007 (
            .O(N__40133),
            .I(N__40064));
    LocalMux I__9006 (
            .O(N__40126),
            .I(N__40064));
    InMux I__9005 (
            .O(N__40125),
            .I(N__40058));
    InMux I__9004 (
            .O(N__40124),
            .I(N__40052));
    InMux I__9003 (
            .O(N__40123),
            .I(N__40052));
    InMux I__9002 (
            .O(N__40122),
            .I(N__40037));
    InMux I__9001 (
            .O(N__40121),
            .I(N__40037));
    InMux I__9000 (
            .O(N__40120),
            .I(N__40037));
    InMux I__8999 (
            .O(N__40119),
            .I(N__40037));
    InMux I__8998 (
            .O(N__40118),
            .I(N__40037));
    InMux I__8997 (
            .O(N__40117),
            .I(N__40037));
    InMux I__8996 (
            .O(N__40116),
            .I(N__40037));
    InMux I__8995 (
            .O(N__40115),
            .I(N__40032));
    InMux I__8994 (
            .O(N__40114),
            .I(N__40032));
    LocalMux I__8993 (
            .O(N__40111),
            .I(N__40029));
    InMux I__8992 (
            .O(N__40110),
            .I(N__40020));
    InMux I__8991 (
            .O(N__40109),
            .I(N__40020));
    InMux I__8990 (
            .O(N__40108),
            .I(N__40020));
    InMux I__8989 (
            .O(N__40107),
            .I(N__40020));
    LocalMux I__8988 (
            .O(N__40102),
            .I(N__40009));
    LocalMux I__8987 (
            .O(N__40097),
            .I(N__40009));
    LocalMux I__8986 (
            .O(N__40080),
            .I(N__40009));
    LocalMux I__8985 (
            .O(N__40071),
            .I(N__40009));
    Span4Mux_h I__8984 (
            .O(N__40064),
            .I(N__40009));
    InMux I__8983 (
            .O(N__40063),
            .I(N__40004));
    InMux I__8982 (
            .O(N__40062),
            .I(N__40004));
    InMux I__8981 (
            .O(N__40061),
            .I(N__40000));
    LocalMux I__8980 (
            .O(N__40058),
            .I(N__39992));
    InMux I__8979 (
            .O(N__40057),
            .I(N__39988));
    LocalMux I__8978 (
            .O(N__40052),
            .I(N__39981));
    LocalMux I__8977 (
            .O(N__40037),
            .I(N__39981));
    LocalMux I__8976 (
            .O(N__40032),
            .I(N__39981));
    Span4Mux_v I__8975 (
            .O(N__40029),
            .I(N__39964));
    LocalMux I__8974 (
            .O(N__40020),
            .I(N__39964));
    Span4Mux_v I__8973 (
            .O(N__40009),
            .I(N__39964));
    LocalMux I__8972 (
            .O(N__40004),
            .I(N__39964));
    InMux I__8971 (
            .O(N__40003),
            .I(N__39954));
    LocalMux I__8970 (
            .O(N__40000),
            .I(N__39951));
    InMux I__8969 (
            .O(N__39999),
            .I(N__39940));
    InMux I__8968 (
            .O(N__39998),
            .I(N__39940));
    InMux I__8967 (
            .O(N__39997),
            .I(N__39940));
    InMux I__8966 (
            .O(N__39996),
            .I(N__39940));
    InMux I__8965 (
            .O(N__39995),
            .I(N__39940));
    Span12Mux_s11_v I__8964 (
            .O(N__39992),
            .I(N__39937));
    InMux I__8963 (
            .O(N__39991),
            .I(N__39934));
    LocalMux I__8962 (
            .O(N__39988),
            .I(N__39929));
    Span4Mux_v I__8961 (
            .O(N__39981),
            .I(N__39929));
    InMux I__8960 (
            .O(N__39980),
            .I(N__39926));
    InMux I__8959 (
            .O(N__39979),
            .I(N__39911));
    InMux I__8958 (
            .O(N__39978),
            .I(N__39911));
    InMux I__8957 (
            .O(N__39977),
            .I(N__39911));
    InMux I__8956 (
            .O(N__39976),
            .I(N__39911));
    InMux I__8955 (
            .O(N__39975),
            .I(N__39911));
    InMux I__8954 (
            .O(N__39974),
            .I(N__39911));
    InMux I__8953 (
            .O(N__39973),
            .I(N__39911));
    Span4Mux_h I__8952 (
            .O(N__39964),
            .I(N__39908));
    InMux I__8951 (
            .O(N__39963),
            .I(N__39893));
    InMux I__8950 (
            .O(N__39962),
            .I(N__39893));
    InMux I__8949 (
            .O(N__39961),
            .I(N__39893));
    InMux I__8948 (
            .O(N__39960),
            .I(N__39893));
    InMux I__8947 (
            .O(N__39959),
            .I(N__39893));
    InMux I__8946 (
            .O(N__39958),
            .I(N__39893));
    InMux I__8945 (
            .O(N__39957),
            .I(N__39893));
    LocalMux I__8944 (
            .O(N__39954),
            .I(N__39886));
    Span12Mux_h I__8943 (
            .O(N__39951),
            .I(N__39886));
    LocalMux I__8942 (
            .O(N__39940),
            .I(N__39886));
    Odrv12 I__8941 (
            .O(N__39937),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__8940 (
            .O(N__39934),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__8939 (
            .O(N__39929),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__8938 (
            .O(N__39926),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__8937 (
            .O(N__39911),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__8936 (
            .O(N__39908),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__8935 (
            .O(N__39893),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__8934 (
            .O(N__39886),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__8933 (
            .O(N__39869),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    CascadeMux I__8932 (
            .O(N__39866),
            .I(N__39861));
    CascadeMux I__8931 (
            .O(N__39865),
            .I(N__39858));
    InMux I__8930 (
            .O(N__39864),
            .I(N__39854));
    InMux I__8929 (
            .O(N__39861),
            .I(N__39851));
    InMux I__8928 (
            .O(N__39858),
            .I(N__39848));
    InMux I__8927 (
            .O(N__39857),
            .I(N__39845));
    LocalMux I__8926 (
            .O(N__39854),
            .I(N__39842));
    LocalMux I__8925 (
            .O(N__39851),
            .I(N__39839));
    LocalMux I__8924 (
            .O(N__39848),
            .I(N__39836));
    LocalMux I__8923 (
            .O(N__39845),
            .I(N__39833));
    Span4Mux_h I__8922 (
            .O(N__39842),
            .I(N__39828));
    Span4Mux_h I__8921 (
            .O(N__39839),
            .I(N__39828));
    Span4Mux_h I__8920 (
            .O(N__39836),
            .I(N__39825));
    Span12Mux_v I__8919 (
            .O(N__39833),
            .I(N__39822));
    Span4Mux_h I__8918 (
            .O(N__39828),
            .I(N__39819));
    Span4Mux_h I__8917 (
            .O(N__39825),
            .I(N__39816));
    Odrv12 I__8916 (
            .O(N__39822),
            .I(\current_shift_inst.N_1310_i ));
    Odrv4 I__8915 (
            .O(N__39819),
            .I(\current_shift_inst.N_1310_i ));
    Odrv4 I__8914 (
            .O(N__39816),
            .I(\current_shift_inst.N_1310_i ));
    InMux I__8913 (
            .O(N__39809),
            .I(N__39806));
    LocalMux I__8912 (
            .O(N__39806),
            .I(N__39803));
    Odrv4 I__8911 (
            .O(N__39803),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__8910 (
            .O(N__39800),
            .I(N__39797));
    InMux I__8909 (
            .O(N__39797),
            .I(N__39794));
    LocalMux I__8908 (
            .O(N__39794),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    InMux I__8907 (
            .O(N__39791),
            .I(N__39788));
    LocalMux I__8906 (
            .O(N__39788),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    CascadeMux I__8905 (
            .O(N__39785),
            .I(N__39782));
    InMux I__8904 (
            .O(N__39782),
            .I(N__39779));
    LocalMux I__8903 (
            .O(N__39779),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__8902 (
            .O(N__39776),
            .I(N__39773));
    LocalMux I__8901 (
            .O(N__39773),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    CascadeMux I__8900 (
            .O(N__39770),
            .I(N__39767));
    InMux I__8899 (
            .O(N__39767),
            .I(N__39764));
    LocalMux I__8898 (
            .O(N__39764),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    InMux I__8897 (
            .O(N__39761),
            .I(N__39758));
    LocalMux I__8896 (
            .O(N__39758),
            .I(N__39755));
    Odrv4 I__8895 (
            .O(N__39755),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    CascadeMux I__8894 (
            .O(N__39752),
            .I(N__39749));
    InMux I__8893 (
            .O(N__39749),
            .I(N__39746));
    LocalMux I__8892 (
            .O(N__39746),
            .I(N__39743));
    Odrv4 I__8891 (
            .O(N__39743),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    CascadeMux I__8890 (
            .O(N__39740),
            .I(N__39737));
    InMux I__8889 (
            .O(N__39737),
            .I(N__39734));
    LocalMux I__8888 (
            .O(N__39734),
            .I(N__39731));
    Odrv4 I__8887 (
            .O(N__39731),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__8886 (
            .O(N__39728),
            .I(N__39725));
    InMux I__8885 (
            .O(N__39725),
            .I(N__39722));
    LocalMux I__8884 (
            .O(N__39722),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__8883 (
            .O(N__39719),
            .I(N__39716));
    LocalMux I__8882 (
            .O(N__39716),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    CascadeMux I__8881 (
            .O(N__39713),
            .I(N__39710));
    InMux I__8880 (
            .O(N__39710),
            .I(N__39707));
    LocalMux I__8879 (
            .O(N__39707),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__8878 (
            .O(N__39704),
            .I(N__39701));
    LocalMux I__8877 (
            .O(N__39701),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    CascadeMux I__8876 (
            .O(N__39698),
            .I(N__39695));
    InMux I__8875 (
            .O(N__39695),
            .I(N__39692));
    LocalMux I__8874 (
            .O(N__39692),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__8873 (
            .O(N__39689),
            .I(N__39686));
    LocalMux I__8872 (
            .O(N__39686),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__8871 (
            .O(N__39683),
            .I(N__39680));
    InMux I__8870 (
            .O(N__39680),
            .I(N__39677));
    LocalMux I__8869 (
            .O(N__39677),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__8868 (
            .O(N__39674),
            .I(N__39671));
    LocalMux I__8867 (
            .O(N__39671),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    InMux I__8866 (
            .O(N__39668),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    SRMux I__8865 (
            .O(N__39665),
            .I(N__39661));
    SRMux I__8864 (
            .O(N__39664),
            .I(N__39658));
    LocalMux I__8863 (
            .O(N__39661),
            .I(N__39652));
    LocalMux I__8862 (
            .O(N__39658),
            .I(N__39652));
    SRMux I__8861 (
            .O(N__39657),
            .I(N__39648));
    Span4Mux_v I__8860 (
            .O(N__39652),
            .I(N__39645));
    SRMux I__8859 (
            .O(N__39651),
            .I(N__39642));
    LocalMux I__8858 (
            .O(N__39648),
            .I(N__39639));
    Span4Mux_h I__8857 (
            .O(N__39645),
            .I(N__39634));
    LocalMux I__8856 (
            .O(N__39642),
            .I(N__39634));
    Span4Mux_h I__8855 (
            .O(N__39639),
            .I(N__39631));
    Span4Mux_h I__8854 (
            .O(N__39634),
            .I(N__39628));
    Odrv4 I__8853 (
            .O(N__39631),
            .I(\phase_controller_inst1.stoper_tr.un1_stoper_state12_1_0_i ));
    Odrv4 I__8852 (
            .O(N__39628),
            .I(\phase_controller_inst1.stoper_tr.un1_stoper_state12_1_0_i ));
    InMux I__8851 (
            .O(N__39623),
            .I(N__39620));
    LocalMux I__8850 (
            .O(N__39620),
            .I(N__39617));
    Span4Mux_h I__8849 (
            .O(N__39617),
            .I(N__39614));
    Odrv4 I__8848 (
            .O(N__39614),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    CascadeMux I__8847 (
            .O(N__39611),
            .I(N__39608));
    InMux I__8846 (
            .O(N__39608),
            .I(N__39605));
    LocalMux I__8845 (
            .O(N__39605),
            .I(N__39602));
    Span4Mux_h I__8844 (
            .O(N__39602),
            .I(N__39599));
    Odrv4 I__8843 (
            .O(N__39599),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    CascadeMux I__8842 (
            .O(N__39596),
            .I(N__39593));
    InMux I__8841 (
            .O(N__39593),
            .I(N__39590));
    LocalMux I__8840 (
            .O(N__39590),
            .I(N__39587));
    Span4Mux_v I__8839 (
            .O(N__39587),
            .I(N__39584));
    Odrv4 I__8838 (
            .O(N__39584),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__8837 (
            .O(N__39581),
            .I(N__39578));
    LocalMux I__8836 (
            .O(N__39578),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__8835 (
            .O(N__39575),
            .I(N__39572));
    InMux I__8834 (
            .O(N__39572),
            .I(N__39569));
    LocalMux I__8833 (
            .O(N__39569),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__8832 (
            .O(N__39566),
            .I(N__39563));
    LocalMux I__8831 (
            .O(N__39563),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__8830 (
            .O(N__39560),
            .I(N__39557));
    InMux I__8829 (
            .O(N__39557),
            .I(N__39554));
    LocalMux I__8828 (
            .O(N__39554),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__8827 (
            .O(N__39551),
            .I(N__39548));
    LocalMux I__8826 (
            .O(N__39548),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    InMux I__8825 (
            .O(N__39545),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__8824 (
            .O(N__39542),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__8823 (
            .O(N__39539),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__8822 (
            .O(N__39536),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__8821 (
            .O(N__39533),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__8820 (
            .O(N__39530),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__8819 (
            .O(N__39527),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__8818 (
            .O(N__39524),
            .I(bfn_17_16_0_));
    InMux I__8817 (
            .O(N__39521),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    CascadeMux I__8816 (
            .O(N__39518),
            .I(N__39515));
    InMux I__8815 (
            .O(N__39515),
            .I(N__39512));
    LocalMux I__8814 (
            .O(N__39512),
            .I(N__39509));
    Span4Mux_h I__8813 (
            .O(N__39509),
            .I(N__39506));
    Odrv4 I__8812 (
            .O(N__39506),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    InMux I__8811 (
            .O(N__39503),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__8810 (
            .O(N__39500),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__8809 (
            .O(N__39497),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__8808 (
            .O(N__39494),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__8807 (
            .O(N__39491),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__8806 (
            .O(N__39488),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__8805 (
            .O(N__39485),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__8804 (
            .O(N__39482),
            .I(bfn_17_15_0_));
    InMux I__8803 (
            .O(N__39479),
            .I(N__39473));
    InMux I__8802 (
            .O(N__39478),
            .I(N__39473));
    LocalMux I__8801 (
            .O(N__39473),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__8800 (
            .O(N__39470),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__8799 (
            .O(N__39467),
            .I(N__39463));
    InMux I__8798 (
            .O(N__39466),
            .I(N__39460));
    LocalMux I__8797 (
            .O(N__39463),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    LocalMux I__8796 (
            .O(N__39460),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__8795 (
            .O(N__39455),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__8794 (
            .O(N__39452),
            .I(N__39448));
    InMux I__8793 (
            .O(N__39451),
            .I(N__39445));
    LocalMux I__8792 (
            .O(N__39448),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    LocalMux I__8791 (
            .O(N__39445),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__8790 (
            .O(N__39440),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__8789 (
            .O(N__39437),
            .I(N__39433));
    InMux I__8788 (
            .O(N__39436),
            .I(N__39428));
    InMux I__8787 (
            .O(N__39433),
            .I(N__39428));
    LocalMux I__8786 (
            .O(N__39428),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__8785 (
            .O(N__39425),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__8784 (
            .O(N__39422),
            .I(N__39416));
    InMux I__8783 (
            .O(N__39421),
            .I(N__39416));
    LocalMux I__8782 (
            .O(N__39416),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__8781 (
            .O(N__39413),
            .I(bfn_17_13_0_));
    InMux I__8780 (
            .O(N__39410),
            .I(N__39407));
    LocalMux I__8779 (
            .O(N__39407),
            .I(N__39403));
    InMux I__8778 (
            .O(N__39406),
            .I(N__39400));
    Odrv4 I__8777 (
            .O(N__39403),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    LocalMux I__8776 (
            .O(N__39400),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__8775 (
            .O(N__39395),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__8774 (
            .O(N__39392),
            .I(N__39389));
    LocalMux I__8773 (
            .O(N__39389),
            .I(N__39385));
    CascadeMux I__8772 (
            .O(N__39388),
            .I(N__39382));
    Span4Mux_h I__8771 (
            .O(N__39385),
            .I(N__39379));
    InMux I__8770 (
            .O(N__39382),
            .I(N__39376));
    Odrv4 I__8769 (
            .O(N__39379),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    LocalMux I__8768 (
            .O(N__39376),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__8767 (
            .O(N__39371),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__8766 (
            .O(N__39368),
            .I(N__39365));
    LocalMux I__8765 (
            .O(N__39365),
            .I(N__39362));
    Span4Mux_h I__8764 (
            .O(N__39362),
            .I(N__39358));
    InMux I__8763 (
            .O(N__39361),
            .I(N__39355));
    Odrv4 I__8762 (
            .O(N__39358),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    LocalMux I__8761 (
            .O(N__39355),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__8760 (
            .O(N__39350),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__8759 (
            .O(N__39347),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__8758 (
            .O(N__39344),
            .I(N__39339));
    InMux I__8757 (
            .O(N__39343),
            .I(N__39334));
    InMux I__8756 (
            .O(N__39342),
            .I(N__39331));
    LocalMux I__8755 (
            .O(N__39339),
            .I(N__39328));
    InMux I__8754 (
            .O(N__39338),
            .I(N__39325));
    InMux I__8753 (
            .O(N__39337),
            .I(N__39322));
    LocalMux I__8752 (
            .O(N__39334),
            .I(N__39319));
    LocalMux I__8751 (
            .O(N__39331),
            .I(N__39316));
    Span4Mux_h I__8750 (
            .O(N__39328),
            .I(N__39313));
    LocalMux I__8749 (
            .O(N__39325),
            .I(N__39308));
    LocalMux I__8748 (
            .O(N__39322),
            .I(N__39308));
    Span4Mux_h I__8747 (
            .O(N__39319),
            .I(N__39303));
    Span4Mux_h I__8746 (
            .O(N__39316),
            .I(N__39303));
    Odrv4 I__8745 (
            .O(N__39313),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv12 I__8744 (
            .O(N__39308),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__8743 (
            .O(N__39303),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    CEMux I__8742 (
            .O(N__39296),
            .I(N__39278));
    CEMux I__8741 (
            .O(N__39295),
            .I(N__39278));
    CEMux I__8740 (
            .O(N__39294),
            .I(N__39278));
    CEMux I__8739 (
            .O(N__39293),
            .I(N__39278));
    CEMux I__8738 (
            .O(N__39292),
            .I(N__39278));
    CEMux I__8737 (
            .O(N__39291),
            .I(N__39278));
    GlobalMux I__8736 (
            .O(N__39278),
            .I(N__39275));
    gio2CtrlBuf I__8735 (
            .O(N__39275),
            .I(\delay_measurement_inst.delay_tr_timer.N_434_i_g ));
    InMux I__8734 (
            .O(N__39272),
            .I(N__39269));
    LocalMux I__8733 (
            .O(N__39269),
            .I(N__39265));
    InMux I__8732 (
            .O(N__39268),
            .I(N__39262));
    Span4Mux_v I__8731 (
            .O(N__39265),
            .I(N__39256));
    LocalMux I__8730 (
            .O(N__39262),
            .I(N__39256));
    InMux I__8729 (
            .O(N__39261),
            .I(N__39253));
    Odrv4 I__8728 (
            .O(N__39256),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    LocalMux I__8727 (
            .O(N__39253),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    InMux I__8726 (
            .O(N__39248),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__8725 (
            .O(N__39245),
            .I(N__39242));
    InMux I__8724 (
            .O(N__39242),
            .I(N__39239));
    LocalMux I__8723 (
            .O(N__39239),
            .I(N__39235));
    CascadeMux I__8722 (
            .O(N__39238),
            .I(N__39231));
    Span4Mux_v I__8721 (
            .O(N__39235),
            .I(N__39228));
    InMux I__8720 (
            .O(N__39234),
            .I(N__39225));
    InMux I__8719 (
            .O(N__39231),
            .I(N__39222));
    Odrv4 I__8718 (
            .O(N__39228),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__8717 (
            .O(N__39225),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__8716 (
            .O(N__39222),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__8715 (
            .O(N__39215),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__8714 (
            .O(N__39212),
            .I(N__39209));
    LocalMux I__8713 (
            .O(N__39209),
            .I(N__39206));
    Span4Mux_v I__8712 (
            .O(N__39206),
            .I(N__39201));
    InMux I__8711 (
            .O(N__39205),
            .I(N__39196));
    InMux I__8710 (
            .O(N__39204),
            .I(N__39196));
    Odrv4 I__8709 (
            .O(N__39201),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    LocalMux I__8708 (
            .O(N__39196),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__8707 (
            .O(N__39191),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__8706 (
            .O(N__39188),
            .I(N__39185));
    LocalMux I__8705 (
            .O(N__39185),
            .I(N__39181));
    CascadeMux I__8704 (
            .O(N__39184),
            .I(N__39178));
    Span4Mux_v I__8703 (
            .O(N__39181),
            .I(N__39174));
    InMux I__8702 (
            .O(N__39178),
            .I(N__39169));
    InMux I__8701 (
            .O(N__39177),
            .I(N__39169));
    Odrv4 I__8700 (
            .O(N__39174),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    LocalMux I__8699 (
            .O(N__39169),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__8698 (
            .O(N__39164),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__8697 (
            .O(N__39161),
            .I(N__39158));
    LocalMux I__8696 (
            .O(N__39158),
            .I(N__39153));
    InMux I__8695 (
            .O(N__39157),
            .I(N__39148));
    InMux I__8694 (
            .O(N__39156),
            .I(N__39148));
    Span4Mux_v I__8693 (
            .O(N__39153),
            .I(N__39145));
    LocalMux I__8692 (
            .O(N__39148),
            .I(N__39142));
    Odrv4 I__8691 (
            .O(N__39145),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__8690 (
            .O(N__39142),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__8689 (
            .O(N__39137),
            .I(bfn_17_12_0_));
    InMux I__8688 (
            .O(N__39134),
            .I(N__39131));
    LocalMux I__8687 (
            .O(N__39131),
            .I(N__39127));
    InMux I__8686 (
            .O(N__39130),
            .I(N__39124));
    Odrv12 I__8685 (
            .O(N__39127),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    LocalMux I__8684 (
            .O(N__39124),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__8683 (
            .O(N__39119),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__8682 (
            .O(N__39116),
            .I(N__39113));
    InMux I__8681 (
            .O(N__39113),
            .I(N__39109));
    InMux I__8680 (
            .O(N__39112),
            .I(N__39106));
    LocalMux I__8679 (
            .O(N__39109),
            .I(N__39103));
    LocalMux I__8678 (
            .O(N__39106),
            .I(N__39100));
    Odrv12 I__8677 (
            .O(N__39103),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    Odrv4 I__8676 (
            .O(N__39100),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__8675 (
            .O(N__39095),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__8674 (
            .O(N__39092),
            .I(N__39088));
    CascadeMux I__8673 (
            .O(N__39091),
            .I(N__39085));
    LocalMux I__8672 (
            .O(N__39088),
            .I(N__39082));
    InMux I__8671 (
            .O(N__39085),
            .I(N__39079));
    Sp12to4 I__8670 (
            .O(N__39082),
            .I(N__39074));
    LocalMux I__8669 (
            .O(N__39079),
            .I(N__39074));
    Odrv12 I__8668 (
            .O(N__39074),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__8667 (
            .O(N__39071),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__8666 (
            .O(N__39068),
            .I(N__39065));
    LocalMux I__8665 (
            .O(N__39065),
            .I(N__39062));
    Span4Mux_v I__8664 (
            .O(N__39062),
            .I(N__39057));
    InMux I__8663 (
            .O(N__39061),
            .I(N__39052));
    InMux I__8662 (
            .O(N__39060),
            .I(N__39052));
    Odrv4 I__8661 (
            .O(N__39057),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    LocalMux I__8660 (
            .O(N__39052),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__8659 (
            .O(N__39047),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__8658 (
            .O(N__39044),
            .I(N__39041));
    InMux I__8657 (
            .O(N__39041),
            .I(N__39038));
    LocalMux I__8656 (
            .O(N__39038),
            .I(N__39034));
    CascadeMux I__8655 (
            .O(N__39037),
            .I(N__39030));
    Span4Mux_h I__8654 (
            .O(N__39034),
            .I(N__39027));
    InMux I__8653 (
            .O(N__39033),
            .I(N__39024));
    InMux I__8652 (
            .O(N__39030),
            .I(N__39021));
    Odrv4 I__8651 (
            .O(N__39027),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    LocalMux I__8650 (
            .O(N__39024),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    LocalMux I__8649 (
            .O(N__39021),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__8648 (
            .O(N__39014),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__8647 (
            .O(N__39011),
            .I(N__39008));
    InMux I__8646 (
            .O(N__39008),
            .I(N__39005));
    LocalMux I__8645 (
            .O(N__39005),
            .I(N__39001));
    CascadeMux I__8644 (
            .O(N__39004),
            .I(N__38996));
    Span4Mux_v I__8643 (
            .O(N__39001),
            .I(N__38993));
    InMux I__8642 (
            .O(N__39000),
            .I(N__38990));
    InMux I__8641 (
            .O(N__38999),
            .I(N__38985));
    InMux I__8640 (
            .O(N__38996),
            .I(N__38985));
    Odrv4 I__8639 (
            .O(N__38993),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    LocalMux I__8638 (
            .O(N__38990),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    LocalMux I__8637 (
            .O(N__38985),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    InMux I__8636 (
            .O(N__38978),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__8635 (
            .O(N__38975),
            .I(N__38972));
    LocalMux I__8634 (
            .O(N__38972),
            .I(N__38969));
    Span4Mux_h I__8633 (
            .O(N__38969),
            .I(N__38965));
    InMux I__8632 (
            .O(N__38968),
            .I(N__38962));
    Odrv4 I__8631 (
            .O(N__38965),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__8630 (
            .O(N__38962),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__8629 (
            .O(N__38957),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__8628 (
            .O(N__38954),
            .I(N__38951));
    LocalMux I__8627 (
            .O(N__38951),
            .I(N__38948));
    Span4Mux_h I__8626 (
            .O(N__38948),
            .I(N__38944));
    InMux I__8625 (
            .O(N__38947),
            .I(N__38941));
    Odrv4 I__8624 (
            .O(N__38944),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    LocalMux I__8623 (
            .O(N__38941),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__8622 (
            .O(N__38936),
            .I(bfn_17_11_0_));
    InMux I__8621 (
            .O(N__38933),
            .I(N__38930));
    LocalMux I__8620 (
            .O(N__38930),
            .I(N__38927));
    Span4Mux_h I__8619 (
            .O(N__38927),
            .I(N__38923));
    InMux I__8618 (
            .O(N__38926),
            .I(N__38920));
    Odrv4 I__8617 (
            .O(N__38923),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    LocalMux I__8616 (
            .O(N__38920),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__8615 (
            .O(N__38915),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__8614 (
            .O(N__38912),
            .I(N__38909));
    LocalMux I__8613 (
            .O(N__38909),
            .I(N__38905));
    CascadeMux I__8612 (
            .O(N__38908),
            .I(N__38902));
    Span4Mux_v I__8611 (
            .O(N__38905),
            .I(N__38899));
    InMux I__8610 (
            .O(N__38902),
            .I(N__38896));
    Odrv4 I__8609 (
            .O(N__38899),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__8608 (
            .O(N__38896),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__8607 (
            .O(N__38891),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__8606 (
            .O(N__38888),
            .I(N__38884));
    CascadeMux I__8605 (
            .O(N__38887),
            .I(N__38881));
    InMux I__8604 (
            .O(N__38884),
            .I(N__38878));
    InMux I__8603 (
            .O(N__38881),
            .I(N__38875));
    LocalMux I__8602 (
            .O(N__38878),
            .I(N__38870));
    LocalMux I__8601 (
            .O(N__38875),
            .I(N__38867));
    InMux I__8600 (
            .O(N__38874),
            .I(N__38862));
    InMux I__8599 (
            .O(N__38873),
            .I(N__38862));
    Odrv4 I__8598 (
            .O(N__38870),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    Odrv4 I__8597 (
            .O(N__38867),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    LocalMux I__8596 (
            .O(N__38862),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    InMux I__8595 (
            .O(N__38855),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__8594 (
            .O(N__38852),
            .I(N__38849));
    LocalMux I__8593 (
            .O(N__38849),
            .I(N__38846));
    Span4Mux_h I__8592 (
            .O(N__38846),
            .I(N__38843));
    Odrv4 I__8591 (
            .O(N__38843),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__8590 (
            .O(N__38840),
            .I(N__38834));
    InMux I__8589 (
            .O(N__38839),
            .I(N__38834));
    LocalMux I__8588 (
            .O(N__38834),
            .I(N__38831));
    Span4Mux_v I__8587 (
            .O(N__38831),
            .I(N__38827));
    InMux I__8586 (
            .O(N__38830),
            .I(N__38824));
    Odrv4 I__8585 (
            .O(N__38827),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__8584 (
            .O(N__38824),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__8583 (
            .O(N__38819),
            .I(N__38815));
    InMux I__8582 (
            .O(N__38818),
            .I(N__38812));
    LocalMux I__8581 (
            .O(N__38815),
            .I(N__38807));
    LocalMux I__8580 (
            .O(N__38812),
            .I(N__38807));
    Odrv4 I__8579 (
            .O(N__38807),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__8578 (
            .O(N__38804),
            .I(N__38801));
    LocalMux I__8577 (
            .O(N__38801),
            .I(N__38797));
    InMux I__8576 (
            .O(N__38800),
            .I(N__38794));
    Span4Mux_v I__8575 (
            .O(N__38797),
            .I(N__38788));
    LocalMux I__8574 (
            .O(N__38794),
            .I(N__38788));
    InMux I__8573 (
            .O(N__38793),
            .I(N__38785));
    Span4Mux_v I__8572 (
            .O(N__38788),
            .I(N__38780));
    LocalMux I__8571 (
            .O(N__38785),
            .I(N__38780));
    Span4Mux_h I__8570 (
            .O(N__38780),
            .I(N__38777));
    Odrv4 I__8569 (
            .O(N__38777),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__8568 (
            .O(N__38774),
            .I(N__38771));
    LocalMux I__8567 (
            .O(N__38771),
            .I(N__38767));
    InMux I__8566 (
            .O(N__38770),
            .I(N__38764));
    Odrv4 I__8565 (
            .O(N__38767),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__8564 (
            .O(N__38764),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__8563 (
            .O(N__38759),
            .I(N__38756));
    LocalMux I__8562 (
            .O(N__38756),
            .I(N__38753));
    Span4Mux_h I__8561 (
            .O(N__38753),
            .I(N__38750));
    Odrv4 I__8560 (
            .O(N__38750),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__8559 (
            .O(N__38747),
            .I(N__38743));
    InMux I__8558 (
            .O(N__38746),
            .I(N__38740));
    LocalMux I__8557 (
            .O(N__38743),
            .I(N__38736));
    LocalMux I__8556 (
            .O(N__38740),
            .I(N__38733));
    InMux I__8555 (
            .O(N__38739),
            .I(N__38730));
    Span4Mux_v I__8554 (
            .O(N__38736),
            .I(N__38727));
    Span4Mux_h I__8553 (
            .O(N__38733),
            .I(N__38722));
    LocalMux I__8552 (
            .O(N__38730),
            .I(N__38722));
    Odrv4 I__8551 (
            .O(N__38727),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__8550 (
            .O(N__38722),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__8549 (
            .O(N__38717),
            .I(N__38714));
    LocalMux I__8548 (
            .O(N__38714),
            .I(N__38711));
    Span4Mux_v I__8547 (
            .O(N__38711),
            .I(N__38707));
    InMux I__8546 (
            .O(N__38710),
            .I(N__38704));
    Odrv4 I__8545 (
            .O(N__38707),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__8544 (
            .O(N__38704),
            .I(\current_shift_inst.un4_control_input1_19 ));
    CascadeMux I__8543 (
            .O(N__38699),
            .I(N__38696));
    InMux I__8542 (
            .O(N__38696),
            .I(N__38693));
    LocalMux I__8541 (
            .O(N__38693),
            .I(N__38690));
    Span4Mux_v I__8540 (
            .O(N__38690),
            .I(N__38687));
    Odrv4 I__8539 (
            .O(N__38687),
            .I(\current_shift_inst.un38_control_input_cry_18_c_RNOZ0 ));
    CascadeMux I__8538 (
            .O(N__38684),
            .I(N__38681));
    InMux I__8537 (
            .O(N__38681),
            .I(N__38678));
    LocalMux I__8536 (
            .O(N__38678),
            .I(N__38675));
    Span4Mux_h I__8535 (
            .O(N__38675),
            .I(N__38672));
    Span4Mux_v I__8534 (
            .O(N__38672),
            .I(N__38668));
    InMux I__8533 (
            .O(N__38671),
            .I(N__38665));
    Odrv4 I__8532 (
            .O(N__38668),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__8531 (
            .O(N__38665),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    CascadeMux I__8530 (
            .O(N__38660),
            .I(N__38657));
    InMux I__8529 (
            .O(N__38657),
            .I(N__38654));
    LocalMux I__8528 (
            .O(N__38654),
            .I(N__38651));
    Span4Mux_v I__8527 (
            .O(N__38651),
            .I(N__38647));
    CascadeMux I__8526 (
            .O(N__38650),
            .I(N__38643));
    Span4Mux_h I__8525 (
            .O(N__38647),
            .I(N__38640));
    InMux I__8524 (
            .O(N__38646),
            .I(N__38637));
    InMux I__8523 (
            .O(N__38643),
            .I(N__38634));
    Odrv4 I__8522 (
            .O(N__38640),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__8521 (
            .O(N__38637),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__8520 (
            .O(N__38634),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__8519 (
            .O(N__38627),
            .I(N__38624));
    LocalMux I__8518 (
            .O(N__38624),
            .I(N__38621));
    Span4Mux_v I__8517 (
            .O(N__38621),
            .I(N__38617));
    InMux I__8516 (
            .O(N__38620),
            .I(N__38614));
    Odrv4 I__8515 (
            .O(N__38617),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__8514 (
            .O(N__38614),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__8513 (
            .O(N__38609),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__8512 (
            .O(N__38606),
            .I(N__38603));
    LocalMux I__8511 (
            .O(N__38603),
            .I(N__38600));
    Span4Mux_h I__8510 (
            .O(N__38600),
            .I(N__38597));
    Span4Mux_v I__8509 (
            .O(N__38597),
            .I(N__38593));
    InMux I__8508 (
            .O(N__38596),
            .I(N__38590));
    Odrv4 I__8507 (
            .O(N__38593),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    LocalMux I__8506 (
            .O(N__38590),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__8505 (
            .O(N__38585),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__8504 (
            .O(N__38582),
            .I(N__38579));
    InMux I__8503 (
            .O(N__38579),
            .I(N__38576));
    LocalMux I__8502 (
            .O(N__38576),
            .I(N__38573));
    Span4Mux_v I__8501 (
            .O(N__38573),
            .I(N__38567));
    InMux I__8500 (
            .O(N__38572),
            .I(N__38562));
    InMux I__8499 (
            .O(N__38571),
            .I(N__38562));
    InMux I__8498 (
            .O(N__38570),
            .I(N__38559));
    Odrv4 I__8497 (
            .O(N__38567),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    LocalMux I__8496 (
            .O(N__38562),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    LocalMux I__8495 (
            .O(N__38559),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    InMux I__8494 (
            .O(N__38552),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__8493 (
            .O(N__38549),
            .I(N__38545));
    InMux I__8492 (
            .O(N__38548),
            .I(N__38542));
    LocalMux I__8491 (
            .O(N__38545),
            .I(N__38537));
    LocalMux I__8490 (
            .O(N__38542),
            .I(N__38537));
    Span4Mux_v I__8489 (
            .O(N__38537),
            .I(N__38533));
    InMux I__8488 (
            .O(N__38536),
            .I(N__38530));
    Odrv4 I__8487 (
            .O(N__38533),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__8486 (
            .O(N__38530),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__8485 (
            .O(N__38525),
            .I(N__38521));
    InMux I__8484 (
            .O(N__38524),
            .I(N__38518));
    LocalMux I__8483 (
            .O(N__38521),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__8482 (
            .O(N__38518),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__8481 (
            .O(N__38513),
            .I(N__38509));
    InMux I__8480 (
            .O(N__38512),
            .I(N__38505));
    LocalMux I__8479 (
            .O(N__38509),
            .I(N__38502));
    InMux I__8478 (
            .O(N__38508),
            .I(N__38499));
    LocalMux I__8477 (
            .O(N__38505),
            .I(N__38492));
    Span4Mux_v I__8476 (
            .O(N__38502),
            .I(N__38492));
    LocalMux I__8475 (
            .O(N__38499),
            .I(N__38492));
    Odrv4 I__8474 (
            .O(N__38492),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__8473 (
            .O(N__38489),
            .I(N__38485));
    InMux I__8472 (
            .O(N__38488),
            .I(N__38482));
    LocalMux I__8471 (
            .O(N__38485),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__8470 (
            .O(N__38482),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__8469 (
            .O(N__38477),
            .I(N__38474));
    LocalMux I__8468 (
            .O(N__38474),
            .I(N__38469));
    InMux I__8467 (
            .O(N__38473),
            .I(N__38464));
    InMux I__8466 (
            .O(N__38472),
            .I(N__38464));
    Odrv12 I__8465 (
            .O(N__38469),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__8464 (
            .O(N__38464),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__8463 (
            .O(N__38459),
            .I(N__38456));
    LocalMux I__8462 (
            .O(N__38456),
            .I(N__38452));
    InMux I__8461 (
            .O(N__38455),
            .I(N__38449));
    Odrv4 I__8460 (
            .O(N__38452),
            .I(\current_shift_inst.un4_control_input1_17 ));
    LocalMux I__8459 (
            .O(N__38449),
            .I(\current_shift_inst.un4_control_input1_17 ));
    InMux I__8458 (
            .O(N__38444),
            .I(N__38441));
    LocalMux I__8457 (
            .O(N__38441),
            .I(N__38438));
    Odrv12 I__8456 (
            .O(N__38438),
            .I(\current_shift_inst.un38_control_input_cry_16_c_RNOZ0 ));
    InMux I__8455 (
            .O(N__38435),
            .I(N__38432));
    LocalMux I__8454 (
            .O(N__38432),
            .I(N__38428));
    InMux I__8453 (
            .O(N__38431),
            .I(N__38425));
    Span4Mux_v I__8452 (
            .O(N__38428),
            .I(N__38422));
    LocalMux I__8451 (
            .O(N__38425),
            .I(N__38419));
    Span4Mux_v I__8450 (
            .O(N__38422),
            .I(N__38415));
    Span4Mux_h I__8449 (
            .O(N__38419),
            .I(N__38412));
    InMux I__8448 (
            .O(N__38418),
            .I(N__38409));
    Odrv4 I__8447 (
            .O(N__38415),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__8446 (
            .O(N__38412),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__8445 (
            .O(N__38409),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__8444 (
            .O(N__38402),
            .I(N__38399));
    LocalMux I__8443 (
            .O(N__38399),
            .I(N__38396));
    Span4Mux_h I__8442 (
            .O(N__38396),
            .I(N__38392));
    InMux I__8441 (
            .O(N__38395),
            .I(N__38389));
    Odrv4 I__8440 (
            .O(N__38392),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__8439 (
            .O(N__38389),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__8438 (
            .O(N__38384),
            .I(N__38380));
    InMux I__8437 (
            .O(N__38383),
            .I(N__38377));
    LocalMux I__8436 (
            .O(N__38380),
            .I(N__38374));
    LocalMux I__8435 (
            .O(N__38377),
            .I(N__38370));
    Span4Mux_h I__8434 (
            .O(N__38374),
            .I(N__38367));
    InMux I__8433 (
            .O(N__38373),
            .I(N__38364));
    Odrv12 I__8432 (
            .O(N__38370),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__8431 (
            .O(N__38367),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__8430 (
            .O(N__38364),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__8429 (
            .O(N__38357),
            .I(N__38354));
    LocalMux I__8428 (
            .O(N__38354),
            .I(N__38350));
    InMux I__8427 (
            .O(N__38353),
            .I(N__38347));
    Odrv4 I__8426 (
            .O(N__38350),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__8425 (
            .O(N__38347),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__8424 (
            .O(N__38342),
            .I(N__38339));
    LocalMux I__8423 (
            .O(N__38339),
            .I(N__38336));
    Span4Mux_h I__8422 (
            .O(N__38336),
            .I(N__38333));
    Span4Mux_h I__8421 (
            .O(N__38333),
            .I(N__38330));
    Odrv4 I__8420 (
            .O(N__38330),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    InMux I__8419 (
            .O(N__38327),
            .I(N__38324));
    LocalMux I__8418 (
            .O(N__38324),
            .I(N__38321));
    Span4Mux_h I__8417 (
            .O(N__38321),
            .I(N__38318));
    Span4Mux_v I__8416 (
            .O(N__38318),
            .I(N__38315));
    Span4Mux_v I__8415 (
            .O(N__38315),
            .I(N__38312));
    Odrv4 I__8414 (
            .O(N__38312),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__8413 (
            .O(N__38309),
            .I(N__38305));
    InMux I__8412 (
            .O(N__38308),
            .I(N__38302));
    LocalMux I__8411 (
            .O(N__38305),
            .I(N__38299));
    LocalMux I__8410 (
            .O(N__38302),
            .I(N__38296));
    Span4Mux_v I__8409 (
            .O(N__38299),
            .I(N__38292));
    Span4Mux_h I__8408 (
            .O(N__38296),
            .I(N__38289));
    InMux I__8407 (
            .O(N__38295),
            .I(N__38286));
    Odrv4 I__8406 (
            .O(N__38292),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__8405 (
            .O(N__38289),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__8404 (
            .O(N__38286),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__8403 (
            .O(N__38279),
            .I(N__38275));
    InMux I__8402 (
            .O(N__38278),
            .I(N__38272));
    LocalMux I__8401 (
            .O(N__38275),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__8400 (
            .O(N__38272),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__8399 (
            .O(N__38267),
            .I(N__38264));
    LocalMux I__8398 (
            .O(N__38264),
            .I(N__38260));
    InMux I__8397 (
            .O(N__38263),
            .I(N__38256));
    Span4Mux_v I__8396 (
            .O(N__38260),
            .I(N__38253));
    InMux I__8395 (
            .O(N__38259),
            .I(N__38250));
    LocalMux I__8394 (
            .O(N__38256),
            .I(N__38247));
    Sp12to4 I__8393 (
            .O(N__38253),
            .I(N__38242));
    LocalMux I__8392 (
            .O(N__38250),
            .I(N__38242));
    Odrv4 I__8391 (
            .O(N__38247),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv12 I__8390 (
            .O(N__38242),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__8389 (
            .O(N__38237),
            .I(N__38233));
    InMux I__8388 (
            .O(N__38236),
            .I(N__38230));
    LocalMux I__8387 (
            .O(N__38233),
            .I(N__38227));
    LocalMux I__8386 (
            .O(N__38230),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__8385 (
            .O(N__38227),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__8384 (
            .O(N__38222),
            .I(N__38219));
    LocalMux I__8383 (
            .O(N__38219),
            .I(N__38216));
    Span4Mux_h I__8382 (
            .O(N__38216),
            .I(N__38213));
    Odrv4 I__8381 (
            .O(N__38213),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__8380 (
            .O(N__38210),
            .I(N__38204));
    InMux I__8379 (
            .O(N__38209),
            .I(N__38204));
    LocalMux I__8378 (
            .O(N__38204),
            .I(N__38200));
    InMux I__8377 (
            .O(N__38203),
            .I(N__38197));
    Span4Mux_h I__8376 (
            .O(N__38200),
            .I(N__38194));
    LocalMux I__8375 (
            .O(N__38197),
            .I(N__38191));
    Span4Mux_v I__8374 (
            .O(N__38194),
            .I(N__38188));
    Span4Mux_v I__8373 (
            .O(N__38191),
            .I(N__38185));
    Odrv4 I__8372 (
            .O(N__38188),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__8371 (
            .O(N__38185),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CEMux I__8370 (
            .O(N__38180),
            .I(N__38162));
    CEMux I__8369 (
            .O(N__38179),
            .I(N__38162));
    CEMux I__8368 (
            .O(N__38178),
            .I(N__38162));
    CEMux I__8367 (
            .O(N__38177),
            .I(N__38162));
    CEMux I__8366 (
            .O(N__38176),
            .I(N__38162));
    CEMux I__8365 (
            .O(N__38175),
            .I(N__38162));
    GlobalMux I__8364 (
            .O(N__38162),
            .I(N__38159));
    gio2CtrlBuf I__8363 (
            .O(N__38159),
            .I(\current_shift_inst.timer_s1.N_166_i_g ));
    InMux I__8362 (
            .O(N__38156),
            .I(N__38150));
    InMux I__8361 (
            .O(N__38155),
            .I(N__38150));
    LocalMux I__8360 (
            .O(N__38150),
            .I(N__38147));
    Span4Mux_v I__8359 (
            .O(N__38147),
            .I(N__38144));
    Span4Mux_h I__8358 (
            .O(N__38144),
            .I(N__38140));
    InMux I__8357 (
            .O(N__38143),
            .I(N__38137));
    Odrv4 I__8356 (
            .O(N__38140),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__8355 (
            .O(N__38137),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__8354 (
            .O(N__38132),
            .I(N__38126));
    InMux I__8353 (
            .O(N__38131),
            .I(N__38126));
    LocalMux I__8352 (
            .O(N__38126),
            .I(\current_shift_inst.un4_control_input1_22 ));
    CascadeMux I__8351 (
            .O(N__38123),
            .I(N__38119));
    InMux I__8350 (
            .O(N__38122),
            .I(N__38115));
    InMux I__8349 (
            .O(N__38119),
            .I(N__38110));
    InMux I__8348 (
            .O(N__38118),
            .I(N__38110));
    LocalMux I__8347 (
            .O(N__38115),
            .I(N__38107));
    LocalMux I__8346 (
            .O(N__38110),
            .I(N__38104));
    Span4Mux_h I__8345 (
            .O(N__38107),
            .I(N__38101));
    Span4Mux_h I__8344 (
            .O(N__38104),
            .I(N__38098));
    Odrv4 I__8343 (
            .O(N__38101),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__8342 (
            .O(N__38098),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__8341 (
            .O(N__38093),
            .I(N__38090));
    LocalMux I__8340 (
            .O(N__38090),
            .I(N__38087));
    Span4Mux_v I__8339 (
            .O(N__38087),
            .I(N__38083));
    InMux I__8338 (
            .O(N__38086),
            .I(N__38080));
    Odrv4 I__8337 (
            .O(N__38083),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__8336 (
            .O(N__38080),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__8335 (
            .O(N__38075),
            .I(N__38069));
    InMux I__8334 (
            .O(N__38074),
            .I(N__38069));
    LocalMux I__8333 (
            .O(N__38069),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__8332 (
            .O(N__38066),
            .I(N__38060));
    InMux I__8331 (
            .O(N__38065),
            .I(N__38060));
    LocalMux I__8330 (
            .O(N__38060),
            .I(N__38057));
    Span4Mux_h I__8329 (
            .O(N__38057),
            .I(N__38053));
    InMux I__8328 (
            .O(N__38056),
            .I(N__38050));
    Odrv4 I__8327 (
            .O(N__38053),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__8326 (
            .O(N__38050),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__8325 (
            .O(N__38045),
            .I(N__38042));
    LocalMux I__8324 (
            .O(N__38042),
            .I(N__38039));
    Span4Mux_h I__8323 (
            .O(N__38039),
            .I(N__38036));
    Odrv4 I__8322 (
            .O(N__38036),
            .I(\current_shift_inst.un38_control_input_cry_17_c_RNOZ0 ));
    InMux I__8321 (
            .O(N__38033),
            .I(N__38030));
    LocalMux I__8320 (
            .O(N__38030),
            .I(N__38026));
    InMux I__8319 (
            .O(N__38029),
            .I(N__38023));
    Span4Mux_v I__8318 (
            .O(N__38026),
            .I(N__38018));
    LocalMux I__8317 (
            .O(N__38023),
            .I(N__38018));
    Span4Mux_h I__8316 (
            .O(N__38018),
            .I(N__38014));
    InMux I__8315 (
            .O(N__38017),
            .I(N__38011));
    Odrv4 I__8314 (
            .O(N__38014),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__8313 (
            .O(N__38011),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__8312 (
            .O(N__38006),
            .I(N__38003));
    LocalMux I__8311 (
            .O(N__38003),
            .I(N__37999));
    InMux I__8310 (
            .O(N__38002),
            .I(N__37996));
    Odrv4 I__8309 (
            .O(N__37999),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__8308 (
            .O(N__37996),
            .I(\current_shift_inst.un4_control_input1_15 ));
    CascadeMux I__8307 (
            .O(N__37991),
            .I(N__37988));
    InMux I__8306 (
            .O(N__37988),
            .I(N__37985));
    LocalMux I__8305 (
            .O(N__37985),
            .I(N__37982));
    Span12Mux_v I__8304 (
            .O(N__37982),
            .I(N__37979));
    Odrv12 I__8303 (
            .O(N__37979),
            .I(\current_shift_inst.un38_control_input_cry_14_c_RNOZ0 ));
    InMux I__8302 (
            .O(N__37976),
            .I(N__37972));
    InMux I__8301 (
            .O(N__37975),
            .I(N__37969));
    LocalMux I__8300 (
            .O(N__37972),
            .I(N__37966));
    LocalMux I__8299 (
            .O(N__37969),
            .I(N__37963));
    Span4Mux_h I__8298 (
            .O(N__37966),
            .I(N__37957));
    Span4Mux_h I__8297 (
            .O(N__37963),
            .I(N__37957));
    InMux I__8296 (
            .O(N__37962),
            .I(N__37954));
    Odrv4 I__8295 (
            .O(N__37957),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    LocalMux I__8294 (
            .O(N__37954),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__8293 (
            .O(N__37949),
            .I(N__37946));
    LocalMux I__8292 (
            .O(N__37946),
            .I(N__37942));
    InMux I__8291 (
            .O(N__37945),
            .I(N__37939));
    Odrv4 I__8290 (
            .O(N__37942),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__8289 (
            .O(N__37939),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__8288 (
            .O(N__37934),
            .I(N__37930));
    InMux I__8287 (
            .O(N__37933),
            .I(N__37927));
    LocalMux I__8286 (
            .O(N__37930),
            .I(N__37924));
    LocalMux I__8285 (
            .O(N__37927),
            .I(N__37921));
    Span4Mux_h I__8284 (
            .O(N__37924),
            .I(N__37917));
    Span4Mux_h I__8283 (
            .O(N__37921),
            .I(N__37914));
    InMux I__8282 (
            .O(N__37920),
            .I(N__37911));
    Odrv4 I__8281 (
            .O(N__37917),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv4 I__8280 (
            .O(N__37914),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__8279 (
            .O(N__37911),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__8278 (
            .O(N__37904),
            .I(N__37900));
    InMux I__8277 (
            .O(N__37903),
            .I(N__37897));
    LocalMux I__8276 (
            .O(N__37900),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__8275 (
            .O(N__37897),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__8274 (
            .O(N__37892),
            .I(N__37888));
    InMux I__8273 (
            .O(N__37891),
            .I(N__37885));
    LocalMux I__8272 (
            .O(N__37888),
            .I(N__37882));
    LocalMux I__8271 (
            .O(N__37885),
            .I(N__37878));
    Span4Mux_v I__8270 (
            .O(N__37882),
            .I(N__37875));
    InMux I__8269 (
            .O(N__37881),
            .I(N__37872));
    Odrv4 I__8268 (
            .O(N__37878),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__8267 (
            .O(N__37875),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__8266 (
            .O(N__37872),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__8265 (
            .O(N__37865),
            .I(N__37861));
    InMux I__8264 (
            .O(N__37864),
            .I(N__37858));
    LocalMux I__8263 (
            .O(N__37861),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__8262 (
            .O(N__37858),
            .I(\current_shift_inst.un4_control_input1_13 ));
    InMux I__8261 (
            .O(N__37853),
            .I(N__37850));
    LocalMux I__8260 (
            .O(N__37850),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__8259 (
            .O(N__37847),
            .I(N__37843));
    InMux I__8258 (
            .O(N__37846),
            .I(N__37840));
    LocalMux I__8257 (
            .O(N__37843),
            .I(\current_shift_inst.un4_control_input1_16 ));
    LocalMux I__8256 (
            .O(N__37840),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__8255 (
            .O(N__37835),
            .I(N__37830));
    InMux I__8254 (
            .O(N__37834),
            .I(N__37825));
    InMux I__8253 (
            .O(N__37833),
            .I(N__37825));
    LocalMux I__8252 (
            .O(N__37830),
            .I(N__37822));
    LocalMux I__8251 (
            .O(N__37825),
            .I(N__37819));
    Span4Mux_v I__8250 (
            .O(N__37822),
            .I(N__37816));
    Span4Mux_h I__8249 (
            .O(N__37819),
            .I(N__37813));
    Odrv4 I__8248 (
            .O(N__37816),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__8247 (
            .O(N__37813),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__8246 (
            .O(N__37808),
            .I(N__37804));
    InMux I__8245 (
            .O(N__37807),
            .I(N__37801));
    LocalMux I__8244 (
            .O(N__37804),
            .I(N__37798));
    LocalMux I__8243 (
            .O(N__37801),
            .I(N__37795));
    Span4Mux_h I__8242 (
            .O(N__37798),
            .I(N__37791));
    Span4Mux_h I__8241 (
            .O(N__37795),
            .I(N__37788));
    InMux I__8240 (
            .O(N__37794),
            .I(N__37785));
    Odrv4 I__8239 (
            .O(N__37791),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__8238 (
            .O(N__37788),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__8237 (
            .O(N__37785),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__8236 (
            .O(N__37778),
            .I(N__37774));
    InMux I__8235 (
            .O(N__37777),
            .I(N__37771));
    LocalMux I__8234 (
            .O(N__37774),
            .I(\current_shift_inst.un4_control_input1_12 ));
    LocalMux I__8233 (
            .O(N__37771),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__8232 (
            .O(N__37766),
            .I(N__37763));
    LocalMux I__8231 (
            .O(N__37763),
            .I(N__37759));
    InMux I__8230 (
            .O(N__37762),
            .I(N__37755));
    Span4Mux_v I__8229 (
            .O(N__37759),
            .I(N__37752));
    InMux I__8228 (
            .O(N__37758),
            .I(N__37749));
    LocalMux I__8227 (
            .O(N__37755),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__8226 (
            .O(N__37752),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__8225 (
            .O(N__37749),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__8224 (
            .O(N__37742),
            .I(N__37738));
    InMux I__8223 (
            .O(N__37741),
            .I(N__37735));
    LocalMux I__8222 (
            .O(N__37738),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__8221 (
            .O(N__37735),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__8220 (
            .O(N__37730),
            .I(N__37727));
    LocalMux I__8219 (
            .O(N__37727),
            .I(N__37717));
    InMux I__8218 (
            .O(N__37726),
            .I(N__37702));
    InMux I__8217 (
            .O(N__37725),
            .I(N__37702));
    InMux I__8216 (
            .O(N__37724),
            .I(N__37702));
    InMux I__8215 (
            .O(N__37723),
            .I(N__37702));
    InMux I__8214 (
            .O(N__37722),
            .I(N__37702));
    InMux I__8213 (
            .O(N__37721),
            .I(N__37702));
    InMux I__8212 (
            .O(N__37720),
            .I(N__37702));
    Span4Mux_h I__8211 (
            .O(N__37717),
            .I(N__37688));
    LocalMux I__8210 (
            .O(N__37702),
            .I(N__37688));
    InMux I__8209 (
            .O(N__37701),
            .I(N__37673));
    InMux I__8208 (
            .O(N__37700),
            .I(N__37673));
    InMux I__8207 (
            .O(N__37699),
            .I(N__37673));
    InMux I__8206 (
            .O(N__37698),
            .I(N__37673));
    InMux I__8205 (
            .O(N__37697),
            .I(N__37673));
    InMux I__8204 (
            .O(N__37696),
            .I(N__37673));
    InMux I__8203 (
            .O(N__37695),
            .I(N__37673));
    InMux I__8202 (
            .O(N__37694),
            .I(N__37668));
    InMux I__8201 (
            .O(N__37693),
            .I(N__37668));
    Odrv4 I__8200 (
            .O(N__37688),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__8199 (
            .O(N__37673),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__8198 (
            .O(N__37668),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__8197 (
            .O(N__37661),
            .I(N__37657));
    InMux I__8196 (
            .O(N__37660),
            .I(N__37654));
    LocalMux I__8195 (
            .O(N__37657),
            .I(N__37651));
    LocalMux I__8194 (
            .O(N__37654),
            .I(N__37647));
    Span4Mux_h I__8193 (
            .O(N__37651),
            .I(N__37644));
    InMux I__8192 (
            .O(N__37650),
            .I(N__37641));
    Odrv4 I__8191 (
            .O(N__37647),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__8190 (
            .O(N__37644),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__8189 (
            .O(N__37641),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__8188 (
            .O(N__37634),
            .I(N__37630));
    InMux I__8187 (
            .O(N__37633),
            .I(N__37627));
    LocalMux I__8186 (
            .O(N__37630),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__8185 (
            .O(N__37627),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__8184 (
            .O(N__37622),
            .I(N__37609));
    InMux I__8183 (
            .O(N__37621),
            .I(N__37609));
    InMux I__8182 (
            .O(N__37620),
            .I(N__37609));
    InMux I__8181 (
            .O(N__37619),
            .I(N__37606));
    InMux I__8180 (
            .O(N__37618),
            .I(N__37599));
    InMux I__8179 (
            .O(N__37617),
            .I(N__37599));
    InMux I__8178 (
            .O(N__37616),
            .I(N__37599));
    LocalMux I__8177 (
            .O(N__37609),
            .I(N__37596));
    LocalMux I__8176 (
            .O(N__37606),
            .I(N__37593));
    LocalMux I__8175 (
            .O(N__37599),
            .I(N__37582));
    Span12Mux_v I__8174 (
            .O(N__37596),
            .I(N__37579));
    Span4Mux_h I__8173 (
            .O(N__37593),
            .I(N__37576));
    InMux I__8172 (
            .O(N__37592),
            .I(N__37573));
    InMux I__8171 (
            .O(N__37591),
            .I(N__37562));
    InMux I__8170 (
            .O(N__37590),
            .I(N__37562));
    InMux I__8169 (
            .O(N__37589),
            .I(N__37562));
    InMux I__8168 (
            .O(N__37588),
            .I(N__37562));
    InMux I__8167 (
            .O(N__37587),
            .I(N__37562));
    InMux I__8166 (
            .O(N__37586),
            .I(N__37557));
    InMux I__8165 (
            .O(N__37585),
            .I(N__37557));
    Odrv4 I__8164 (
            .O(N__37582),
            .I(\phase_controller_inst1.stoper_tr.N_249 ));
    Odrv12 I__8163 (
            .O(N__37579),
            .I(\phase_controller_inst1.stoper_tr.N_249 ));
    Odrv4 I__8162 (
            .O(N__37576),
            .I(\phase_controller_inst1.stoper_tr.N_249 ));
    LocalMux I__8161 (
            .O(N__37573),
            .I(\phase_controller_inst1.stoper_tr.N_249 ));
    LocalMux I__8160 (
            .O(N__37562),
            .I(\phase_controller_inst1.stoper_tr.N_249 ));
    LocalMux I__8159 (
            .O(N__37557),
            .I(\phase_controller_inst1.stoper_tr.N_249 ));
    CascadeMux I__8158 (
            .O(N__37544),
            .I(N__37541));
    InMux I__8157 (
            .O(N__37541),
            .I(N__37536));
    InMux I__8156 (
            .O(N__37540),
            .I(N__37533));
    CascadeMux I__8155 (
            .O(N__37539),
            .I(N__37530));
    LocalMux I__8154 (
            .O(N__37536),
            .I(N__37527));
    LocalMux I__8153 (
            .O(N__37533),
            .I(N__37524));
    InMux I__8152 (
            .O(N__37530),
            .I(N__37520));
    Span4Mux_h I__8151 (
            .O(N__37527),
            .I(N__37517));
    Sp12to4 I__8150 (
            .O(N__37524),
            .I(N__37514));
    InMux I__8149 (
            .O(N__37523),
            .I(N__37511));
    LocalMux I__8148 (
            .O(N__37520),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    Odrv4 I__8147 (
            .O(N__37517),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    Odrv12 I__8146 (
            .O(N__37514),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    LocalMux I__8145 (
            .O(N__37511),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    CascadeMux I__8144 (
            .O(N__37502),
            .I(N__37499));
    InMux I__8143 (
            .O(N__37499),
            .I(N__37494));
    CascadeMux I__8142 (
            .O(N__37498),
            .I(N__37489));
    CascadeMux I__8141 (
            .O(N__37497),
            .I(N__37485));
    LocalMux I__8140 (
            .O(N__37494),
            .I(N__37482));
    InMux I__8139 (
            .O(N__37493),
            .I(N__37479));
    InMux I__8138 (
            .O(N__37492),
            .I(N__37474));
    InMux I__8137 (
            .O(N__37489),
            .I(N__37474));
    InMux I__8136 (
            .O(N__37488),
            .I(N__37469));
    InMux I__8135 (
            .O(N__37485),
            .I(N__37469));
    Span4Mux_v I__8134 (
            .O(N__37482),
            .I(N__37466));
    LocalMux I__8133 (
            .O(N__37479),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2 ));
    LocalMux I__8132 (
            .O(N__37474),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2 ));
    LocalMux I__8131 (
            .O(N__37469),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2 ));
    Odrv4 I__8130 (
            .O(N__37466),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2 ));
    InMux I__8129 (
            .O(N__37457),
            .I(N__37454));
    LocalMux I__8128 (
            .O(N__37454),
            .I(N__37451));
    Span4Mux_v I__8127 (
            .O(N__37451),
            .I(N__37446));
    InMux I__8126 (
            .O(N__37450),
            .I(N__37441));
    InMux I__8125 (
            .O(N__37449),
            .I(N__37441));
    Odrv4 I__8124 (
            .O(N__37446),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    LocalMux I__8123 (
            .O(N__37441),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__8122 (
            .O(N__37436),
            .I(N__37432));
    InMux I__8121 (
            .O(N__37435),
            .I(N__37429));
    LocalMux I__8120 (
            .O(N__37432),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__8119 (
            .O(N__37429),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__8118 (
            .O(N__37424),
            .I(N__37421));
    LocalMux I__8117 (
            .O(N__37421),
            .I(N__37418));
    Span4Mux_h I__8116 (
            .O(N__37418),
            .I(N__37415));
    Odrv4 I__8115 (
            .O(N__37415),
            .I(\current_shift_inst.un38_control_input_cry_11_c_RNOZ0 ));
    InMux I__8114 (
            .O(N__37412),
            .I(N__37408));
    InMux I__8113 (
            .O(N__37411),
            .I(N__37405));
    LocalMux I__8112 (
            .O(N__37408),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__8111 (
            .O(N__37405),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__8110 (
            .O(N__37400),
            .I(N__37396));
    InMux I__8109 (
            .O(N__37399),
            .I(N__37393));
    LocalMux I__8108 (
            .O(N__37396),
            .I(N__37388));
    LocalMux I__8107 (
            .O(N__37393),
            .I(N__37388));
    Span4Mux_h I__8106 (
            .O(N__37388),
            .I(N__37384));
    InMux I__8105 (
            .O(N__37387),
            .I(N__37381));
    Odrv4 I__8104 (
            .O(N__37384),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__8103 (
            .O(N__37381),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__8102 (
            .O(N__37376),
            .I(N__37372));
    InMux I__8101 (
            .O(N__37375),
            .I(N__37369));
    LocalMux I__8100 (
            .O(N__37372),
            .I(N__37364));
    LocalMux I__8099 (
            .O(N__37369),
            .I(N__37364));
    Span4Mux_h I__8098 (
            .O(N__37364),
            .I(N__37360));
    InMux I__8097 (
            .O(N__37363),
            .I(N__37357));
    Odrv4 I__8096 (
            .O(N__37360),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__8095 (
            .O(N__37357),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__8094 (
            .O(N__37352),
            .I(N__37348));
    InMux I__8093 (
            .O(N__37351),
            .I(N__37345));
    LocalMux I__8092 (
            .O(N__37348),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__8091 (
            .O(N__37345),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__8090 (
            .O(N__37340),
            .I(N__37336));
    CascadeMux I__8089 (
            .O(N__37339),
            .I(N__37333));
    LocalMux I__8088 (
            .O(N__37336),
            .I(N__37329));
    InMux I__8087 (
            .O(N__37333),
            .I(N__37324));
    InMux I__8086 (
            .O(N__37332),
            .I(N__37324));
    Span4Mux_h I__8085 (
            .O(N__37329),
            .I(N__37321));
    LocalMux I__8084 (
            .O(N__37324),
            .I(N__37318));
    Odrv4 I__8083 (
            .O(N__37321),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__8082 (
            .O(N__37318),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__8081 (
            .O(N__37313),
            .I(N__37309));
    InMux I__8080 (
            .O(N__37312),
            .I(N__37306));
    LocalMux I__8079 (
            .O(N__37309),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__8078 (
            .O(N__37306),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__8077 (
            .O(N__37301),
            .I(N__37297));
    InMux I__8076 (
            .O(N__37300),
            .I(N__37294));
    LocalMux I__8075 (
            .O(N__37297),
            .I(N__37291));
    LocalMux I__8074 (
            .O(N__37294),
            .I(N__37287));
    Span4Mux_h I__8073 (
            .O(N__37291),
            .I(N__37284));
    InMux I__8072 (
            .O(N__37290),
            .I(N__37281));
    Odrv4 I__8071 (
            .O(N__37287),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__8070 (
            .O(N__37284),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__8069 (
            .O(N__37281),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__8068 (
            .O(N__37274),
            .I(N__37271));
    LocalMux I__8067 (
            .O(N__37271),
            .I(N__37267));
    InMux I__8066 (
            .O(N__37270),
            .I(N__37264));
    Odrv12 I__8065 (
            .O(N__37267),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__8064 (
            .O(N__37264),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__8063 (
            .O(N__37259),
            .I(N__37255));
    InMux I__8062 (
            .O(N__37258),
            .I(N__37252));
    LocalMux I__8061 (
            .O(N__37255),
            .I(N__37249));
    LocalMux I__8060 (
            .O(N__37252),
            .I(N__37246));
    Span4Mux_v I__8059 (
            .O(N__37249),
            .I(N__37240));
    Span4Mux_v I__8058 (
            .O(N__37246),
            .I(N__37240));
    InMux I__8057 (
            .O(N__37245),
            .I(N__37237));
    Odrv4 I__8056 (
            .O(N__37240),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    LocalMux I__8055 (
            .O(N__37237),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__8054 (
            .O(N__37232),
            .I(N__37229));
    LocalMux I__8053 (
            .O(N__37229),
            .I(N__37225));
    InMux I__8052 (
            .O(N__37228),
            .I(N__37222));
    Odrv4 I__8051 (
            .O(N__37225),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__8050 (
            .O(N__37222),
            .I(\current_shift_inst.un4_control_input1_5 ));
    CascadeMux I__8049 (
            .O(N__37217),
            .I(N__37213));
    InMux I__8048 (
            .O(N__37216),
            .I(N__37210));
    InMux I__8047 (
            .O(N__37213),
            .I(N__37207));
    LocalMux I__8046 (
            .O(N__37210),
            .I(N__37204));
    LocalMux I__8045 (
            .O(N__37207),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_1Z0Z_9 ));
    Odrv4 I__8044 (
            .O(N__37204),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_1Z0Z_9 ));
    CascadeMux I__8043 (
            .O(N__37199),
            .I(N__37196));
    InMux I__8042 (
            .O(N__37196),
            .I(N__37192));
    InMux I__8041 (
            .O(N__37195),
            .I(N__37189));
    LocalMux I__8040 (
            .O(N__37192),
            .I(N__37186));
    LocalMux I__8039 (
            .O(N__37189),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9 ));
    Odrv4 I__8038 (
            .O(N__37186),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9 ));
    InMux I__8037 (
            .O(N__37181),
            .I(N__37177));
    CascadeMux I__8036 (
            .O(N__37180),
            .I(N__37174));
    LocalMux I__8035 (
            .O(N__37177),
            .I(N__37171));
    InMux I__8034 (
            .O(N__37174),
            .I(N__37167));
    Span4Mux_h I__8033 (
            .O(N__37171),
            .I(N__37164));
    InMux I__8032 (
            .O(N__37170),
            .I(N__37161));
    LocalMux I__8031 (
            .O(N__37167),
            .I(elapsed_time_ns_1_RNIAE2591_0_2));
    Odrv4 I__8030 (
            .O(N__37164),
            .I(elapsed_time_ns_1_RNIAE2591_0_2));
    LocalMux I__8029 (
            .O(N__37161),
            .I(elapsed_time_ns_1_RNIAE2591_0_2));
    CascadeMux I__8028 (
            .O(N__37154),
            .I(N__37150));
    InMux I__8027 (
            .O(N__37153),
            .I(N__37147));
    InMux I__8026 (
            .O(N__37150),
            .I(N__37143));
    LocalMux I__8025 (
            .O(N__37147),
            .I(N__37140));
    InMux I__8024 (
            .O(N__37146),
            .I(N__37137));
    LocalMux I__8023 (
            .O(N__37143),
            .I(N__37134));
    Odrv4 I__8022 (
            .O(N__37140),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_0_2 ));
    LocalMux I__8021 (
            .O(N__37137),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_0_2 ));
    Odrv4 I__8020 (
            .O(N__37134),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_0_2 ));
    CascadeMux I__8019 (
            .O(N__37127),
            .I(N__37124));
    InMux I__8018 (
            .O(N__37124),
            .I(N__37121));
    LocalMux I__8017 (
            .O(N__37121),
            .I(N__37117));
    CascadeMux I__8016 (
            .O(N__37120),
            .I(N__37114));
    Span4Mux_v I__8015 (
            .O(N__37117),
            .I(N__37109));
    InMux I__8014 (
            .O(N__37114),
            .I(N__37106));
    InMux I__8013 (
            .O(N__37113),
            .I(N__37103));
    InMux I__8012 (
            .O(N__37112),
            .I(N__37100));
    Odrv4 I__8011 (
            .O(N__37109),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2 ));
    LocalMux I__8010 (
            .O(N__37106),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2 ));
    LocalMux I__8009 (
            .O(N__37103),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2 ));
    LocalMux I__8008 (
            .O(N__37100),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2 ));
    InMux I__8007 (
            .O(N__37091),
            .I(N__37088));
    LocalMux I__8006 (
            .O(N__37088),
            .I(N__37083));
    InMux I__8005 (
            .O(N__37087),
            .I(N__37080));
    InMux I__8004 (
            .O(N__37086),
            .I(N__37075));
    Span12Mux_v I__8003 (
            .O(N__37083),
            .I(N__37070));
    LocalMux I__8002 (
            .O(N__37080),
            .I(N__37070));
    InMux I__8001 (
            .O(N__37079),
            .I(N__37067));
    InMux I__8000 (
            .O(N__37078),
            .I(N__37064));
    LocalMux I__7999 (
            .O(N__37075),
            .I(N__37061));
    Span12Mux_s11_h I__7998 (
            .O(N__37070),
            .I(N__37056));
    LocalMux I__7997 (
            .O(N__37067),
            .I(N__37056));
    LocalMux I__7996 (
            .O(N__37064),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    Odrv4 I__7995 (
            .O(N__37061),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    Odrv12 I__7994 (
            .O(N__37056),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    CascadeMux I__7993 (
            .O(N__37049),
            .I(N__37046));
    InMux I__7992 (
            .O(N__37046),
            .I(N__37043));
    LocalMux I__7991 (
            .O(N__37043),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2 ));
    CascadeMux I__7990 (
            .O(N__37040),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2_cascade_ ));
    CascadeMux I__7989 (
            .O(N__37037),
            .I(N__37034));
    InMux I__7988 (
            .O(N__37034),
            .I(N__37030));
    CascadeMux I__7987 (
            .O(N__37033),
            .I(N__37026));
    LocalMux I__7986 (
            .O(N__37030),
            .I(N__37023));
    CascadeMux I__7985 (
            .O(N__37029),
            .I(N__37015));
    InMux I__7984 (
            .O(N__37026),
            .I(N__37012));
    Span4Mux_h I__7983 (
            .O(N__37023),
            .I(N__37009));
    InMux I__7982 (
            .O(N__37022),
            .I(N__37006));
    InMux I__7981 (
            .O(N__37021),
            .I(N__37003));
    InMux I__7980 (
            .O(N__37020),
            .I(N__37000));
    InMux I__7979 (
            .O(N__37019),
            .I(N__36995));
    InMux I__7978 (
            .O(N__37018),
            .I(N__36995));
    InMux I__7977 (
            .O(N__37015),
            .I(N__36992));
    LocalMux I__7976 (
            .O(N__37012),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    Odrv4 I__7975 (
            .O(N__37009),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__7974 (
            .O(N__37006),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__7973 (
            .O(N__37003),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__7972 (
            .O(N__37000),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__7971 (
            .O(N__36995),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__7970 (
            .O(N__36992),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    InMux I__7969 (
            .O(N__36977),
            .I(N__36974));
    LocalMux I__7968 (
            .O(N__36974),
            .I(N__36971));
    Span4Mux_h I__7967 (
            .O(N__36971),
            .I(N__36965));
    InMux I__7966 (
            .O(N__36970),
            .I(N__36962));
    InMux I__7965 (
            .O(N__36969),
            .I(N__36959));
    InMux I__7964 (
            .O(N__36968),
            .I(N__36956));
    Odrv4 I__7963 (
            .O(N__36965),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9 ));
    LocalMux I__7962 (
            .O(N__36962),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9 ));
    LocalMux I__7961 (
            .O(N__36959),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9 ));
    LocalMux I__7960 (
            .O(N__36956),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9 ));
    InMux I__7959 (
            .O(N__36947),
            .I(N__36944));
    LocalMux I__7958 (
            .O(N__36944),
            .I(N__36939));
    InMux I__7957 (
            .O(N__36943),
            .I(N__36936));
    InMux I__7956 (
            .O(N__36942),
            .I(N__36933));
    Odrv4 I__7955 (
            .O(N__36939),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    LocalMux I__7954 (
            .O(N__36936),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    LocalMux I__7953 (
            .O(N__36933),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    InMux I__7952 (
            .O(N__36926),
            .I(N__36923));
    LocalMux I__7951 (
            .O(N__36923),
            .I(N__36919));
    InMux I__7950 (
            .O(N__36922),
            .I(N__36914));
    Span4Mux_v I__7949 (
            .O(N__36919),
            .I(N__36911));
    InMux I__7948 (
            .O(N__36918),
            .I(N__36906));
    InMux I__7947 (
            .O(N__36917),
            .I(N__36906));
    LocalMux I__7946 (
            .O(N__36914),
            .I(elapsed_time_ns_1_RNI1OL2M1_0_9));
    Odrv4 I__7945 (
            .O(N__36911),
            .I(elapsed_time_ns_1_RNI1OL2M1_0_9));
    LocalMux I__7944 (
            .O(N__36906),
            .I(elapsed_time_ns_1_RNI1OL2M1_0_9));
    InMux I__7943 (
            .O(N__36899),
            .I(N__36895));
    InMux I__7942 (
            .O(N__36898),
            .I(N__36892));
    LocalMux I__7941 (
            .O(N__36895),
            .I(\phase_controller_inst1.stoper_tr.N_244 ));
    LocalMux I__7940 (
            .O(N__36892),
            .I(\phase_controller_inst1.stoper_tr.N_244 ));
    InMux I__7939 (
            .O(N__36887),
            .I(N__36884));
    LocalMux I__7938 (
            .O(N__36884),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_0_6 ));
    CascadeMux I__7937 (
            .O(N__36881),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9_cascade_ ));
    CascadeMux I__7936 (
            .O(N__36878),
            .I(\phase_controller_inst1.stoper_tr.N_249_cascade_ ));
    CascadeMux I__7935 (
            .O(N__36875),
            .I(N__36872));
    InMux I__7934 (
            .O(N__36872),
            .I(N__36868));
    InMux I__7933 (
            .O(N__36871),
            .I(N__36864));
    LocalMux I__7932 (
            .O(N__36868),
            .I(N__36861));
    CascadeMux I__7931 (
            .O(N__36867),
            .I(N__36858));
    LocalMux I__7930 (
            .O(N__36864),
            .I(N__36855));
    Span4Mux_h I__7929 (
            .O(N__36861),
            .I(N__36852));
    InMux I__7928 (
            .O(N__36858),
            .I(N__36849));
    Odrv4 I__7927 (
            .O(N__36855),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    Odrv4 I__7926 (
            .O(N__36852),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    LocalMux I__7925 (
            .O(N__36849),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    InMux I__7924 (
            .O(N__36842),
            .I(N__36838));
    InMux I__7923 (
            .O(N__36841),
            .I(N__36833));
    LocalMux I__7922 (
            .O(N__36838),
            .I(N__36830));
    InMux I__7921 (
            .O(N__36837),
            .I(N__36827));
    InMux I__7920 (
            .O(N__36836),
            .I(N__36824));
    LocalMux I__7919 (
            .O(N__36833),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    Odrv4 I__7918 (
            .O(N__36830),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    LocalMux I__7917 (
            .O(N__36827),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    LocalMux I__7916 (
            .O(N__36824),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    InMux I__7915 (
            .O(N__36815),
            .I(N__36810));
    InMux I__7914 (
            .O(N__36814),
            .I(N__36807));
    InMux I__7913 (
            .O(N__36813),
            .I(N__36804));
    LocalMux I__7912 (
            .O(N__36810),
            .I(N__36801));
    LocalMux I__7911 (
            .O(N__36807),
            .I(N__36798));
    LocalMux I__7910 (
            .O(N__36804),
            .I(N__36795));
    Span4Mux_h I__7909 (
            .O(N__36801),
            .I(N__36789));
    Span4Mux_h I__7908 (
            .O(N__36798),
            .I(N__36789));
    Span4Mux_h I__7907 (
            .O(N__36795),
            .I(N__36786));
    InMux I__7906 (
            .O(N__36794),
            .I(N__36783));
    Odrv4 I__7905 (
            .O(N__36789),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6));
    Odrv4 I__7904 (
            .O(N__36786),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6));
    LocalMux I__7903 (
            .O(N__36783),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6));
    InMux I__7902 (
            .O(N__36776),
            .I(N__36771));
    CascadeMux I__7901 (
            .O(N__36775),
            .I(N__36767));
    InMux I__7900 (
            .O(N__36774),
            .I(N__36764));
    LocalMux I__7899 (
            .O(N__36771),
            .I(N__36761));
    InMux I__7898 (
            .O(N__36770),
            .I(N__36758));
    InMux I__7897 (
            .O(N__36767),
            .I(N__36755));
    LocalMux I__7896 (
            .O(N__36764),
            .I(N__36752));
    Span4Mux_h I__7895 (
            .O(N__36761),
            .I(N__36748));
    LocalMux I__7894 (
            .O(N__36758),
            .I(N__36743));
    LocalMux I__7893 (
            .O(N__36755),
            .I(N__36743));
    Span4Mux_h I__7892 (
            .O(N__36752),
            .I(N__36740));
    InMux I__7891 (
            .O(N__36751),
            .I(N__36737));
    Odrv4 I__7890 (
            .O(N__36748),
            .I(\phase_controller_inst1.stoper_tr.N_250 ));
    Odrv12 I__7889 (
            .O(N__36743),
            .I(\phase_controller_inst1.stoper_tr.N_250 ));
    Odrv4 I__7888 (
            .O(N__36740),
            .I(\phase_controller_inst1.stoper_tr.N_250 ));
    LocalMux I__7887 (
            .O(N__36737),
            .I(\phase_controller_inst1.stoper_tr.N_250 ));
    CascadeMux I__7886 (
            .O(N__36728),
            .I(N__36725));
    InMux I__7885 (
            .O(N__36725),
            .I(N__36719));
    InMux I__7884 (
            .O(N__36724),
            .I(N__36719));
    LocalMux I__7883 (
            .O(N__36719),
            .I(N__36716));
    Span4Mux_v I__7882 (
            .O(N__36716),
            .I(N__36711));
    InMux I__7881 (
            .O(N__36715),
            .I(N__36706));
    InMux I__7880 (
            .O(N__36714),
            .I(N__36706));
    Span4Mux_v I__7879 (
            .O(N__36711),
            .I(N__36703));
    LocalMux I__7878 (
            .O(N__36706),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__7877 (
            .O(N__36703),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__7876 (
            .O(N__36698),
            .I(N__36693));
    InMux I__7875 (
            .O(N__36697),
            .I(N__36687));
    InMux I__7874 (
            .O(N__36696),
            .I(N__36687));
    LocalMux I__7873 (
            .O(N__36693),
            .I(N__36684));
    InMux I__7872 (
            .O(N__36692),
            .I(N__36681));
    LocalMux I__7871 (
            .O(N__36687),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__7870 (
            .O(N__36684),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__7869 (
            .O(N__36681),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__7868 (
            .O(N__36674),
            .I(N__36665));
    InMux I__7867 (
            .O(N__36673),
            .I(N__36665));
    InMux I__7866 (
            .O(N__36672),
            .I(N__36665));
    LocalMux I__7865 (
            .O(N__36665),
            .I(N__36662));
    Span4Mux_v I__7864 (
            .O(N__36662),
            .I(N__36659));
    Span4Mux_v I__7863 (
            .O(N__36659),
            .I(N__36656));
    Odrv4 I__7862 (
            .O(N__36656),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    IoInMux I__7861 (
            .O(N__36653),
            .I(N__36650));
    LocalMux I__7860 (
            .O(N__36650),
            .I(N__36647));
    Span4Mux_s0_v I__7859 (
            .O(N__36647),
            .I(N__36644));
    Span4Mux_h I__7858 (
            .O(N__36644),
            .I(N__36641));
    Span4Mux_v I__7857 (
            .O(N__36641),
            .I(N__36638));
    Span4Mux_v I__7856 (
            .O(N__36638),
            .I(N__36635));
    Odrv4 I__7855 (
            .O(N__36635),
            .I(\delay_measurement_inst.delay_tr_timer.N_434_i ));
    CascadeMux I__7854 (
            .O(N__36632),
            .I(N__36627));
    InMux I__7853 (
            .O(N__36631),
            .I(N__36624));
    InMux I__7852 (
            .O(N__36630),
            .I(N__36620));
    InMux I__7851 (
            .O(N__36627),
            .I(N__36617));
    LocalMux I__7850 (
            .O(N__36624),
            .I(N__36614));
    InMux I__7849 (
            .O(N__36623),
            .I(N__36611));
    LocalMux I__7848 (
            .O(N__36620),
            .I(N__36606));
    LocalMux I__7847 (
            .O(N__36617),
            .I(N__36606));
    Span12Mux_h I__7846 (
            .O(N__36614),
            .I(N__36603));
    LocalMux I__7845 (
            .O(N__36611),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv12 I__7844 (
            .O(N__36606),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv12 I__7843 (
            .O(N__36603),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__7842 (
            .O(N__36596),
            .I(N__36593));
    LocalMux I__7841 (
            .O(N__36593),
            .I(N__36590));
    Span4Mux_v I__7840 (
            .O(N__36590),
            .I(N__36585));
    InMux I__7839 (
            .O(N__36589),
            .I(N__36580));
    InMux I__7838 (
            .O(N__36588),
            .I(N__36580));
    Span4Mux_h I__7837 (
            .O(N__36585),
            .I(N__36577));
    LocalMux I__7836 (
            .O(N__36580),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__7835 (
            .O(N__36577),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__7834 (
            .O(N__36572),
            .I(N__36569));
    LocalMux I__7833 (
            .O(N__36569),
            .I(N__36566));
    Span4Mux_h I__7832 (
            .O(N__36566),
            .I(N__36563));
    Span4Mux_h I__7831 (
            .O(N__36563),
            .I(N__36560));
    Span4Mux_v I__7830 (
            .O(N__36560),
            .I(N__36557));
    Odrv4 I__7829 (
            .O(N__36557),
            .I(\phase_controller_inst1.N_55 ));
    CascadeMux I__7828 (
            .O(N__36554),
            .I(N__36550));
    InMux I__7827 (
            .O(N__36553),
            .I(N__36544));
    InMux I__7826 (
            .O(N__36550),
            .I(N__36534));
    InMux I__7825 (
            .O(N__36549),
            .I(N__36534));
    InMux I__7824 (
            .O(N__36548),
            .I(N__36531));
    CascadeMux I__7823 (
            .O(N__36547),
            .I(N__36526));
    LocalMux I__7822 (
            .O(N__36544),
            .I(N__36521));
    CascadeMux I__7821 (
            .O(N__36543),
            .I(N__36503));
    InMux I__7820 (
            .O(N__36542),
            .I(N__36493));
    InMux I__7819 (
            .O(N__36541),
            .I(N__36493));
    InMux I__7818 (
            .O(N__36540),
            .I(N__36493));
    InMux I__7817 (
            .O(N__36539),
            .I(N__36493));
    LocalMux I__7816 (
            .O(N__36534),
            .I(N__36488));
    LocalMux I__7815 (
            .O(N__36531),
            .I(N__36488));
    InMux I__7814 (
            .O(N__36530),
            .I(N__36485));
    InMux I__7813 (
            .O(N__36529),
            .I(N__36480));
    InMux I__7812 (
            .O(N__36526),
            .I(N__36480));
    InMux I__7811 (
            .O(N__36525),
            .I(N__36477));
    InMux I__7810 (
            .O(N__36524),
            .I(N__36474));
    Span4Mux_v I__7809 (
            .O(N__36521),
            .I(N__36471));
    InMux I__7808 (
            .O(N__36520),
            .I(N__36466));
    InMux I__7807 (
            .O(N__36519),
            .I(N__36466));
    InMux I__7806 (
            .O(N__36518),
            .I(N__36459));
    InMux I__7805 (
            .O(N__36517),
            .I(N__36459));
    InMux I__7804 (
            .O(N__36516),
            .I(N__36459));
    InMux I__7803 (
            .O(N__36515),
            .I(N__36454));
    InMux I__7802 (
            .O(N__36514),
            .I(N__36454));
    InMux I__7801 (
            .O(N__36513),
            .I(N__36443));
    InMux I__7800 (
            .O(N__36512),
            .I(N__36443));
    InMux I__7799 (
            .O(N__36511),
            .I(N__36443));
    InMux I__7798 (
            .O(N__36510),
            .I(N__36443));
    InMux I__7797 (
            .O(N__36509),
            .I(N__36443));
    InMux I__7796 (
            .O(N__36508),
            .I(N__36434));
    InMux I__7795 (
            .O(N__36507),
            .I(N__36434));
    InMux I__7794 (
            .O(N__36506),
            .I(N__36434));
    InMux I__7793 (
            .O(N__36503),
            .I(N__36434));
    InMux I__7792 (
            .O(N__36502),
            .I(N__36431));
    LocalMux I__7791 (
            .O(N__36493),
            .I(N__36426));
    Span4Mux_h I__7790 (
            .O(N__36488),
            .I(N__36426));
    LocalMux I__7789 (
            .O(N__36485),
            .I(N__36421));
    LocalMux I__7788 (
            .O(N__36480),
            .I(N__36421));
    LocalMux I__7787 (
            .O(N__36477),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__7786 (
            .O(N__36474),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__7785 (
            .O(N__36471),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__7784 (
            .O(N__36466),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__7783 (
            .O(N__36459),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__7782 (
            .O(N__36454),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__7781 (
            .O(N__36443),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__7780 (
            .O(N__36434),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__7779 (
            .O(N__36431),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__7778 (
            .O(N__36426),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__7777 (
            .O(N__36421),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    CascadeMux I__7776 (
            .O(N__36398),
            .I(N__36393));
    CascadeMux I__7775 (
            .O(N__36397),
            .I(N__36390));
    CascadeMux I__7774 (
            .O(N__36396),
            .I(N__36386));
    InMux I__7773 (
            .O(N__36393),
            .I(N__36378));
    InMux I__7772 (
            .O(N__36390),
            .I(N__36378));
    InMux I__7771 (
            .O(N__36389),
            .I(N__36378));
    InMux I__7770 (
            .O(N__36386),
            .I(N__36371));
    InMux I__7769 (
            .O(N__36385),
            .I(N__36371));
    LocalMux I__7768 (
            .O(N__36378),
            .I(N__36367));
    InMux I__7767 (
            .O(N__36377),
            .I(N__36364));
    CascadeMux I__7766 (
            .O(N__36376),
            .I(N__36359));
    LocalMux I__7765 (
            .O(N__36371),
            .I(N__36356));
    InMux I__7764 (
            .O(N__36370),
            .I(N__36353));
    Span4Mux_v I__7763 (
            .O(N__36367),
            .I(N__36348));
    LocalMux I__7762 (
            .O(N__36364),
            .I(N__36348));
    InMux I__7761 (
            .O(N__36363),
            .I(N__36343));
    InMux I__7760 (
            .O(N__36362),
            .I(N__36343));
    InMux I__7759 (
            .O(N__36359),
            .I(N__36340));
    Odrv4 I__7758 (
            .O(N__36356),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    LocalMux I__7757 (
            .O(N__36353),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    Odrv4 I__7756 (
            .O(N__36348),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    LocalMux I__7755 (
            .O(N__36343),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    LocalMux I__7754 (
            .O(N__36340),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    CascadeMux I__7753 (
            .O(N__36329),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_ ));
    InMux I__7752 (
            .O(N__36326),
            .I(N__36323));
    LocalMux I__7751 (
            .O(N__36323),
            .I(N__36318));
    InMux I__7750 (
            .O(N__36322),
            .I(N__36315));
    CascadeMux I__7749 (
            .O(N__36321),
            .I(N__36311));
    Span4Mux_v I__7748 (
            .O(N__36318),
            .I(N__36304));
    LocalMux I__7747 (
            .O(N__36315),
            .I(N__36301));
    InMux I__7746 (
            .O(N__36314),
            .I(N__36298));
    InMux I__7745 (
            .O(N__36311),
            .I(N__36293));
    InMux I__7744 (
            .O(N__36310),
            .I(N__36293));
    InMux I__7743 (
            .O(N__36309),
            .I(N__36288));
    InMux I__7742 (
            .O(N__36308),
            .I(N__36288));
    InMux I__7741 (
            .O(N__36307),
            .I(N__36285));
    Span4Mux_h I__7740 (
            .O(N__36304),
            .I(N__36282));
    Odrv4 I__7739 (
            .O(N__36301),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    LocalMux I__7738 (
            .O(N__36298),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    LocalMux I__7737 (
            .O(N__36293),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    LocalMux I__7736 (
            .O(N__36288),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    LocalMux I__7735 (
            .O(N__36285),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    Odrv4 I__7734 (
            .O(N__36282),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    CascadeMux I__7733 (
            .O(N__36269),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_));
    InMux I__7732 (
            .O(N__36266),
            .I(N__36261));
    InMux I__7731 (
            .O(N__36265),
            .I(N__36256));
    InMux I__7730 (
            .O(N__36264),
            .I(N__36256));
    LocalMux I__7729 (
            .O(N__36261),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ));
    LocalMux I__7728 (
            .O(N__36256),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ));
    InMux I__7727 (
            .O(N__36251),
            .I(N__36244));
    InMux I__7726 (
            .O(N__36250),
            .I(N__36244));
    InMux I__7725 (
            .O(N__36249),
            .I(N__36241));
    LocalMux I__7724 (
            .O(N__36244),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ));
    LocalMux I__7723 (
            .O(N__36241),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ));
    InMux I__7722 (
            .O(N__36236),
            .I(N__36233));
    LocalMux I__7721 (
            .O(N__36233),
            .I(N__36229));
    InMux I__7720 (
            .O(N__36232),
            .I(N__36226));
    Odrv4 I__7719 (
            .O(N__36229),
            .I(elapsed_time_ns_1_RNI0GIF91_0_26));
    LocalMux I__7718 (
            .O(N__36226),
            .I(elapsed_time_ns_1_RNI0GIF91_0_26));
    InMux I__7717 (
            .O(N__36221),
            .I(N__36218));
    LocalMux I__7716 (
            .O(N__36218),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6 ));
    CascadeMux I__7715 (
            .O(N__36215),
            .I(N__36212));
    InMux I__7714 (
            .O(N__36212),
            .I(N__36209));
    LocalMux I__7713 (
            .O(N__36209),
            .I(elapsed_time_ns_1_RNITCIF91_0_23));
    CascadeMux I__7712 (
            .O(N__36206),
            .I(elapsed_time_ns_1_RNITCIF91_0_23_cascade_));
    InMux I__7711 (
            .O(N__36203),
            .I(N__36200));
    LocalMux I__7710 (
            .O(N__36200),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_0_15 ));
    CascadeMux I__7709 (
            .O(N__36197),
            .I(N__36194));
    InMux I__7708 (
            .O(N__36194),
            .I(N__36190));
    InMux I__7707 (
            .O(N__36193),
            .I(N__36187));
    LocalMux I__7706 (
            .O(N__36190),
            .I(elapsed_time_ns_1_RNI1HIF91_0_27));
    LocalMux I__7705 (
            .O(N__36187),
            .I(elapsed_time_ns_1_RNI1HIF91_0_27));
    InMux I__7704 (
            .O(N__36182),
            .I(N__36179));
    LocalMux I__7703 (
            .O(N__36179),
            .I(N__36173));
    CascadeMux I__7702 (
            .O(N__36178),
            .I(N__36168));
    CascadeMux I__7701 (
            .O(N__36177),
            .I(N__36164));
    CascadeMux I__7700 (
            .O(N__36176),
            .I(N__36160));
    Span4Mux_h I__7699 (
            .O(N__36173),
            .I(N__36157));
    CascadeMux I__7698 (
            .O(N__36172),
            .I(N__36149));
    CascadeMux I__7697 (
            .O(N__36171),
            .I(N__36146));
    InMux I__7696 (
            .O(N__36168),
            .I(N__36141));
    InMux I__7695 (
            .O(N__36167),
            .I(N__36138));
    InMux I__7694 (
            .O(N__36164),
            .I(N__36135));
    InMux I__7693 (
            .O(N__36163),
            .I(N__36130));
    InMux I__7692 (
            .O(N__36160),
            .I(N__36130));
    Span4Mux_v I__7691 (
            .O(N__36157),
            .I(N__36121));
    InMux I__7690 (
            .O(N__36156),
            .I(N__36114));
    InMux I__7689 (
            .O(N__36155),
            .I(N__36114));
    InMux I__7688 (
            .O(N__36154),
            .I(N__36114));
    InMux I__7687 (
            .O(N__36153),
            .I(N__36107));
    InMux I__7686 (
            .O(N__36152),
            .I(N__36107));
    InMux I__7685 (
            .O(N__36149),
            .I(N__36107));
    InMux I__7684 (
            .O(N__36146),
            .I(N__36100));
    InMux I__7683 (
            .O(N__36145),
            .I(N__36100));
    InMux I__7682 (
            .O(N__36144),
            .I(N__36100));
    LocalMux I__7681 (
            .O(N__36141),
            .I(N__36091));
    LocalMux I__7680 (
            .O(N__36138),
            .I(N__36091));
    LocalMux I__7679 (
            .O(N__36135),
            .I(N__36091));
    LocalMux I__7678 (
            .O(N__36130),
            .I(N__36091));
    InMux I__7677 (
            .O(N__36129),
            .I(N__36088));
    InMux I__7676 (
            .O(N__36128),
            .I(N__36081));
    InMux I__7675 (
            .O(N__36127),
            .I(N__36081));
    InMux I__7674 (
            .O(N__36126),
            .I(N__36081));
    InMux I__7673 (
            .O(N__36125),
            .I(N__36076));
    InMux I__7672 (
            .O(N__36124),
            .I(N__36076));
    Odrv4 I__7671 (
            .O(N__36121),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__7670 (
            .O(N__36114),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__7669 (
            .O(N__36107),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__7668 (
            .O(N__36100),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    Odrv4 I__7667 (
            .O(N__36091),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__7666 (
            .O(N__36088),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__7665 (
            .O(N__36081),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__7664 (
            .O(N__36076),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    CascadeMux I__7663 (
            .O(N__36059),
            .I(N__36056));
    InMux I__7662 (
            .O(N__36056),
            .I(N__36052));
    InMux I__7661 (
            .O(N__36055),
            .I(N__36049));
    LocalMux I__7660 (
            .O(N__36052),
            .I(elapsed_time_ns_1_RNIUDIF91_0_24));
    LocalMux I__7659 (
            .O(N__36049),
            .I(elapsed_time_ns_1_RNIUDIF91_0_24));
    CascadeMux I__7658 (
            .O(N__36044),
            .I(\delay_measurement_inst.delay_tr_timer.N_367_cascade_ ));
    InMux I__7657 (
            .O(N__36041),
            .I(N__36037));
    InMux I__7656 (
            .O(N__36040),
            .I(N__36033));
    LocalMux I__7655 (
            .O(N__36037),
            .I(N__36030));
    InMux I__7654 (
            .O(N__36036),
            .I(N__36027));
    LocalMux I__7653 (
            .O(N__36033),
            .I(N__36020));
    Span4Mux_h I__7652 (
            .O(N__36030),
            .I(N__36020));
    LocalMux I__7651 (
            .O(N__36027),
            .I(N__36020));
    Odrv4 I__7650 (
            .O(N__36020),
            .I(\delay_measurement_inst.delay_tr_timer.N_378 ));
    InMux I__7649 (
            .O(N__36017),
            .I(N__36014));
    LocalMux I__7648 (
            .O(N__36014),
            .I(N__36011));
    Span12Mux_v I__7647 (
            .O(N__36011),
            .I(N__36006));
    InMux I__7646 (
            .O(N__36010),
            .I(N__36001));
    InMux I__7645 (
            .O(N__36009),
            .I(N__36001));
    Odrv12 I__7644 (
            .O(N__36006),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__7643 (
            .O(N__36001),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__7642 (
            .O(N__35996),
            .I(N__35993));
    LocalMux I__7641 (
            .O(N__35993),
            .I(\delay_measurement_inst.delay_tr_timer.N_349 ));
    InMux I__7640 (
            .O(N__35990),
            .I(N__35987));
    LocalMux I__7639 (
            .O(N__35987),
            .I(elapsed_time_ns_1_RNIVEIF91_0_25));
    CascadeMux I__7638 (
            .O(N__35984),
            .I(elapsed_time_ns_1_RNIVEIF91_0_25_cascade_));
    InMux I__7637 (
            .O(N__35981),
            .I(N__35978));
    LocalMux I__7636 (
            .O(N__35978),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_o5_6Z0Z_15 ));
    CascadeMux I__7635 (
            .O(N__35975),
            .I(N__35972));
    InMux I__7634 (
            .O(N__35972),
            .I(N__35968));
    InMux I__7633 (
            .O(N__35971),
            .I(N__35965));
    LocalMux I__7632 (
            .O(N__35968),
            .I(elapsed_time_ns_1_RNI2IIF91_0_28));
    LocalMux I__7631 (
            .O(N__35965),
            .I(elapsed_time_ns_1_RNI2IIF91_0_28));
    CascadeMux I__7630 (
            .O(N__35960),
            .I(N__35957));
    InMux I__7629 (
            .O(N__35957),
            .I(N__35954));
    LocalMux I__7628 (
            .O(N__35954),
            .I(N__35951));
    Span4Mux_v I__7627 (
            .O(N__35951),
            .I(N__35947));
    InMux I__7626 (
            .O(N__35950),
            .I(N__35944));
    Odrv4 I__7625 (
            .O(N__35947),
            .I(\delay_measurement_inst.delay_tr_timer.N_345 ));
    LocalMux I__7624 (
            .O(N__35944),
            .I(\delay_measurement_inst.delay_tr_timer.N_345 ));
    InMux I__7623 (
            .O(N__35939),
            .I(N__35936));
    LocalMux I__7622 (
            .O(N__35936),
            .I(\delay_measurement_inst.delay_tr_timer.N_348 ));
    InMux I__7621 (
            .O(N__35933),
            .I(N__35930));
    LocalMux I__7620 (
            .O(N__35930),
            .I(\delay_measurement_inst.delay_tr_timer.N_347 ));
    CascadeMux I__7619 (
            .O(N__35927),
            .I(\delay_measurement_inst.delay_tr_timer.N_347_cascade_ ));
    CascadeMux I__7618 (
            .O(N__35924),
            .I(N__35921));
    InMux I__7617 (
            .O(N__35921),
            .I(N__35915));
    InMux I__7616 (
            .O(N__35920),
            .I(N__35915));
    LocalMux I__7615 (
            .O(N__35915),
            .I(N__35911));
    InMux I__7614 (
            .O(N__35914),
            .I(N__35908));
    Span4Mux_h I__7613 (
            .O(N__35911),
            .I(N__35905));
    LocalMux I__7612 (
            .O(N__35908),
            .I(\delay_measurement_inst.delay_tr_timer.N_365 ));
    Odrv4 I__7611 (
            .O(N__35905),
            .I(\delay_measurement_inst.delay_tr_timer.N_365 ));
    InMux I__7610 (
            .O(N__35900),
            .I(N__35897));
    LocalMux I__7609 (
            .O(N__35897),
            .I(N__35894));
    Odrv4 I__7608 (
            .O(N__35894),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__7607 (
            .O(N__35891),
            .I(N__35888));
    LocalMux I__7606 (
            .O(N__35888),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__7605 (
            .O(N__35885),
            .I(N__35882));
    InMux I__7604 (
            .O(N__35882),
            .I(N__35879));
    LocalMux I__7603 (
            .O(N__35879),
            .I(N__35874));
    InMux I__7602 (
            .O(N__35878),
            .I(N__35871));
    CascadeMux I__7601 (
            .O(N__35877),
            .I(N__35868));
    Span4Mux_h I__7600 (
            .O(N__35874),
            .I(N__35864));
    LocalMux I__7599 (
            .O(N__35871),
            .I(N__35861));
    InMux I__7598 (
            .O(N__35868),
            .I(N__35858));
    InMux I__7597 (
            .O(N__35867),
            .I(N__35855));
    Span4Mux_h I__7596 (
            .O(N__35864),
            .I(N__35850));
    Span4Mux_v I__7595 (
            .O(N__35861),
            .I(N__35850));
    LocalMux I__7594 (
            .O(N__35858),
            .I(N__35845));
    LocalMux I__7593 (
            .O(N__35855),
            .I(N__35845));
    Span4Mux_v I__7592 (
            .O(N__35850),
            .I(N__35842));
    Span4Mux_h I__7591 (
            .O(N__35845),
            .I(N__35839));
    Odrv4 I__7590 (
            .O(N__35842),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__7589 (
            .O(N__35839),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__7588 (
            .O(N__35834),
            .I(N__35822));
    CascadeMux I__7587 (
            .O(N__35833),
            .I(N__35815));
    InMux I__7586 (
            .O(N__35832),
            .I(N__35801));
    InMux I__7585 (
            .O(N__35831),
            .I(N__35801));
    InMux I__7584 (
            .O(N__35830),
            .I(N__35801));
    InMux I__7583 (
            .O(N__35829),
            .I(N__35801));
    InMux I__7582 (
            .O(N__35828),
            .I(N__35796));
    InMux I__7581 (
            .O(N__35827),
            .I(N__35796));
    InMux I__7580 (
            .O(N__35826),
            .I(N__35791));
    InMux I__7579 (
            .O(N__35825),
            .I(N__35791));
    LocalMux I__7578 (
            .O(N__35822),
            .I(N__35788));
    InMux I__7577 (
            .O(N__35821),
            .I(N__35779));
    InMux I__7576 (
            .O(N__35820),
            .I(N__35779));
    InMux I__7575 (
            .O(N__35819),
            .I(N__35779));
    InMux I__7574 (
            .O(N__35818),
            .I(N__35779));
    InMux I__7573 (
            .O(N__35815),
            .I(N__35767));
    InMux I__7572 (
            .O(N__35814),
            .I(N__35767));
    InMux I__7571 (
            .O(N__35813),
            .I(N__35767));
    InMux I__7570 (
            .O(N__35812),
            .I(N__35767));
    InMux I__7569 (
            .O(N__35811),
            .I(N__35767));
    InMux I__7568 (
            .O(N__35810),
            .I(N__35764));
    LocalMux I__7567 (
            .O(N__35801),
            .I(N__35751));
    LocalMux I__7566 (
            .O(N__35796),
            .I(N__35751));
    LocalMux I__7565 (
            .O(N__35791),
            .I(N__35751));
    Span4Mux_v I__7564 (
            .O(N__35788),
            .I(N__35748));
    LocalMux I__7563 (
            .O(N__35779),
            .I(N__35745));
    InMux I__7562 (
            .O(N__35778),
            .I(N__35742));
    LocalMux I__7561 (
            .O(N__35767),
            .I(N__35731));
    LocalMux I__7560 (
            .O(N__35764),
            .I(N__35731));
    InMux I__7559 (
            .O(N__35763),
            .I(N__35718));
    InMux I__7558 (
            .O(N__35762),
            .I(N__35718));
    InMux I__7557 (
            .O(N__35761),
            .I(N__35718));
    InMux I__7556 (
            .O(N__35760),
            .I(N__35718));
    InMux I__7555 (
            .O(N__35759),
            .I(N__35718));
    InMux I__7554 (
            .O(N__35758),
            .I(N__35718));
    Span4Mux_v I__7553 (
            .O(N__35751),
            .I(N__35715));
    Sp12to4 I__7552 (
            .O(N__35748),
            .I(N__35712));
    Span4Mux_v I__7551 (
            .O(N__35745),
            .I(N__35707));
    LocalMux I__7550 (
            .O(N__35742),
            .I(N__35707));
    InMux I__7549 (
            .O(N__35741),
            .I(N__35694));
    InMux I__7548 (
            .O(N__35740),
            .I(N__35694));
    InMux I__7547 (
            .O(N__35739),
            .I(N__35694));
    InMux I__7546 (
            .O(N__35738),
            .I(N__35694));
    InMux I__7545 (
            .O(N__35737),
            .I(N__35694));
    InMux I__7544 (
            .O(N__35736),
            .I(N__35694));
    Span4Mux_h I__7543 (
            .O(N__35731),
            .I(N__35691));
    LocalMux I__7542 (
            .O(N__35718),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__7541 (
            .O(N__35715),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__7540 (
            .O(N__35712),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__7539 (
            .O(N__35707),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__7538 (
            .O(N__35694),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__7537 (
            .O(N__35691),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__7536 (
            .O(N__35678),
            .I(N__35666));
    InMux I__7535 (
            .O(N__35677),
            .I(N__35666));
    InMux I__7534 (
            .O(N__35676),
            .I(N__35661));
    InMux I__7533 (
            .O(N__35675),
            .I(N__35661));
    CascadeMux I__7532 (
            .O(N__35674),
            .I(N__35658));
    CascadeMux I__7531 (
            .O(N__35673),
            .I(N__35655));
    CascadeMux I__7530 (
            .O(N__35672),
            .I(N__35639));
    CascadeMux I__7529 (
            .O(N__35671),
            .I(N__35636));
    LocalMux I__7528 (
            .O(N__35666),
            .I(N__35626));
    LocalMux I__7527 (
            .O(N__35661),
            .I(N__35623));
    InMux I__7526 (
            .O(N__35658),
            .I(N__35610));
    InMux I__7525 (
            .O(N__35655),
            .I(N__35610));
    InMux I__7524 (
            .O(N__35654),
            .I(N__35610));
    InMux I__7523 (
            .O(N__35653),
            .I(N__35610));
    InMux I__7522 (
            .O(N__35652),
            .I(N__35610));
    InMux I__7521 (
            .O(N__35651),
            .I(N__35610));
    InMux I__7520 (
            .O(N__35650),
            .I(N__35599));
    InMux I__7519 (
            .O(N__35649),
            .I(N__35599));
    InMux I__7518 (
            .O(N__35648),
            .I(N__35599));
    InMux I__7517 (
            .O(N__35647),
            .I(N__35599));
    InMux I__7516 (
            .O(N__35646),
            .I(N__35599));
    InMux I__7515 (
            .O(N__35645),
            .I(N__35590));
    InMux I__7514 (
            .O(N__35644),
            .I(N__35590));
    InMux I__7513 (
            .O(N__35643),
            .I(N__35590));
    InMux I__7512 (
            .O(N__35642),
            .I(N__35590));
    InMux I__7511 (
            .O(N__35639),
            .I(N__35575));
    InMux I__7510 (
            .O(N__35636),
            .I(N__35575));
    InMux I__7509 (
            .O(N__35635),
            .I(N__35575));
    InMux I__7508 (
            .O(N__35634),
            .I(N__35575));
    InMux I__7507 (
            .O(N__35633),
            .I(N__35575));
    InMux I__7506 (
            .O(N__35632),
            .I(N__35570));
    InMux I__7505 (
            .O(N__35631),
            .I(N__35570));
    InMux I__7504 (
            .O(N__35630),
            .I(N__35565));
    InMux I__7503 (
            .O(N__35629),
            .I(N__35565));
    Span4Mux_v I__7502 (
            .O(N__35626),
            .I(N__35562));
    Span4Mux_v I__7501 (
            .O(N__35623),
            .I(N__35557));
    LocalMux I__7500 (
            .O(N__35610),
            .I(N__35557));
    LocalMux I__7499 (
            .O(N__35599),
            .I(N__35552));
    LocalMux I__7498 (
            .O(N__35590),
            .I(N__35552));
    InMux I__7497 (
            .O(N__35589),
            .I(N__35543));
    InMux I__7496 (
            .O(N__35588),
            .I(N__35543));
    InMux I__7495 (
            .O(N__35587),
            .I(N__35543));
    InMux I__7494 (
            .O(N__35586),
            .I(N__35543));
    LocalMux I__7493 (
            .O(N__35575),
            .I(N__35538));
    LocalMux I__7492 (
            .O(N__35570),
            .I(N__35538));
    LocalMux I__7491 (
            .O(N__35565),
            .I(N__35535));
    Span4Mux_h I__7490 (
            .O(N__35562),
            .I(N__35528));
    Span4Mux_v I__7489 (
            .O(N__35557),
            .I(N__35528));
    Span4Mux_v I__7488 (
            .O(N__35552),
            .I(N__35528));
    LocalMux I__7487 (
            .O(N__35543),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__7486 (
            .O(N__35538),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__7485 (
            .O(N__35535),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__7484 (
            .O(N__35528),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    CascadeMux I__7483 (
            .O(N__35519),
            .I(N__35501));
    CascadeMux I__7482 (
            .O(N__35518),
            .I(N__35498));
    CascadeMux I__7481 (
            .O(N__35517),
            .I(N__35495));
    CascadeMux I__7480 (
            .O(N__35516),
            .I(N__35489));
    CascadeMux I__7479 (
            .O(N__35515),
            .I(N__35486));
    CascadeMux I__7478 (
            .O(N__35514),
            .I(N__35483));
    CascadeMux I__7477 (
            .O(N__35513),
            .I(N__35480));
    CascadeMux I__7476 (
            .O(N__35512),
            .I(N__35477));
    CascadeMux I__7475 (
            .O(N__35511),
            .I(N__35472));
    CascadeMux I__7474 (
            .O(N__35510),
            .I(N__35469));
    CascadeMux I__7473 (
            .O(N__35509),
            .I(N__35466));
    CascadeMux I__7472 (
            .O(N__35508),
            .I(N__35463));
    CascadeMux I__7471 (
            .O(N__35507),
            .I(N__35459));
    InMux I__7470 (
            .O(N__35506),
            .I(N__35446));
    InMux I__7469 (
            .O(N__35505),
            .I(N__35446));
    InMux I__7468 (
            .O(N__35504),
            .I(N__35446));
    InMux I__7467 (
            .O(N__35501),
            .I(N__35446));
    InMux I__7466 (
            .O(N__35498),
            .I(N__35446));
    InMux I__7465 (
            .O(N__35495),
            .I(N__35446));
    CascadeMux I__7464 (
            .O(N__35494),
            .I(N__35440));
    CascadeMux I__7463 (
            .O(N__35493),
            .I(N__35436));
    CascadeMux I__7462 (
            .O(N__35492),
            .I(N__35433));
    InMux I__7461 (
            .O(N__35489),
            .I(N__35426));
    InMux I__7460 (
            .O(N__35486),
            .I(N__35426));
    InMux I__7459 (
            .O(N__35483),
            .I(N__35419));
    InMux I__7458 (
            .O(N__35480),
            .I(N__35419));
    InMux I__7457 (
            .O(N__35477),
            .I(N__35419));
    InMux I__7456 (
            .O(N__35476),
            .I(N__35410));
    InMux I__7455 (
            .O(N__35475),
            .I(N__35410));
    InMux I__7454 (
            .O(N__35472),
            .I(N__35410));
    InMux I__7453 (
            .O(N__35469),
            .I(N__35410));
    InMux I__7452 (
            .O(N__35466),
            .I(N__35405));
    InMux I__7451 (
            .O(N__35463),
            .I(N__35405));
    InMux I__7450 (
            .O(N__35462),
            .I(N__35400));
    InMux I__7449 (
            .O(N__35459),
            .I(N__35400));
    LocalMux I__7448 (
            .O(N__35446),
            .I(N__35397));
    InMux I__7447 (
            .O(N__35445),
            .I(N__35388));
    InMux I__7446 (
            .O(N__35444),
            .I(N__35388));
    InMux I__7445 (
            .O(N__35443),
            .I(N__35388));
    InMux I__7444 (
            .O(N__35440),
            .I(N__35388));
    InMux I__7443 (
            .O(N__35439),
            .I(N__35377));
    InMux I__7442 (
            .O(N__35436),
            .I(N__35377));
    InMux I__7441 (
            .O(N__35433),
            .I(N__35377));
    InMux I__7440 (
            .O(N__35432),
            .I(N__35377));
    InMux I__7439 (
            .O(N__35431),
            .I(N__35377));
    LocalMux I__7438 (
            .O(N__35426),
            .I(N__35372));
    LocalMux I__7437 (
            .O(N__35419),
            .I(N__35372));
    LocalMux I__7436 (
            .O(N__35410),
            .I(N__35365));
    LocalMux I__7435 (
            .O(N__35405),
            .I(N__35365));
    LocalMux I__7434 (
            .O(N__35400),
            .I(N__35365));
    Span4Mux_v I__7433 (
            .O(N__35397),
            .I(N__35360));
    LocalMux I__7432 (
            .O(N__35388),
            .I(N__35360));
    LocalMux I__7431 (
            .O(N__35377),
            .I(N__35355));
    Span4Mux_h I__7430 (
            .O(N__35372),
            .I(N__35355));
    Span4Mux_h I__7429 (
            .O(N__35365),
            .I(N__35352));
    Span4Mux_h I__7428 (
            .O(N__35360),
            .I(N__35349));
    Span4Mux_h I__7427 (
            .O(N__35355),
            .I(N__35346));
    Odrv4 I__7426 (
            .O(N__35352),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    Odrv4 I__7425 (
            .O(N__35349),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    Odrv4 I__7424 (
            .O(N__35346),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    InMux I__7423 (
            .O(N__35339),
            .I(N__35336));
    LocalMux I__7422 (
            .O(N__35336),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    CascadeMux I__7421 (
            .O(N__35333),
            .I(N__35330));
    InMux I__7420 (
            .O(N__35330),
            .I(N__35325));
    InMux I__7419 (
            .O(N__35329),
            .I(N__35322));
    CascadeMux I__7418 (
            .O(N__35328),
            .I(N__35318));
    LocalMux I__7417 (
            .O(N__35325),
            .I(N__35315));
    LocalMux I__7416 (
            .O(N__35322),
            .I(N__35312));
    InMux I__7415 (
            .O(N__35321),
            .I(N__35307));
    InMux I__7414 (
            .O(N__35318),
            .I(N__35307));
    Span4Mux_v I__7413 (
            .O(N__35315),
            .I(N__35303));
    Span4Mux_v I__7412 (
            .O(N__35312),
            .I(N__35300));
    LocalMux I__7411 (
            .O(N__35307),
            .I(N__35297));
    InMux I__7410 (
            .O(N__35306),
            .I(N__35294));
    Span4Mux_h I__7409 (
            .O(N__35303),
            .I(N__35291));
    Sp12to4 I__7408 (
            .O(N__35300),
            .I(N__35286));
    Span12Mux_s8_v I__7407 (
            .O(N__35297),
            .I(N__35286));
    LocalMux I__7406 (
            .O(N__35294),
            .I(N__35283));
    Odrv4 I__7405 (
            .O(N__35291),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv12 I__7404 (
            .O(N__35286),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__7403 (
            .O(N__35283),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__7402 (
            .O(N__35276),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ));
    InMux I__7401 (
            .O(N__35273),
            .I(N__35269));
    InMux I__7400 (
            .O(N__35272),
            .I(N__35266));
    LocalMux I__7399 (
            .O(N__35269),
            .I(N__35261));
    LocalMux I__7398 (
            .O(N__35266),
            .I(N__35261));
    Odrv4 I__7397 (
            .O(N__35261),
            .I(\delay_measurement_inst.delay_tr_timer.N_380 ));
    InMux I__7396 (
            .O(N__35258),
            .I(N__35255));
    LocalMux I__7395 (
            .O(N__35255),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ));
    InMux I__7394 (
            .O(N__35252),
            .I(N__35246));
    InMux I__7393 (
            .O(N__35251),
            .I(N__35246));
    LocalMux I__7392 (
            .O(N__35246),
            .I(\delay_measurement_inst.delay_tr_timer.N_341 ));
    InMux I__7391 (
            .O(N__35243),
            .I(N__35240));
    LocalMux I__7390 (
            .O(N__35240),
            .I(\delay_measurement_inst.delay_tr_timer.N_367 ));
    InMux I__7389 (
            .O(N__35237),
            .I(N__35234));
    LocalMux I__7388 (
            .O(N__35234),
            .I(N__35231));
    Odrv4 I__7387 (
            .O(N__35231),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    CascadeMux I__7386 (
            .O(N__35228),
            .I(N__35225));
    InMux I__7385 (
            .O(N__35225),
            .I(N__35222));
    LocalMux I__7384 (
            .O(N__35222),
            .I(N__35218));
    InMux I__7383 (
            .O(N__35221),
            .I(N__35214));
    Span4Mux_v I__7382 (
            .O(N__35218),
            .I(N__35211));
    InMux I__7381 (
            .O(N__35217),
            .I(N__35208));
    LocalMux I__7380 (
            .O(N__35214),
            .I(N__35203));
    Span4Mux_h I__7379 (
            .O(N__35211),
            .I(N__35198));
    LocalMux I__7378 (
            .O(N__35208),
            .I(N__35198));
    InMux I__7377 (
            .O(N__35207),
            .I(N__35193));
    InMux I__7376 (
            .O(N__35206),
            .I(N__35193));
    Span4Mux_v I__7375 (
            .O(N__35203),
            .I(N__35188));
    Span4Mux_h I__7374 (
            .O(N__35198),
            .I(N__35188));
    LocalMux I__7373 (
            .O(N__35193),
            .I(N__35185));
    Odrv4 I__7372 (
            .O(N__35188),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__7371 (
            .O(N__35185),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__7370 (
            .O(N__35180),
            .I(N__35177));
    LocalMux I__7369 (
            .O(N__35177),
            .I(N__35174));
    Odrv4 I__7368 (
            .O(N__35174),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    CascadeMux I__7367 (
            .O(N__35171),
            .I(N__35167));
    InMux I__7366 (
            .O(N__35170),
            .I(N__35163));
    InMux I__7365 (
            .O(N__35167),
            .I(N__35160));
    InMux I__7364 (
            .O(N__35166),
            .I(N__35157));
    LocalMux I__7363 (
            .O(N__35163),
            .I(N__35153));
    LocalMux I__7362 (
            .O(N__35160),
            .I(N__35150));
    LocalMux I__7361 (
            .O(N__35157),
            .I(N__35146));
    InMux I__7360 (
            .O(N__35156),
            .I(N__35143));
    Span4Mux_v I__7359 (
            .O(N__35153),
            .I(N__35140));
    Span12Mux_h I__7358 (
            .O(N__35150),
            .I(N__35137));
    InMux I__7357 (
            .O(N__35149),
            .I(N__35134));
    Span4Mux_h I__7356 (
            .O(N__35146),
            .I(N__35129));
    LocalMux I__7355 (
            .O(N__35143),
            .I(N__35129));
    Odrv4 I__7354 (
            .O(N__35140),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv12 I__7353 (
            .O(N__35137),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__7352 (
            .O(N__35134),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__7351 (
            .O(N__35129),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__7350 (
            .O(N__35120),
            .I(N__35117));
    LocalMux I__7349 (
            .O(N__35117),
            .I(N__35114));
    Odrv4 I__7348 (
            .O(N__35114),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__7347 (
            .O(N__35111),
            .I(N__35107));
    InMux I__7346 (
            .O(N__35110),
            .I(N__35104));
    LocalMux I__7345 (
            .O(N__35107),
            .I(N__35101));
    LocalMux I__7344 (
            .O(N__35104),
            .I(N__35096));
    Span4Mux_h I__7343 (
            .O(N__35101),
            .I(N__35093));
    InMux I__7342 (
            .O(N__35100),
            .I(N__35090));
    InMux I__7341 (
            .O(N__35099),
            .I(N__35087));
    Span4Mux_v I__7340 (
            .O(N__35096),
            .I(N__35080));
    Span4Mux_v I__7339 (
            .O(N__35093),
            .I(N__35080));
    LocalMux I__7338 (
            .O(N__35090),
            .I(N__35080));
    LocalMux I__7337 (
            .O(N__35087),
            .I(N__35076));
    Span4Mux_h I__7336 (
            .O(N__35080),
            .I(N__35073));
    InMux I__7335 (
            .O(N__35079),
            .I(N__35070));
    Odrv12 I__7334 (
            .O(N__35076),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__7333 (
            .O(N__35073),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__7332 (
            .O(N__35070),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__7331 (
            .O(N__35063),
            .I(N__35060));
    LocalMux I__7330 (
            .O(N__35060),
            .I(N__35057));
    Odrv4 I__7329 (
            .O(N__35057),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    CascadeMux I__7328 (
            .O(N__35054),
            .I(N__35051));
    InMux I__7327 (
            .O(N__35051),
            .I(N__35048));
    LocalMux I__7326 (
            .O(N__35048),
            .I(N__35044));
    InMux I__7325 (
            .O(N__35047),
            .I(N__35039));
    Span4Mux_v I__7324 (
            .O(N__35044),
            .I(N__35035));
    InMux I__7323 (
            .O(N__35043),
            .I(N__35032));
    CascadeMux I__7322 (
            .O(N__35042),
            .I(N__35029));
    LocalMux I__7321 (
            .O(N__35039),
            .I(N__35026));
    InMux I__7320 (
            .O(N__35038),
            .I(N__35023));
    Span4Mux_h I__7319 (
            .O(N__35035),
            .I(N__35018));
    LocalMux I__7318 (
            .O(N__35032),
            .I(N__35018));
    InMux I__7317 (
            .O(N__35029),
            .I(N__35015));
    Span4Mux_v I__7316 (
            .O(N__35026),
            .I(N__35012));
    LocalMux I__7315 (
            .O(N__35023),
            .I(N__35009));
    Span4Mux_h I__7314 (
            .O(N__35018),
            .I(N__35006));
    LocalMux I__7313 (
            .O(N__35015),
            .I(N__35003));
    Odrv4 I__7312 (
            .O(N__35012),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv12 I__7311 (
            .O(N__35009),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__7310 (
            .O(N__35006),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv12 I__7309 (
            .O(N__35003),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__7308 (
            .O(N__34994),
            .I(N__34990));
    InMux I__7307 (
            .O(N__34993),
            .I(N__34987));
    LocalMux I__7306 (
            .O(N__34990),
            .I(N__34983));
    LocalMux I__7305 (
            .O(N__34987),
            .I(N__34980));
    InMux I__7304 (
            .O(N__34986),
            .I(N__34977));
    Span4Mux_h I__7303 (
            .O(N__34983),
            .I(N__34974));
    Span4Mux_v I__7302 (
            .O(N__34980),
            .I(N__34971));
    LocalMux I__7301 (
            .O(N__34977),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv4 I__7300 (
            .O(N__34974),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv4 I__7299 (
            .O(N__34971),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    CascadeMux I__7298 (
            .O(N__34964),
            .I(N__34956));
    CascadeMux I__7297 (
            .O(N__34963),
            .I(N__34950));
    CascadeMux I__7296 (
            .O(N__34962),
            .I(N__34944));
    CascadeMux I__7295 (
            .O(N__34961),
            .I(N__34939));
    CascadeMux I__7294 (
            .O(N__34960),
            .I(N__34934));
    CascadeMux I__7293 (
            .O(N__34959),
            .I(N__34930));
    InMux I__7292 (
            .O(N__34956),
            .I(N__34927));
    CascadeMux I__7291 (
            .O(N__34955),
            .I(N__34923));
    CascadeMux I__7290 (
            .O(N__34954),
            .I(N__34920));
    CascadeMux I__7289 (
            .O(N__34953),
            .I(N__34917));
    InMux I__7288 (
            .O(N__34950),
            .I(N__34909));
    CascadeMux I__7287 (
            .O(N__34949),
            .I(N__34906));
    CascadeMux I__7286 (
            .O(N__34948),
            .I(N__34902));
    InMux I__7285 (
            .O(N__34947),
            .I(N__34894));
    InMux I__7284 (
            .O(N__34944),
            .I(N__34891));
    CascadeMux I__7283 (
            .O(N__34943),
            .I(N__34887));
    InMux I__7282 (
            .O(N__34942),
            .I(N__34869));
    InMux I__7281 (
            .O(N__34939),
            .I(N__34851));
    InMux I__7280 (
            .O(N__34938),
            .I(N__34851));
    InMux I__7279 (
            .O(N__34937),
            .I(N__34851));
    InMux I__7278 (
            .O(N__34934),
            .I(N__34851));
    InMux I__7277 (
            .O(N__34933),
            .I(N__34851));
    InMux I__7276 (
            .O(N__34930),
            .I(N__34851));
    LocalMux I__7275 (
            .O(N__34927),
            .I(N__34848));
    InMux I__7274 (
            .O(N__34926),
            .I(N__34839));
    InMux I__7273 (
            .O(N__34923),
            .I(N__34839));
    InMux I__7272 (
            .O(N__34920),
            .I(N__34839));
    InMux I__7271 (
            .O(N__34917),
            .I(N__34839));
    InMux I__7270 (
            .O(N__34916),
            .I(N__34834));
    InMux I__7269 (
            .O(N__34915),
            .I(N__34834));
    InMux I__7268 (
            .O(N__34914),
            .I(N__34826));
    InMux I__7267 (
            .O(N__34913),
            .I(N__34826));
    InMux I__7266 (
            .O(N__34912),
            .I(N__34826));
    LocalMux I__7265 (
            .O(N__34909),
            .I(N__34823));
    InMux I__7264 (
            .O(N__34906),
            .I(N__34806));
    InMux I__7263 (
            .O(N__34905),
            .I(N__34806));
    InMux I__7262 (
            .O(N__34902),
            .I(N__34806));
    InMux I__7261 (
            .O(N__34901),
            .I(N__34806));
    InMux I__7260 (
            .O(N__34900),
            .I(N__34806));
    InMux I__7259 (
            .O(N__34899),
            .I(N__34806));
    InMux I__7258 (
            .O(N__34898),
            .I(N__34806));
    InMux I__7257 (
            .O(N__34897),
            .I(N__34806));
    LocalMux I__7256 (
            .O(N__34894),
            .I(N__34801));
    LocalMux I__7255 (
            .O(N__34891),
            .I(N__34801));
    InMux I__7254 (
            .O(N__34890),
            .I(N__34798));
    InMux I__7253 (
            .O(N__34887),
            .I(N__34787));
    InMux I__7252 (
            .O(N__34886),
            .I(N__34787));
    InMux I__7251 (
            .O(N__34885),
            .I(N__34787));
    InMux I__7250 (
            .O(N__34884),
            .I(N__34787));
    InMux I__7249 (
            .O(N__34883),
            .I(N__34787));
    InMux I__7248 (
            .O(N__34882),
            .I(N__34782));
    InMux I__7247 (
            .O(N__34881),
            .I(N__34782));
    InMux I__7246 (
            .O(N__34880),
            .I(N__34771));
    InMux I__7245 (
            .O(N__34879),
            .I(N__34771));
    InMux I__7244 (
            .O(N__34878),
            .I(N__34771));
    InMux I__7243 (
            .O(N__34877),
            .I(N__34771));
    InMux I__7242 (
            .O(N__34876),
            .I(N__34771));
    InMux I__7241 (
            .O(N__34875),
            .I(N__34766));
    InMux I__7240 (
            .O(N__34874),
            .I(N__34766));
    InMux I__7239 (
            .O(N__34873),
            .I(N__34763));
    InMux I__7238 (
            .O(N__34872),
            .I(N__34760));
    LocalMux I__7237 (
            .O(N__34869),
            .I(N__34757));
    InMux I__7236 (
            .O(N__34868),
            .I(N__34746));
    InMux I__7235 (
            .O(N__34867),
            .I(N__34746));
    InMux I__7234 (
            .O(N__34866),
            .I(N__34746));
    InMux I__7233 (
            .O(N__34865),
            .I(N__34746));
    InMux I__7232 (
            .O(N__34864),
            .I(N__34746));
    LocalMux I__7231 (
            .O(N__34851),
            .I(N__34739));
    Span4Mux_v I__7230 (
            .O(N__34848),
            .I(N__34739));
    LocalMux I__7229 (
            .O(N__34839),
            .I(N__34739));
    LocalMux I__7228 (
            .O(N__34834),
            .I(N__34736));
    InMux I__7227 (
            .O(N__34833),
            .I(N__34733));
    LocalMux I__7226 (
            .O(N__34826),
            .I(N__34726));
    Span4Mux_v I__7225 (
            .O(N__34823),
            .I(N__34726));
    LocalMux I__7224 (
            .O(N__34806),
            .I(N__34726));
    Span4Mux_h I__7223 (
            .O(N__34801),
            .I(N__34711));
    LocalMux I__7222 (
            .O(N__34798),
            .I(N__34711));
    LocalMux I__7221 (
            .O(N__34787),
            .I(N__34711));
    LocalMux I__7220 (
            .O(N__34782),
            .I(N__34711));
    LocalMux I__7219 (
            .O(N__34771),
            .I(N__34711));
    LocalMux I__7218 (
            .O(N__34766),
            .I(N__34711));
    LocalMux I__7217 (
            .O(N__34763),
            .I(N__34711));
    LocalMux I__7216 (
            .O(N__34760),
            .I(N__34708));
    Span4Mux_h I__7215 (
            .O(N__34757),
            .I(N__34703));
    LocalMux I__7214 (
            .O(N__34746),
            .I(N__34703));
    Span4Mux_v I__7213 (
            .O(N__34739),
            .I(N__34698));
    Span4Mux_v I__7212 (
            .O(N__34736),
            .I(N__34698));
    LocalMux I__7211 (
            .O(N__34733),
            .I(N__34691));
    Span4Mux_h I__7210 (
            .O(N__34726),
            .I(N__34691));
    Span4Mux_v I__7209 (
            .O(N__34711),
            .I(N__34691));
    Odrv4 I__7208 (
            .O(N__34708),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__7207 (
            .O(N__34703),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__7206 (
            .O(N__34698),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__7205 (
            .O(N__34691),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__7204 (
            .O(N__34682),
            .I(N__34679));
    LocalMux I__7203 (
            .O(N__34679),
            .I(N__34676));
    Span4Mux_h I__7202 (
            .O(N__34676),
            .I(N__34673));
    Odrv4 I__7201 (
            .O(N__34673),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_10 ));
    CascadeMux I__7200 (
            .O(N__34670),
            .I(N__34667));
    InMux I__7199 (
            .O(N__34667),
            .I(N__34664));
    LocalMux I__7198 (
            .O(N__34664),
            .I(N__34661));
    Odrv4 I__7197 (
            .O(N__34661),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ));
    InMux I__7196 (
            .O(N__34658),
            .I(N__34655));
    LocalMux I__7195 (
            .O(N__34655),
            .I(N__34652));
    Odrv4 I__7194 (
            .O(N__34652),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    CascadeMux I__7193 (
            .O(N__34649),
            .I(N__34646));
    InMux I__7192 (
            .O(N__34646),
            .I(N__34641));
    InMux I__7191 (
            .O(N__34645),
            .I(N__34638));
    InMux I__7190 (
            .O(N__34644),
            .I(N__34635));
    LocalMux I__7189 (
            .O(N__34641),
            .I(N__34632));
    LocalMux I__7188 (
            .O(N__34638),
            .I(N__34627));
    LocalMux I__7187 (
            .O(N__34635),
            .I(N__34622));
    Span4Mux_v I__7186 (
            .O(N__34632),
            .I(N__34622));
    InMux I__7185 (
            .O(N__34631),
            .I(N__34619));
    InMux I__7184 (
            .O(N__34630),
            .I(N__34616));
    Span4Mux_v I__7183 (
            .O(N__34627),
            .I(N__34611));
    Span4Mux_h I__7182 (
            .O(N__34622),
            .I(N__34611));
    LocalMux I__7181 (
            .O(N__34619),
            .I(N__34608));
    LocalMux I__7180 (
            .O(N__34616),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__7179 (
            .O(N__34611),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__7178 (
            .O(N__34608),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__7177 (
            .O(N__34601),
            .I(N__34598));
    LocalMux I__7176 (
            .O(N__34598),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    CascadeMux I__7175 (
            .O(N__34595),
            .I(N__34592));
    InMux I__7174 (
            .O(N__34592),
            .I(N__34589));
    LocalMux I__7173 (
            .O(N__34589),
            .I(N__34585));
    CascadeMux I__7172 (
            .O(N__34588),
            .I(N__34581));
    Span4Mux_v I__7171 (
            .O(N__34585),
            .I(N__34578));
    InMux I__7170 (
            .O(N__34584),
            .I(N__34575));
    InMux I__7169 (
            .O(N__34581),
            .I(N__34572));
    Span4Mux_h I__7168 (
            .O(N__34578),
            .I(N__34567));
    LocalMux I__7167 (
            .O(N__34575),
            .I(N__34567));
    LocalMux I__7166 (
            .O(N__34572),
            .I(N__34563));
    Span4Mux_h I__7165 (
            .O(N__34567),
            .I(N__34560));
    InMux I__7164 (
            .O(N__34566),
            .I(N__34557));
    Span4Mux_h I__7163 (
            .O(N__34563),
            .I(N__34552));
    Span4Mux_v I__7162 (
            .O(N__34560),
            .I(N__34552));
    LocalMux I__7161 (
            .O(N__34557),
            .I(N__34549));
    Odrv4 I__7160 (
            .O(N__34552),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__7159 (
            .O(N__34549),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    CascadeMux I__7158 (
            .O(N__34544),
            .I(N__34541));
    InMux I__7157 (
            .O(N__34541),
            .I(N__34538));
    LocalMux I__7156 (
            .O(N__34538),
            .I(N__34535));
    Odrv4 I__7155 (
            .O(N__34535),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__7154 (
            .O(N__34532),
            .I(N__34529));
    LocalMux I__7153 (
            .O(N__34529),
            .I(N__34524));
    InMux I__7152 (
            .O(N__34528),
            .I(N__34521));
    CascadeMux I__7151 (
            .O(N__34527),
            .I(N__34518));
    Span4Mux_h I__7150 (
            .O(N__34524),
            .I(N__34512));
    LocalMux I__7149 (
            .O(N__34521),
            .I(N__34512));
    InMux I__7148 (
            .O(N__34518),
            .I(N__34507));
    InMux I__7147 (
            .O(N__34517),
            .I(N__34507));
    Span4Mux_v I__7146 (
            .O(N__34512),
            .I(N__34504));
    LocalMux I__7145 (
            .O(N__34507),
            .I(N__34501));
    Span4Mux_h I__7144 (
            .O(N__34504),
            .I(N__34498));
    Span4Mux_h I__7143 (
            .O(N__34501),
            .I(N__34495));
    Odrv4 I__7142 (
            .O(N__34498),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__7141 (
            .O(N__34495),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__7140 (
            .O(N__34490),
            .I(N__34487));
    LocalMux I__7139 (
            .O(N__34487),
            .I(N__34482));
    InMux I__7138 (
            .O(N__34486),
            .I(N__34479));
    InMux I__7137 (
            .O(N__34485),
            .I(N__34475));
    Span4Mux_h I__7136 (
            .O(N__34482),
            .I(N__34470));
    LocalMux I__7135 (
            .O(N__34479),
            .I(N__34470));
    InMux I__7134 (
            .O(N__34478),
            .I(N__34467));
    LocalMux I__7133 (
            .O(N__34475),
            .I(N__34464));
    Span4Mux_h I__7132 (
            .O(N__34470),
            .I(N__34461));
    LocalMux I__7131 (
            .O(N__34467),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__7130 (
            .O(N__34464),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__7129 (
            .O(N__34461),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__7128 (
            .O(N__34454),
            .I(N__34450));
    InMux I__7127 (
            .O(N__34453),
            .I(N__34447));
    LocalMux I__7126 (
            .O(N__34450),
            .I(N__34444));
    LocalMux I__7125 (
            .O(N__34447),
            .I(N__34441));
    Span4Mux_h I__7124 (
            .O(N__34444),
            .I(N__34438));
    Span4Mux_v I__7123 (
            .O(N__34441),
            .I(N__34432));
    Span4Mux_v I__7122 (
            .O(N__34438),
            .I(N__34432));
    InMux I__7121 (
            .O(N__34437),
            .I(N__34429));
    Odrv4 I__7120 (
            .O(N__34432),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    LocalMux I__7119 (
            .O(N__34429),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__7118 (
            .O(N__34424),
            .I(N__34421));
    LocalMux I__7117 (
            .O(N__34421),
            .I(N__34418));
    Span4Mux_h I__7116 (
            .O(N__34418),
            .I(N__34415));
    Span4Mux_v I__7115 (
            .O(N__34415),
            .I(N__34412));
    Odrv4 I__7114 (
            .O(N__34412),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_6 ));
    CascadeMux I__7113 (
            .O(N__34409),
            .I(N__34406));
    InMux I__7112 (
            .O(N__34406),
            .I(N__34403));
    LocalMux I__7111 (
            .O(N__34403),
            .I(N__34400));
    Odrv4 I__7110 (
            .O(N__34400),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ));
    CascadeMux I__7109 (
            .O(N__34397),
            .I(N__34394));
    InMux I__7108 (
            .O(N__34394),
            .I(N__34391));
    LocalMux I__7107 (
            .O(N__34391),
            .I(N__34387));
    InMux I__7106 (
            .O(N__34390),
            .I(N__34382));
    Span4Mux_v I__7105 (
            .O(N__34387),
            .I(N__34378));
    InMux I__7104 (
            .O(N__34386),
            .I(N__34375));
    InMux I__7103 (
            .O(N__34385),
            .I(N__34372));
    LocalMux I__7102 (
            .O(N__34382),
            .I(N__34369));
    InMux I__7101 (
            .O(N__34381),
            .I(N__34366));
    Span4Mux_h I__7100 (
            .O(N__34378),
            .I(N__34359));
    LocalMux I__7099 (
            .O(N__34375),
            .I(N__34359));
    LocalMux I__7098 (
            .O(N__34372),
            .I(N__34359));
    Odrv4 I__7097 (
            .O(N__34369),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__7096 (
            .O(N__34366),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__7095 (
            .O(N__34359),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__7094 (
            .O(N__34352),
            .I(N__34349));
    LocalMux I__7093 (
            .O(N__34349),
            .I(\current_shift_inst.PI_CTRL.integrator_i_14 ));
    CascadeMux I__7092 (
            .O(N__34346),
            .I(N__34343));
    InMux I__7091 (
            .O(N__34343),
            .I(N__34337));
    InMux I__7090 (
            .O(N__34342),
            .I(N__34334));
    InMux I__7089 (
            .O(N__34341),
            .I(N__34331));
    InMux I__7088 (
            .O(N__34340),
            .I(N__34328));
    LocalMux I__7087 (
            .O(N__34337),
            .I(N__34325));
    LocalMux I__7086 (
            .O(N__34334),
            .I(N__34321));
    LocalMux I__7085 (
            .O(N__34331),
            .I(N__34316));
    LocalMux I__7084 (
            .O(N__34328),
            .I(N__34316));
    Span12Mux_v I__7083 (
            .O(N__34325),
            .I(N__34313));
    InMux I__7082 (
            .O(N__34324),
            .I(N__34310));
    Span4Mux_v I__7081 (
            .O(N__34321),
            .I(N__34307));
    Span4Mux_v I__7080 (
            .O(N__34316),
            .I(N__34304));
    Odrv12 I__7079 (
            .O(N__34313),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__7078 (
            .O(N__34310),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__7077 (
            .O(N__34307),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__7076 (
            .O(N__34304),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    CascadeMux I__7075 (
            .O(N__34295),
            .I(N__34292));
    InMux I__7074 (
            .O(N__34292),
            .I(N__34289));
    LocalMux I__7073 (
            .O(N__34289),
            .I(N__34286));
    Odrv4 I__7072 (
            .O(N__34286),
            .I(\current_shift_inst.PI_CTRL.integrator_i_19 ));
    InMux I__7071 (
            .O(N__34283),
            .I(N__34280));
    LocalMux I__7070 (
            .O(N__34280),
            .I(N__34277));
    Odrv12 I__7069 (
            .O(N__34277),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7 ));
    InMux I__7068 (
            .O(N__34274),
            .I(N__34271));
    LocalMux I__7067 (
            .O(N__34271),
            .I(N__34268));
    Odrv4 I__7066 (
            .O(N__34268),
            .I(\current_shift_inst.PI_CTRL.integrator_i_24 ));
    InMux I__7065 (
            .O(N__34265),
            .I(N__34262));
    LocalMux I__7064 (
            .O(N__34262),
            .I(\current_shift_inst.PI_CTRL.integrator_i_6 ));
    InMux I__7063 (
            .O(N__34259),
            .I(N__34256));
    LocalMux I__7062 (
            .O(N__34256),
            .I(\current_shift_inst.PI_CTRL.integrator_i_10 ));
    InMux I__7061 (
            .O(N__34253),
            .I(N__34250));
    LocalMux I__7060 (
            .O(N__34250),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__7059 (
            .O(N__34247),
            .I(N__34244));
    LocalMux I__7058 (
            .O(N__34244),
            .I(N__34241));
    Span4Mux_h I__7057 (
            .O(N__34241),
            .I(N__34238));
    Span4Mux_h I__7056 (
            .O(N__34238),
            .I(N__34235));
    Odrv4 I__7055 (
            .O(N__34235),
            .I(\current_shift_inst.PI_CTRL.N_74_16 ));
    CascadeMux I__7054 (
            .O(N__34232),
            .I(N__34229));
    InMux I__7053 (
            .O(N__34229),
            .I(N__34224));
    InMux I__7052 (
            .O(N__34228),
            .I(N__34219));
    InMux I__7051 (
            .O(N__34227),
            .I(N__34216));
    LocalMux I__7050 (
            .O(N__34224),
            .I(N__34213));
    InMux I__7049 (
            .O(N__34223),
            .I(N__34210));
    InMux I__7048 (
            .O(N__34222),
            .I(N__34207));
    LocalMux I__7047 (
            .O(N__34219),
            .I(N__34202));
    LocalMux I__7046 (
            .O(N__34216),
            .I(N__34202));
    Span4Mux_v I__7045 (
            .O(N__34213),
            .I(N__34197));
    LocalMux I__7044 (
            .O(N__34210),
            .I(N__34197));
    LocalMux I__7043 (
            .O(N__34207),
            .I(N__34194));
    Span4Mux_v I__7042 (
            .O(N__34202),
            .I(N__34188));
    Span4Mux_h I__7041 (
            .O(N__34197),
            .I(N__34188));
    Span4Mux_v I__7040 (
            .O(N__34194),
            .I(N__34185));
    InMux I__7039 (
            .O(N__34193),
            .I(N__34182));
    Span4Mux_h I__7038 (
            .O(N__34188),
            .I(N__34179));
    Odrv4 I__7037 (
            .O(N__34185),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__7036 (
            .O(N__34182),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__7035 (
            .O(N__34179),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    CascadeMux I__7034 (
            .O(N__34172),
            .I(N__34169));
    InMux I__7033 (
            .O(N__34169),
            .I(N__34166));
    LocalMux I__7032 (
            .O(N__34166),
            .I(N__34163));
    Odrv12 I__7031 (
            .O(N__34163),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ));
    InMux I__7030 (
            .O(N__34160),
            .I(N__34157));
    LocalMux I__7029 (
            .O(N__34157),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__7028 (
            .O(N__34154),
            .I(N__34151));
    LocalMux I__7027 (
            .O(N__34151),
            .I(N__34148));
    Odrv12 I__7026 (
            .O(N__34148),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__7025 (
            .O(N__34145),
            .I(N__34142));
    LocalMux I__7024 (
            .O(N__34142),
            .I(N__34139));
    Odrv12 I__7023 (
            .O(N__34139),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__7022 (
            .O(N__34136),
            .I(N__34133));
    LocalMux I__7021 (
            .O(N__34133),
            .I(N__34130));
    Odrv12 I__7020 (
            .O(N__34130),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__7019 (
            .O(N__34127),
            .I(N__34124));
    LocalMux I__7018 (
            .O(N__34124),
            .I(N__34121));
    Odrv4 I__7017 (
            .O(N__34121),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__7016 (
            .O(N__34118),
            .I(N__34115));
    LocalMux I__7015 (
            .O(N__34115),
            .I(N__34112));
    Odrv12 I__7014 (
            .O(N__34112),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__7013 (
            .O(N__34109),
            .I(N__34106));
    LocalMux I__7012 (
            .O(N__34106),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    ClkMux I__7011 (
            .O(N__34103),
            .I(N__34100));
    GlobalMux I__7010 (
            .O(N__34100),
            .I(N__34097));
    gio2CtrlBuf I__7009 (
            .O(N__34097),
            .I(delay_tr_input_c_g));
    InMux I__7008 (
            .O(N__34094),
            .I(N__34091));
    LocalMux I__7007 (
            .O(N__34091),
            .I(N__34088));
    Odrv4 I__7006 (
            .O(N__34088),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__7005 (
            .O(N__34085),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__7004 (
            .O(N__34082),
            .I(N__34079));
    LocalMux I__7003 (
            .O(N__34079),
            .I(N__34076));
    Odrv4 I__7002 (
            .O(N__34076),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__7001 (
            .O(N__34073),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__7000 (
            .O(N__34070),
            .I(bfn_15_20_0_));
    InMux I__6999 (
            .O(N__34067),
            .I(N__34064));
    LocalMux I__6998 (
            .O(N__34064),
            .I(N__34061));
    Odrv4 I__6997 (
            .O(N__34061),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__6996 (
            .O(N__34058),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__6995 (
            .O(N__34055),
            .I(N__34052));
    LocalMux I__6994 (
            .O(N__34052),
            .I(N__34049));
    Odrv4 I__6993 (
            .O(N__34049),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__6992 (
            .O(N__34046),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__6991 (
            .O(N__34043),
            .I(N__34040));
    LocalMux I__6990 (
            .O(N__34040),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    CascadeMux I__6989 (
            .O(N__34037),
            .I(N__34034));
    InMux I__6988 (
            .O(N__34034),
            .I(N__34028));
    InMux I__6987 (
            .O(N__34033),
            .I(N__34028));
    LocalMux I__6986 (
            .O(N__34028),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__6985 (
            .O(N__34025),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__6984 (
            .O(N__34022),
            .I(N__34019));
    LocalMux I__6983 (
            .O(N__34019),
            .I(N__34016));
    Odrv4 I__6982 (
            .O(N__34016),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__6981 (
            .O(N__34013),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__6980 (
            .O(N__34010),
            .I(\current_shift_inst.un4_control_input1_31 ));
    InMux I__6979 (
            .O(N__34007),
            .I(N__34004));
    LocalMux I__6978 (
            .O(N__34004),
            .I(N__34001));
    Span4Mux_h I__6977 (
            .O(N__34001),
            .I(N__33998));
    Odrv4 I__6976 (
            .O(N__33998),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__6975 (
            .O(N__33995),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ));
    InMux I__6974 (
            .O(N__33992),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__6973 (
            .O(N__33989),
            .I(N__33986));
    LocalMux I__6972 (
            .O(N__33986),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__6971 (
            .O(N__33983),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__6970 (
            .O(N__33980),
            .I(N__33977));
    LocalMux I__6969 (
            .O(N__33977),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__6968 (
            .O(N__33974),
            .I(bfn_15_19_0_));
    CascadeMux I__6967 (
            .O(N__33971),
            .I(N__33968));
    InMux I__6966 (
            .O(N__33968),
            .I(N__33965));
    LocalMux I__6965 (
            .O(N__33965),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__6964 (
            .O(N__33962),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__6963 (
            .O(N__33959),
            .I(N__33956));
    LocalMux I__6962 (
            .O(N__33956),
            .I(N__33953));
    Span4Mux_h I__6961 (
            .O(N__33953),
            .I(N__33950));
    Odrv4 I__6960 (
            .O(N__33950),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__6959 (
            .O(N__33947),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__6958 (
            .O(N__33944),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__6957 (
            .O(N__33941),
            .I(N__33938));
    LocalMux I__6956 (
            .O(N__33938),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__6955 (
            .O(N__33935),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__6954 (
            .O(N__33932),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__6953 (
            .O(N__33929),
            .I(N__33926));
    LocalMux I__6952 (
            .O(N__33926),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__6951 (
            .O(N__33923),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__6950 (
            .O(N__33920),
            .I(N__33917));
    LocalMux I__6949 (
            .O(N__33917),
            .I(N__33914));
    Odrv4 I__6948 (
            .O(N__33914),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__6947 (
            .O(N__33911),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__6946 (
            .O(N__33908),
            .I(N__33905));
    LocalMux I__6945 (
            .O(N__33905),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__6944 (
            .O(N__33902),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__6943 (
            .O(N__33899),
            .I(N__33896));
    LocalMux I__6942 (
            .O(N__33896),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__6941 (
            .O(N__33893),
            .I(bfn_15_18_0_));
    InMux I__6940 (
            .O(N__33890),
            .I(N__33887));
    LocalMux I__6939 (
            .O(N__33887),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__6938 (
            .O(N__33884),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__6937 (
            .O(N__33881),
            .I(N__33878));
    LocalMux I__6936 (
            .O(N__33878),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__6935 (
            .O(N__33875),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__6934 (
            .O(N__33872),
            .I(N__33869));
    LocalMux I__6933 (
            .O(N__33869),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__6932 (
            .O(N__33866),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__6931 (
            .O(N__33863),
            .I(N__33860));
    LocalMux I__6930 (
            .O(N__33860),
            .I(N__33857));
    Odrv4 I__6929 (
            .O(N__33857),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__6928 (
            .O(N__33854),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__6927 (
            .O(N__33851),
            .I(N__33848));
    LocalMux I__6926 (
            .O(N__33848),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__6925 (
            .O(N__33845),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__6924 (
            .O(N__33842),
            .I(N__33838));
    CascadeMux I__6923 (
            .O(N__33841),
            .I(N__33835));
    LocalMux I__6922 (
            .O(N__33838),
            .I(N__33832));
    InMux I__6921 (
            .O(N__33835),
            .I(N__33829));
    Span4Mux_h I__6920 (
            .O(N__33832),
            .I(N__33826));
    LocalMux I__6919 (
            .O(N__33829),
            .I(N__33822));
    Span4Mux_v I__6918 (
            .O(N__33826),
            .I(N__33819));
    InMux I__6917 (
            .O(N__33825),
            .I(N__33816));
    Span4Mux_v I__6916 (
            .O(N__33822),
            .I(N__33813));
    Odrv4 I__6915 (
            .O(N__33819),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__6914 (
            .O(N__33816),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__6913 (
            .O(N__33813),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__6912 (
            .O(N__33806),
            .I(N__33803));
    LocalMux I__6911 (
            .O(N__33803),
            .I(N__33800));
    Span4Mux_h I__6910 (
            .O(N__33800),
            .I(N__33795));
    InMux I__6909 (
            .O(N__33799),
            .I(N__33790));
    InMux I__6908 (
            .O(N__33798),
            .I(N__33790));
    Odrv4 I__6907 (
            .O(N__33795),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__6906 (
            .O(N__33790),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    InMux I__6905 (
            .O(N__33785),
            .I(N__33782));
    LocalMux I__6904 (
            .O(N__33782),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    InMux I__6903 (
            .O(N__33779),
            .I(N__33774));
    CascadeMux I__6902 (
            .O(N__33778),
            .I(N__33771));
    InMux I__6901 (
            .O(N__33777),
            .I(N__33768));
    LocalMux I__6900 (
            .O(N__33774),
            .I(N__33765));
    InMux I__6899 (
            .O(N__33771),
            .I(N__33762));
    LocalMux I__6898 (
            .O(N__33768),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv4 I__6897 (
            .O(N__33765),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__6896 (
            .O(N__33762),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__6895 (
            .O(N__33755),
            .I(N__33751));
    CascadeMux I__6894 (
            .O(N__33754),
            .I(N__33748));
    LocalMux I__6893 (
            .O(N__33751),
            .I(N__33745));
    InMux I__6892 (
            .O(N__33748),
            .I(N__33742));
    Odrv12 I__6891 (
            .O(N__33745),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__6890 (
            .O(N__33742),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__6889 (
            .O(N__33737),
            .I(N__33734));
    LocalMux I__6888 (
            .O(N__33734),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__6887 (
            .O(N__33731),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__6886 (
            .O(N__33728),
            .I(N__33725));
    LocalMux I__6885 (
            .O(N__33725),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__6884 (
            .O(N__33722),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__6883 (
            .O(N__33719),
            .I(N__33716));
    LocalMux I__6882 (
            .O(N__33716),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__6881 (
            .O(N__33713),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__6880 (
            .O(N__33710),
            .I(N__33707));
    LocalMux I__6879 (
            .O(N__33707),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__6878 (
            .O(N__33704),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    CascadeMux I__6877 (
            .O(N__33701),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_ ));
    InMux I__6876 (
            .O(N__33698),
            .I(N__33695));
    LocalMux I__6875 (
            .O(N__33695),
            .I(N__33692));
    Span4Mux_v I__6874 (
            .O(N__33692),
            .I(N__33687));
    InMux I__6873 (
            .O(N__33691),
            .I(N__33684));
    InMux I__6872 (
            .O(N__33690),
            .I(N__33681));
    Odrv4 I__6871 (
            .O(N__33687),
            .I(elapsed_time_ns_1_RNIPFL2M1_0_1));
    LocalMux I__6870 (
            .O(N__33684),
            .I(elapsed_time_ns_1_RNIPFL2M1_0_1));
    LocalMux I__6869 (
            .O(N__33681),
            .I(elapsed_time_ns_1_RNIPFL2M1_0_1));
    CascadeMux I__6868 (
            .O(N__33674),
            .I(elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_));
    InMux I__6867 (
            .O(N__33671),
            .I(N__33668));
    LocalMux I__6866 (
            .O(N__33668),
            .I(N__33665));
    Span4Mux_v I__6865 (
            .O(N__33665),
            .I(N__33661));
    InMux I__6864 (
            .O(N__33664),
            .I(N__33658));
    Odrv4 I__6863 (
            .O(N__33661),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_0_1Z0Z_1 ));
    LocalMux I__6862 (
            .O(N__33658),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_0_1Z0Z_1 ));
    CascadeMux I__6861 (
            .O(N__33653),
            .I(elapsed_time_ns_1_RNISCJF91_0_31_cascade_));
    InMux I__6860 (
            .O(N__33650),
            .I(N__33646));
    CascadeMux I__6859 (
            .O(N__33649),
            .I(N__33643));
    LocalMux I__6858 (
            .O(N__33646),
            .I(N__33640));
    InMux I__6857 (
            .O(N__33643),
            .I(N__33637));
    Span4Mux_h I__6856 (
            .O(N__33640),
            .I(N__33634));
    LocalMux I__6855 (
            .O(N__33637),
            .I(N__33630));
    Span4Mux_v I__6854 (
            .O(N__33634),
            .I(N__33627));
    InMux I__6853 (
            .O(N__33633),
            .I(N__33624));
    Span4Mux_v I__6852 (
            .O(N__33630),
            .I(N__33621));
    Odrv4 I__6851 (
            .O(N__33627),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__6850 (
            .O(N__33624),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__6849 (
            .O(N__33621),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__6848 (
            .O(N__33614),
            .I(N__33609));
    InMux I__6847 (
            .O(N__33613),
            .I(N__33604));
    InMux I__6846 (
            .O(N__33612),
            .I(N__33604));
    LocalMux I__6845 (
            .O(N__33609),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6844 (
            .O(N__33604),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__6843 (
            .O(N__33599),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_ ));
    InMux I__6842 (
            .O(N__33596),
            .I(N__33593));
    LocalMux I__6841 (
            .O(N__33593),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    CascadeMux I__6840 (
            .O(N__33590),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15_cascade_));
    CascadeMux I__6839 (
            .O(N__33587),
            .I(\phase_controller_inst1.stoper_tr.N_251_cascade_ ));
    CascadeMux I__6838 (
            .O(N__33584),
            .I(elapsed_time_ns_1_RNIDH2591_0_5_cascade_));
    InMux I__6837 (
            .O(N__33581),
            .I(N__33578));
    LocalMux I__6836 (
            .O(N__33578),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3Z0Z_2 ));
    CascadeMux I__6835 (
            .O(N__33575),
            .I(\phase_controller_inst1.stoper_tr.N_241_cascade_ ));
    InMux I__6834 (
            .O(N__33572),
            .I(N__33569));
    LocalMux I__6833 (
            .O(N__33569),
            .I(N__33566));
    Odrv12 I__6832 (
            .O(N__33566),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ));
    InMux I__6831 (
            .O(N__33563),
            .I(N__33560));
    LocalMux I__6830 (
            .O(N__33560),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ));
    InMux I__6829 (
            .O(N__33557),
            .I(N__33554));
    LocalMux I__6828 (
            .O(N__33554),
            .I(\delay_measurement_inst.delay_tr_timer.N_381 ));
    InMux I__6827 (
            .O(N__33551),
            .I(N__33547));
    InMux I__6826 (
            .O(N__33550),
            .I(N__33544));
    LocalMux I__6825 (
            .O(N__33547),
            .I(\delay_measurement_inst.delay_tr_timer.N_359_1 ));
    LocalMux I__6824 (
            .O(N__33544),
            .I(\delay_measurement_inst.delay_tr_timer.N_359_1 ));
    CascadeMux I__6823 (
            .O(N__33539),
            .I(\delay_measurement_inst.delay_tr_timer.N_381_cascade_ ));
    CascadeMux I__6822 (
            .O(N__33536),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ));
    CascadeMux I__6821 (
            .O(N__33533),
            .I(elapsed_time_ns_1_RNISAHF91_0_13_cascade_));
    CascadeMux I__6820 (
            .O(N__33530),
            .I(N__33527));
    InMux I__6819 (
            .O(N__33527),
            .I(N__33523));
    InMux I__6818 (
            .O(N__33526),
            .I(N__33520));
    LocalMux I__6817 (
            .O(N__33523),
            .I(N__33517));
    LocalMux I__6816 (
            .O(N__33520),
            .I(N__33511));
    Span4Mux_v I__6815 (
            .O(N__33517),
            .I(N__33511));
    InMux I__6814 (
            .O(N__33516),
            .I(N__33508));
    Odrv4 I__6813 (
            .O(N__33511),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    LocalMux I__6812 (
            .O(N__33508),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    InMux I__6811 (
            .O(N__33503),
            .I(N__33500));
    LocalMux I__6810 (
            .O(N__33500),
            .I(N__33497));
    Span4Mux_v I__6809 (
            .O(N__33497),
            .I(N__33494));
    Odrv4 I__6808 (
            .O(N__33494),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ));
    CascadeMux I__6807 (
            .O(N__33491),
            .I(N__33488));
    InMux I__6806 (
            .O(N__33488),
            .I(N__33485));
    LocalMux I__6805 (
            .O(N__33485),
            .I(N__33482));
    Odrv4 I__6804 (
            .O(N__33482),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ));
    CascadeMux I__6803 (
            .O(N__33479),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_ ));
    CascadeMux I__6802 (
            .O(N__33476),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ));
    InMux I__6801 (
            .O(N__33473),
            .I(N__33470));
    LocalMux I__6800 (
            .O(N__33470),
            .I(elapsed_time_ns_1_RNI3JIF91_0_29));
    CascadeMux I__6799 (
            .O(N__33467),
            .I(N__33464));
    InMux I__6798 (
            .O(N__33464),
            .I(N__33460));
    InMux I__6797 (
            .O(N__33463),
            .I(N__33457));
    LocalMux I__6796 (
            .O(N__33460),
            .I(elapsed_time_ns_1_RNIRBJF91_0_30));
    LocalMux I__6795 (
            .O(N__33457),
            .I(elapsed_time_ns_1_RNIRBJF91_0_30));
    InMux I__6794 (
            .O(N__33452),
            .I(N__33446));
    InMux I__6793 (
            .O(N__33451),
            .I(N__33446));
    LocalMux I__6792 (
            .O(N__33446),
            .I(elapsed_time_ns_1_RNIRAIF91_0_21));
    CascadeMux I__6791 (
            .O(N__33443),
            .I(elapsed_time_ns_1_RNI3JIF91_0_29_cascade_));
    InMux I__6790 (
            .O(N__33440),
            .I(N__33436));
    InMux I__6789 (
            .O(N__33439),
            .I(N__33433));
    LocalMux I__6788 (
            .O(N__33436),
            .I(elapsed_time_ns_1_RNIQ9IF91_0_20));
    LocalMux I__6787 (
            .O(N__33433),
            .I(elapsed_time_ns_1_RNIQ9IF91_0_20));
    InMux I__6786 (
            .O(N__33428),
            .I(N__33422));
    InMux I__6785 (
            .O(N__33427),
            .I(N__33422));
    LocalMux I__6784 (
            .O(N__33422),
            .I(N__33419));
    Odrv4 I__6783 (
            .O(N__33419),
            .I(elapsed_time_ns_1_RNISBIF91_0_22));
    CascadeMux I__6782 (
            .O(N__33416),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_o5_7Z0Z_15_cascade_ ));
    InMux I__6781 (
            .O(N__33413),
            .I(N__33410));
    LocalMux I__6780 (
            .O(N__33410),
            .I(N__33407));
    Span4Mux_h I__6779 (
            .O(N__33407),
            .I(N__33404));
    Span4Mux_v I__6778 (
            .O(N__33404),
            .I(N__33401));
    Odrv4 I__6777 (
            .O(N__33401),
            .I(\current_shift_inst.PI_CTRL.integrator_i_27 ));
    CascadeMux I__6776 (
            .O(N__33398),
            .I(N__33395));
    InMux I__6775 (
            .O(N__33395),
            .I(N__33392));
    LocalMux I__6774 (
            .O(N__33392),
            .I(N__33389));
    Span4Mux_h I__6773 (
            .O(N__33389),
            .I(N__33386));
    Span4Mux_v I__6772 (
            .O(N__33386),
            .I(N__33383));
    Odrv4 I__6771 (
            .O(N__33383),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ));
    InMux I__6770 (
            .O(N__33380),
            .I(N__33377));
    LocalMux I__6769 (
            .O(N__33377),
            .I(N__33374));
    Span4Mux_h I__6768 (
            .O(N__33374),
            .I(N__33371));
    Odrv4 I__6767 (
            .O(N__33371),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__6766 (
            .O(N__33368),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ));
    CascadeMux I__6765 (
            .O(N__33365),
            .I(N__33362));
    InMux I__6764 (
            .O(N__33362),
            .I(N__33359));
    LocalMux I__6763 (
            .O(N__33359),
            .I(N__33356));
    Span12Mux_v I__6762 (
            .O(N__33356),
            .I(N__33353));
    Odrv12 I__6761 (
            .O(N__33353),
            .I(\current_shift_inst.PI_CTRL.integrator_i_28 ));
    InMux I__6760 (
            .O(N__33350),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ));
    CascadeMux I__6759 (
            .O(N__33347),
            .I(N__33344));
    InMux I__6758 (
            .O(N__33344),
            .I(N__33341));
    LocalMux I__6757 (
            .O(N__33341),
            .I(N__33338));
    Odrv12 I__6756 (
            .O(N__33338),
            .I(\current_shift_inst.PI_CTRL.integrator_i_29 ));
    InMux I__6755 (
            .O(N__33335),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ));
    InMux I__6754 (
            .O(N__33332),
            .I(N__33327));
    InMux I__6753 (
            .O(N__33331),
            .I(N__33322));
    InMux I__6752 (
            .O(N__33330),
            .I(N__33322));
    LocalMux I__6751 (
            .O(N__33327),
            .I(N__33317));
    LocalMux I__6750 (
            .O(N__33322),
            .I(N__33317));
    Span4Mux_h I__6749 (
            .O(N__33317),
            .I(N__33314));
    Odrv4 I__6748 (
            .O(N__33314),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_0_12 ));
    CascadeMux I__6747 (
            .O(N__33311),
            .I(N__33308));
    InMux I__6746 (
            .O(N__33308),
            .I(N__33305));
    LocalMux I__6745 (
            .O(N__33305),
            .I(N__33302));
    Span4Mux_v I__6744 (
            .O(N__33302),
            .I(N__33299));
    Span4Mux_v I__6743 (
            .O(N__33299),
            .I(N__33296));
    Odrv4 I__6742 (
            .O(N__33296),
            .I(\current_shift_inst.PI_CTRL.integrator_i_30 ));
    InMux I__6741 (
            .O(N__33293),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ));
    InMux I__6740 (
            .O(N__33290),
            .I(bfn_15_11_0_));
    InMux I__6739 (
            .O(N__33287),
            .I(N__33284));
    LocalMux I__6738 (
            .O(N__33284),
            .I(N__33281));
    Odrv4 I__6737 (
            .O(N__33281),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6 ));
    CascadeMux I__6736 (
            .O(N__33278),
            .I(\delay_measurement_inst.delay_tr_timer.N_363_cascade_ ));
    InMux I__6735 (
            .O(N__33275),
            .I(N__33272));
    LocalMux I__6734 (
            .O(N__33272),
            .I(N__33269));
    Span4Mux_v I__6733 (
            .O(N__33269),
            .I(N__33265));
    InMux I__6732 (
            .O(N__33268),
            .I(N__33261));
    Span4Mux_h I__6731 (
            .O(N__33265),
            .I(N__33258));
    InMux I__6730 (
            .O(N__33264),
            .I(N__33255));
    LocalMux I__6729 (
            .O(N__33261),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    Odrv4 I__6728 (
            .O(N__33258),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    LocalMux I__6727 (
            .O(N__33255),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    CascadeMux I__6726 (
            .O(N__33248),
            .I(N__33245));
    InMux I__6725 (
            .O(N__33245),
            .I(N__33242));
    LocalMux I__6724 (
            .O(N__33242),
            .I(N__33239));
    Span4Mux_h I__6723 (
            .O(N__33239),
            .I(N__33236));
    Odrv4 I__6722 (
            .O(N__33236),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ));
    InMux I__6721 (
            .O(N__33233),
            .I(N__33230));
    LocalMux I__6720 (
            .O(N__33230),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ));
    InMux I__6719 (
            .O(N__33227),
            .I(N__33224));
    LocalMux I__6718 (
            .O(N__33224),
            .I(N__33221));
    Odrv4 I__6717 (
            .O(N__33221),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__6716 (
            .O(N__33218),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ));
    InMux I__6715 (
            .O(N__33215),
            .I(N__33212));
    LocalMux I__6714 (
            .O(N__33212),
            .I(N__33209));
    Span4Mux_v I__6713 (
            .O(N__33209),
            .I(N__33206));
    Span4Mux_v I__6712 (
            .O(N__33206),
            .I(N__33203));
    Odrv4 I__6711 (
            .O(N__33203),
            .I(\current_shift_inst.PI_CTRL.integrator_i_20 ));
    CascadeMux I__6710 (
            .O(N__33200),
            .I(N__33197));
    InMux I__6709 (
            .O(N__33197),
            .I(N__33194));
    LocalMux I__6708 (
            .O(N__33194),
            .I(N__33191));
    Odrv4 I__6707 (
            .O(N__33191),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ));
    CascadeMux I__6706 (
            .O(N__33188),
            .I(N__33185));
    InMux I__6705 (
            .O(N__33185),
            .I(N__33182));
    LocalMux I__6704 (
            .O(N__33182),
            .I(N__33179));
    Odrv12 I__6703 (
            .O(N__33179),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__6702 (
            .O(N__33176),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ));
    InMux I__6701 (
            .O(N__33173),
            .I(N__33170));
    LocalMux I__6700 (
            .O(N__33170),
            .I(N__33167));
    Span4Mux_v I__6699 (
            .O(N__33167),
            .I(N__33164));
    Odrv4 I__6698 (
            .O(N__33164),
            .I(\current_shift_inst.PI_CTRL.integrator_i_21 ));
    CascadeMux I__6697 (
            .O(N__33161),
            .I(N__33158));
    InMux I__6696 (
            .O(N__33158),
            .I(N__33155));
    LocalMux I__6695 (
            .O(N__33155),
            .I(N__33152));
    Span4Mux_h I__6694 (
            .O(N__33152),
            .I(N__33149));
    Odrv4 I__6693 (
            .O(N__33149),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ));
    InMux I__6692 (
            .O(N__33146),
            .I(N__33143));
    LocalMux I__6691 (
            .O(N__33143),
            .I(N__33140));
    Odrv12 I__6690 (
            .O(N__33140),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__6689 (
            .O(N__33137),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ));
    InMux I__6688 (
            .O(N__33134),
            .I(N__33131));
    LocalMux I__6687 (
            .O(N__33131),
            .I(N__33128));
    Span4Mux_v I__6686 (
            .O(N__33128),
            .I(N__33125));
    Odrv4 I__6685 (
            .O(N__33125),
            .I(\current_shift_inst.PI_CTRL.integrator_i_22 ));
    CascadeMux I__6684 (
            .O(N__33122),
            .I(N__33119));
    InMux I__6683 (
            .O(N__33119),
            .I(N__33116));
    LocalMux I__6682 (
            .O(N__33116),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ));
    CascadeMux I__6681 (
            .O(N__33113),
            .I(N__33110));
    InMux I__6680 (
            .O(N__33110),
            .I(N__33107));
    LocalMux I__6679 (
            .O(N__33107),
            .I(N__33104));
    Span4Mux_h I__6678 (
            .O(N__33104),
            .I(N__33101));
    Odrv4 I__6677 (
            .O(N__33101),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__6676 (
            .O(N__33098),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ));
    CascadeMux I__6675 (
            .O(N__33095),
            .I(N__33092));
    InMux I__6674 (
            .O(N__33092),
            .I(N__33089));
    LocalMux I__6673 (
            .O(N__33089),
            .I(\current_shift_inst.PI_CTRL.integrator_i_23 ));
    InMux I__6672 (
            .O(N__33086),
            .I(bfn_15_10_0_));
    CascadeMux I__6671 (
            .O(N__33083),
            .I(N__33080));
    InMux I__6670 (
            .O(N__33080),
            .I(N__33077));
    LocalMux I__6669 (
            .O(N__33077),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ));
    InMux I__6668 (
            .O(N__33074),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ));
    InMux I__6667 (
            .O(N__33071),
            .I(N__33068));
    LocalMux I__6666 (
            .O(N__33068),
            .I(N__33065));
    Span4Mux_v I__6665 (
            .O(N__33065),
            .I(N__33062));
    Odrv4 I__6664 (
            .O(N__33062),
            .I(\current_shift_inst.PI_CTRL.integrator_i_25 ));
    InMux I__6663 (
            .O(N__33059),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ));
    InMux I__6662 (
            .O(N__33056),
            .I(N__33053));
    LocalMux I__6661 (
            .O(N__33053),
            .I(\current_shift_inst.PI_CTRL.integrator_i_26 ));
    CascadeMux I__6660 (
            .O(N__33050),
            .I(N__33047));
    InMux I__6659 (
            .O(N__33047),
            .I(N__33044));
    LocalMux I__6658 (
            .O(N__33044),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ));
    InMux I__6657 (
            .O(N__33041),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ));
    InMux I__6656 (
            .O(N__33038),
            .I(N__33035));
    LocalMux I__6655 (
            .O(N__33035),
            .I(N__33032));
    Span4Mux_h I__6654 (
            .O(N__33032),
            .I(N__33029));
    Odrv4 I__6653 (
            .O(N__33029),
            .I(\current_shift_inst.PI_CTRL.integrator_i_12 ));
    CascadeMux I__6652 (
            .O(N__33026),
            .I(N__33023));
    InMux I__6651 (
            .O(N__33023),
            .I(N__33020));
    LocalMux I__6650 (
            .O(N__33020),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ));
    InMux I__6649 (
            .O(N__33017),
            .I(N__33014));
    LocalMux I__6648 (
            .O(N__33014),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__6647 (
            .O(N__33011),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ));
    InMux I__6646 (
            .O(N__33008),
            .I(N__33005));
    LocalMux I__6645 (
            .O(N__33005),
            .I(N__33002));
    Span12Mux_h I__6644 (
            .O(N__33002),
            .I(N__32999));
    Odrv12 I__6643 (
            .O(N__32999),
            .I(\current_shift_inst.PI_CTRL.integrator_i_13 ));
    CascadeMux I__6642 (
            .O(N__32996),
            .I(N__32993));
    InMux I__6641 (
            .O(N__32993),
            .I(N__32990));
    LocalMux I__6640 (
            .O(N__32990),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ));
    CascadeMux I__6639 (
            .O(N__32987),
            .I(N__32984));
    InMux I__6638 (
            .O(N__32984),
            .I(N__32981));
    LocalMux I__6637 (
            .O(N__32981),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__6636 (
            .O(N__32978),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ));
    CascadeMux I__6635 (
            .O(N__32975),
            .I(N__32972));
    InMux I__6634 (
            .O(N__32972),
            .I(N__32969));
    LocalMux I__6633 (
            .O(N__32969),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ));
    CascadeMux I__6632 (
            .O(N__32966),
            .I(N__32963));
    InMux I__6631 (
            .O(N__32963),
            .I(N__32960));
    LocalMux I__6630 (
            .O(N__32960),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__6629 (
            .O(N__32957),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ));
    InMux I__6628 (
            .O(N__32954),
            .I(N__32951));
    LocalMux I__6627 (
            .O(N__32951),
            .I(\current_shift_inst.PI_CTRL.integrator_i_15 ));
    CascadeMux I__6626 (
            .O(N__32948),
            .I(N__32945));
    InMux I__6625 (
            .O(N__32945),
            .I(N__32942));
    LocalMux I__6624 (
            .O(N__32942),
            .I(N__32939));
    Odrv12 I__6623 (
            .O(N__32939),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ));
    InMux I__6622 (
            .O(N__32936),
            .I(N__32933));
    LocalMux I__6621 (
            .O(N__32933),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__6620 (
            .O(N__32930),
            .I(bfn_15_9_0_));
    InMux I__6619 (
            .O(N__32927),
            .I(N__32924));
    LocalMux I__6618 (
            .O(N__32924),
            .I(N__32921));
    Span4Mux_h I__6617 (
            .O(N__32921),
            .I(N__32918));
    Odrv4 I__6616 (
            .O(N__32918),
            .I(\current_shift_inst.PI_CTRL.integrator_i_16 ));
    CascadeMux I__6615 (
            .O(N__32915),
            .I(N__32912));
    InMux I__6614 (
            .O(N__32912),
            .I(N__32909));
    LocalMux I__6613 (
            .O(N__32909),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ));
    InMux I__6612 (
            .O(N__32906),
            .I(N__32903));
    LocalMux I__6611 (
            .O(N__32903),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__6610 (
            .O(N__32900),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ));
    InMux I__6609 (
            .O(N__32897),
            .I(N__32894));
    LocalMux I__6608 (
            .O(N__32894),
            .I(N__32891));
    Span4Mux_h I__6607 (
            .O(N__32891),
            .I(N__32888));
    Odrv4 I__6606 (
            .O(N__32888),
            .I(\current_shift_inst.PI_CTRL.integrator_i_17 ));
    CascadeMux I__6605 (
            .O(N__32885),
            .I(N__32882));
    InMux I__6604 (
            .O(N__32882),
            .I(N__32879));
    LocalMux I__6603 (
            .O(N__32879),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ));
    InMux I__6602 (
            .O(N__32876),
            .I(N__32873));
    LocalMux I__6601 (
            .O(N__32873),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__6600 (
            .O(N__32870),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ));
    InMux I__6599 (
            .O(N__32867),
            .I(N__32864));
    LocalMux I__6598 (
            .O(N__32864),
            .I(N__32861));
    Odrv12 I__6597 (
            .O(N__32861),
            .I(\current_shift_inst.PI_CTRL.integrator_i_18 ));
    CascadeMux I__6596 (
            .O(N__32858),
            .I(N__32855));
    InMux I__6595 (
            .O(N__32855),
            .I(N__32852));
    LocalMux I__6594 (
            .O(N__32852),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ));
    InMux I__6593 (
            .O(N__32849),
            .I(N__32846));
    LocalMux I__6592 (
            .O(N__32846),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__6591 (
            .O(N__32843),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ));
    InMux I__6590 (
            .O(N__32840),
            .I(N__32837));
    LocalMux I__6589 (
            .O(N__32837),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ));
    CascadeMux I__6588 (
            .O(N__32834),
            .I(N__32831));
    InMux I__6587 (
            .O(N__32831),
            .I(N__32828));
    LocalMux I__6586 (
            .O(N__32828),
            .I(N__32825));
    Odrv4 I__6585 (
            .O(N__32825),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ));
    CascadeMux I__6584 (
            .O(N__32822),
            .I(N__32819));
    InMux I__6583 (
            .O(N__32819),
            .I(N__32816));
    LocalMux I__6582 (
            .O(N__32816),
            .I(N__32813));
    Odrv4 I__6581 (
            .O(N__32813),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__6580 (
            .O(N__32810),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ));
    InMux I__6579 (
            .O(N__32807),
            .I(N__32804));
    LocalMux I__6578 (
            .O(N__32804),
            .I(N__32801));
    Span4Mux_h I__6577 (
            .O(N__32801),
            .I(N__32798));
    Odrv4 I__6576 (
            .O(N__32798),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ));
    CascadeMux I__6575 (
            .O(N__32795),
            .I(N__32792));
    InMux I__6574 (
            .O(N__32792),
            .I(N__32789));
    LocalMux I__6573 (
            .O(N__32789),
            .I(N__32786));
    Span12Mux_v I__6572 (
            .O(N__32786),
            .I(N__32783));
    Odrv12 I__6571 (
            .O(N__32783),
            .I(\current_shift_inst.PI_CTRL.integrator_i_5 ));
    InMux I__6570 (
            .O(N__32780),
            .I(N__32777));
    LocalMux I__6569 (
            .O(N__32777),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__6568 (
            .O(N__32774),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ));
    InMux I__6567 (
            .O(N__32771),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ));
    InMux I__6566 (
            .O(N__32768),
            .I(N__32765));
    LocalMux I__6565 (
            .O(N__32765),
            .I(\current_shift_inst.PI_CTRL.integrator_i_7 ));
    CascadeMux I__6564 (
            .O(N__32762),
            .I(N__32759));
    InMux I__6563 (
            .O(N__32759),
            .I(N__32756));
    LocalMux I__6562 (
            .O(N__32756),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ));
    InMux I__6561 (
            .O(N__32753),
            .I(N__32750));
    LocalMux I__6560 (
            .O(N__32750),
            .I(N__32747));
    Odrv4 I__6559 (
            .O(N__32747),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__6558 (
            .O(N__32744),
            .I(bfn_15_8_0_));
    InMux I__6557 (
            .O(N__32741),
            .I(N__32738));
    LocalMux I__6556 (
            .O(N__32738),
            .I(N__32735));
    Odrv12 I__6555 (
            .O(N__32735),
            .I(\current_shift_inst.PI_CTRL.integrator_i_8 ));
    CascadeMux I__6554 (
            .O(N__32732),
            .I(N__32729));
    InMux I__6553 (
            .O(N__32729),
            .I(N__32726));
    LocalMux I__6552 (
            .O(N__32726),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ));
    CascadeMux I__6551 (
            .O(N__32723),
            .I(N__32720));
    InMux I__6550 (
            .O(N__32720),
            .I(N__32717));
    LocalMux I__6549 (
            .O(N__32717),
            .I(N__32714));
    Span4Mux_h I__6548 (
            .O(N__32714),
            .I(N__32711));
    Odrv4 I__6547 (
            .O(N__32711),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__6546 (
            .O(N__32708),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ));
    InMux I__6545 (
            .O(N__32705),
            .I(N__32702));
    LocalMux I__6544 (
            .O(N__32702),
            .I(N__32699));
    Odrv4 I__6543 (
            .O(N__32699),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ));
    CascadeMux I__6542 (
            .O(N__32696),
            .I(N__32693));
    InMux I__6541 (
            .O(N__32693),
            .I(N__32690));
    LocalMux I__6540 (
            .O(N__32690),
            .I(N__32687));
    Span12Mux_v I__6539 (
            .O(N__32687),
            .I(N__32684));
    Odrv12 I__6538 (
            .O(N__32684),
            .I(\current_shift_inst.PI_CTRL.integrator_i_9 ));
    InMux I__6537 (
            .O(N__32681),
            .I(N__32678));
    LocalMux I__6536 (
            .O(N__32678),
            .I(N__32675));
    Odrv4 I__6535 (
            .O(N__32675),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__6534 (
            .O(N__32672),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ));
    CascadeMux I__6533 (
            .O(N__32669),
            .I(N__32666));
    InMux I__6532 (
            .O(N__32666),
            .I(N__32663));
    LocalMux I__6531 (
            .O(N__32663),
            .I(N__32660));
    Span4Mux_h I__6530 (
            .O(N__32660),
            .I(N__32657));
    Odrv4 I__6529 (
            .O(N__32657),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ));
    InMux I__6528 (
            .O(N__32654),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ));
    InMux I__6527 (
            .O(N__32651),
            .I(N__32648));
    LocalMux I__6526 (
            .O(N__32648),
            .I(N__32645));
    Span4Mux_h I__6525 (
            .O(N__32645),
            .I(N__32642));
    Span4Mux_h I__6524 (
            .O(N__32642),
            .I(N__32639));
    Odrv4 I__6523 (
            .O(N__32639),
            .I(\current_shift_inst.PI_CTRL.integrator_i_11 ));
    CascadeMux I__6522 (
            .O(N__32636),
            .I(N__32633));
    InMux I__6521 (
            .O(N__32633),
            .I(N__32630));
    LocalMux I__6520 (
            .O(N__32630),
            .I(N__32627));
    Span4Mux_h I__6519 (
            .O(N__32627),
            .I(N__32624));
    Odrv4 I__6518 (
            .O(N__32624),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ));
    InMux I__6517 (
            .O(N__32621),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ));
    InMux I__6516 (
            .O(N__32618),
            .I(N__32614));
    CascadeMux I__6515 (
            .O(N__32617),
            .I(N__32609));
    LocalMux I__6514 (
            .O(N__32614),
            .I(N__32605));
    InMux I__6513 (
            .O(N__32613),
            .I(N__32602));
    InMux I__6512 (
            .O(N__32612),
            .I(N__32599));
    InMux I__6511 (
            .O(N__32609),
            .I(N__32596));
    InMux I__6510 (
            .O(N__32608),
            .I(N__32593));
    Span4Mux_h I__6509 (
            .O(N__32605),
            .I(N__32590));
    LocalMux I__6508 (
            .O(N__32602),
            .I(N__32587));
    LocalMux I__6507 (
            .O(N__32599),
            .I(N__32582));
    LocalMux I__6506 (
            .O(N__32596),
            .I(N__32582));
    LocalMux I__6505 (
            .O(N__32593),
            .I(N__32575));
    Span4Mux_h I__6504 (
            .O(N__32590),
            .I(N__32575));
    Span4Mux_v I__6503 (
            .O(N__32587),
            .I(N__32575));
    Span4Mux_h I__6502 (
            .O(N__32582),
            .I(N__32572));
    Span4Mux_v I__6501 (
            .O(N__32575),
            .I(N__32569));
    Odrv4 I__6500 (
            .O(N__32572),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__6499 (
            .O(N__32569),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__6498 (
            .O(N__32564),
            .I(N__32561));
    InMux I__6497 (
            .O(N__32561),
            .I(N__32558));
    LocalMux I__6496 (
            .O(N__32558),
            .I(N__32553));
    CascadeMux I__6495 (
            .O(N__32557),
            .I(N__32550));
    InMux I__6494 (
            .O(N__32556),
            .I(N__32546));
    Span4Mux_h I__6493 (
            .O(N__32553),
            .I(N__32543));
    InMux I__6492 (
            .O(N__32550),
            .I(N__32540));
    InMux I__6491 (
            .O(N__32549),
            .I(N__32537));
    LocalMux I__6490 (
            .O(N__32546),
            .I(N__32534));
    Span4Mux_v I__6489 (
            .O(N__32543),
            .I(N__32526));
    LocalMux I__6488 (
            .O(N__32540),
            .I(N__32526));
    LocalMux I__6487 (
            .O(N__32537),
            .I(N__32526));
    Span4Mux_v I__6486 (
            .O(N__32534),
            .I(N__32523));
    InMux I__6485 (
            .O(N__32533),
            .I(N__32520));
    Span4Mux_h I__6484 (
            .O(N__32526),
            .I(N__32517));
    Odrv4 I__6483 (
            .O(N__32523),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__6482 (
            .O(N__32520),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__6481 (
            .O(N__32517),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__6480 (
            .O(N__32510),
            .I(N__32504));
    InMux I__6479 (
            .O(N__32509),
            .I(N__32501));
    InMux I__6478 (
            .O(N__32508),
            .I(N__32498));
    InMux I__6477 (
            .O(N__32507),
            .I(N__32495));
    LocalMux I__6476 (
            .O(N__32504),
            .I(N__32492));
    LocalMux I__6475 (
            .O(N__32501),
            .I(N__32488));
    LocalMux I__6474 (
            .O(N__32498),
            .I(N__32483));
    LocalMux I__6473 (
            .O(N__32495),
            .I(N__32483));
    Span12Mux_h I__6472 (
            .O(N__32492),
            .I(N__32480));
    InMux I__6471 (
            .O(N__32491),
            .I(N__32477));
    Span4Mux_v I__6470 (
            .O(N__32488),
            .I(N__32472));
    Span4Mux_h I__6469 (
            .O(N__32483),
            .I(N__32472));
    Odrv12 I__6468 (
            .O(N__32480),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__6467 (
            .O(N__32477),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__6466 (
            .O(N__32472),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    CascadeMux I__6465 (
            .O(N__32465),
            .I(N__32462));
    InMux I__6464 (
            .O(N__32462),
            .I(N__32458));
    InMux I__6463 (
            .O(N__32461),
            .I(N__32455));
    LocalMux I__6462 (
            .O(N__32458),
            .I(N__32450));
    LocalMux I__6461 (
            .O(N__32455),
            .I(N__32450));
    Span4Mux_h I__6460 (
            .O(N__32450),
            .I(N__32447));
    Odrv4 I__6459 (
            .O(N__32447),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_12 ));
    InMux I__6458 (
            .O(N__32444),
            .I(N__32440));
    InMux I__6457 (
            .O(N__32443),
            .I(N__32437));
    LocalMux I__6456 (
            .O(N__32440),
            .I(N__32434));
    LocalMux I__6455 (
            .O(N__32437),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    Odrv4 I__6454 (
            .O(N__32434),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    CascadeMux I__6453 (
            .O(N__32429),
            .I(N__32426));
    InMux I__6452 (
            .O(N__32426),
            .I(N__32423));
    LocalMux I__6451 (
            .O(N__32423),
            .I(N__32420));
    Span4Mux_h I__6450 (
            .O(N__32420),
            .I(N__32417));
    Odrv4 I__6449 (
            .O(N__32417),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ));
    CascadeMux I__6448 (
            .O(N__32414),
            .I(N__32411));
    InMux I__6447 (
            .O(N__32411),
            .I(N__32408));
    LocalMux I__6446 (
            .O(N__32408),
            .I(N__32403));
    InMux I__6445 (
            .O(N__32407),
            .I(N__32400));
    InMux I__6444 (
            .O(N__32406),
            .I(N__32397));
    Span4Mux_v I__6443 (
            .O(N__32403),
            .I(N__32394));
    LocalMux I__6442 (
            .O(N__32400),
            .I(N__32391));
    LocalMux I__6441 (
            .O(N__32397),
            .I(N__32388));
    Span4Mux_h I__6440 (
            .O(N__32394),
            .I(N__32385));
    Span4Mux_h I__6439 (
            .O(N__32391),
            .I(N__32380));
    Span4Mux_v I__6438 (
            .O(N__32388),
            .I(N__32380));
    Odrv4 I__6437 (
            .O(N__32385),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    Odrv4 I__6436 (
            .O(N__32380),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    InMux I__6435 (
            .O(N__32375),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ));
    InMux I__6434 (
            .O(N__32372),
            .I(N__32369));
    LocalMux I__6433 (
            .O(N__32369),
            .I(N__32366));
    Span12Mux_s9_v I__6432 (
            .O(N__32366),
            .I(N__32363));
    Odrv12 I__6431 (
            .O(N__32363),
            .I(\current_shift_inst.PI_CTRL.integrator_i_1 ));
    CascadeMux I__6430 (
            .O(N__32360),
            .I(N__32357));
    InMux I__6429 (
            .O(N__32357),
            .I(N__32354));
    LocalMux I__6428 (
            .O(N__32354),
            .I(N__32351));
    Span4Mux_h I__6427 (
            .O(N__32351),
            .I(N__32348));
    Odrv4 I__6426 (
            .O(N__32348),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ));
    CascadeMux I__6425 (
            .O(N__32345),
            .I(N__32342));
    InMux I__6424 (
            .O(N__32342),
            .I(N__32339));
    LocalMux I__6423 (
            .O(N__32339),
            .I(N__32333));
    InMux I__6422 (
            .O(N__32338),
            .I(N__32328));
    InMux I__6421 (
            .O(N__32337),
            .I(N__32328));
    CascadeMux I__6420 (
            .O(N__32336),
            .I(N__32325));
    Span4Mux_v I__6419 (
            .O(N__32333),
            .I(N__32322));
    LocalMux I__6418 (
            .O(N__32328),
            .I(N__32319));
    InMux I__6417 (
            .O(N__32325),
            .I(N__32316));
    Span4Mux_h I__6416 (
            .O(N__32322),
            .I(N__32311));
    Span4Mux_v I__6415 (
            .O(N__32319),
            .I(N__32311));
    LocalMux I__6414 (
            .O(N__32316),
            .I(N__32308));
    Span4Mux_h I__6413 (
            .O(N__32311),
            .I(N__32305));
    Odrv12 I__6412 (
            .O(N__32308),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__6411 (
            .O(N__32305),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__6410 (
            .O(N__32300),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ));
    InMux I__6409 (
            .O(N__32297),
            .I(N__32294));
    LocalMux I__6408 (
            .O(N__32294),
            .I(N__32291));
    Span4Mux_h I__6407 (
            .O(N__32291),
            .I(N__32288));
    Odrv4 I__6406 (
            .O(N__32288),
            .I(\current_shift_inst.PI_CTRL.integrator_i_2 ));
    InMux I__6405 (
            .O(N__32285),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ));
    InMux I__6404 (
            .O(N__32282),
            .I(N__32279));
    LocalMux I__6403 (
            .O(N__32279),
            .I(N__32276));
    Span4Mux_h I__6402 (
            .O(N__32276),
            .I(N__32273));
    Odrv4 I__6401 (
            .O(N__32273),
            .I(\current_shift_inst.PI_CTRL.integrator_i_3 ));
    CascadeMux I__6400 (
            .O(N__32270),
            .I(N__32267));
    InMux I__6399 (
            .O(N__32267),
            .I(N__32264));
    LocalMux I__6398 (
            .O(N__32264),
            .I(N__32261));
    Span4Mux_h I__6397 (
            .O(N__32261),
            .I(N__32258));
    Odrv4 I__6396 (
            .O(N__32258),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ));
    CascadeMux I__6395 (
            .O(N__32255),
            .I(N__32252));
    InMux I__6394 (
            .O(N__32252),
            .I(N__32248));
    InMux I__6393 (
            .O(N__32251),
            .I(N__32242));
    LocalMux I__6392 (
            .O(N__32248),
            .I(N__32239));
    InMux I__6391 (
            .O(N__32247),
            .I(N__32236));
    InMux I__6390 (
            .O(N__32246),
            .I(N__32233));
    InMux I__6389 (
            .O(N__32245),
            .I(N__32230));
    LocalMux I__6388 (
            .O(N__32242),
            .I(N__32225));
    Span4Mux_h I__6387 (
            .O(N__32239),
            .I(N__32225));
    LocalMux I__6386 (
            .O(N__32236),
            .I(N__32220));
    LocalMux I__6385 (
            .O(N__32233),
            .I(N__32220));
    LocalMux I__6384 (
            .O(N__32230),
            .I(N__32217));
    Span4Mux_h I__6383 (
            .O(N__32225),
            .I(N__32214));
    Span4Mux_h I__6382 (
            .O(N__32220),
            .I(N__32211));
    Odrv12 I__6381 (
            .O(N__32217),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__6380 (
            .O(N__32214),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__6379 (
            .O(N__32211),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__6378 (
            .O(N__32204),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ));
    InMux I__6377 (
            .O(N__32201),
            .I(N__32198));
    LocalMux I__6376 (
            .O(N__32198),
            .I(N__32195));
    Odrv12 I__6375 (
            .O(N__32195),
            .I(\current_shift_inst.PI_CTRL.integrator_i_4 ));
    CascadeMux I__6374 (
            .O(N__32192),
            .I(N__32189));
    InMux I__6373 (
            .O(N__32189),
            .I(N__32186));
    LocalMux I__6372 (
            .O(N__32186),
            .I(N__32183));
    Odrv12 I__6371 (
            .O(N__32183),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__6370 (
            .O(N__32180),
            .I(N__32171));
    InMux I__6369 (
            .O(N__32179),
            .I(N__32171));
    InMux I__6368 (
            .O(N__32178),
            .I(N__32171));
    LocalMux I__6367 (
            .O(N__32171),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__6366 (
            .O(N__32168),
            .I(N__32165));
    LocalMux I__6365 (
            .O(N__32165),
            .I(N__32162));
    Odrv12 I__6364 (
            .O(N__32162),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3 ));
    CascadeMux I__6363 (
            .O(N__32159),
            .I(N__32156));
    InMux I__6362 (
            .O(N__32156),
            .I(N__32153));
    LocalMux I__6361 (
            .O(N__32153),
            .I(N__32150));
    Span4Mux_v I__6360 (
            .O(N__32150),
            .I(N__32147));
    Odrv4 I__6359 (
            .O(N__32147),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__6358 (
            .O(N__32144),
            .I(N__32141));
    LocalMux I__6357 (
            .O(N__32141),
            .I(N__32138));
    Odrv4 I__6356 (
            .O(N__32138),
            .I(\current_shift_inst.un38_control_input_cry_5_c_RNOZ0 ));
    InMux I__6355 (
            .O(N__32135),
            .I(N__32132));
    LocalMux I__6354 (
            .O(N__32132),
            .I(N__32129));
    Odrv4 I__6353 (
            .O(N__32129),
            .I(\current_shift_inst.un38_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__6352 (
            .O(N__32126),
            .I(N__32123));
    InMux I__6351 (
            .O(N__32123),
            .I(N__32120));
    LocalMux I__6350 (
            .O(N__32120),
            .I(N__32117));
    Span12Mux_h I__6349 (
            .O(N__32117),
            .I(N__32114));
    Odrv12 I__6348 (
            .O(N__32114),
            .I(\current_shift_inst.un38_control_input_cry_8_c_RNOZ0 ));
    CascadeMux I__6347 (
            .O(N__32111),
            .I(N__32108));
    InMux I__6346 (
            .O(N__32108),
            .I(N__32105));
    LocalMux I__6345 (
            .O(N__32105),
            .I(N__32102));
    Span4Mux_v I__6344 (
            .O(N__32102),
            .I(N__32099));
    Odrv4 I__6343 (
            .O(N__32099),
            .I(\current_shift_inst.un38_control_input_cry_10_c_RNOZ0 ));
    CascadeMux I__6342 (
            .O(N__32096),
            .I(N__32093));
    InMux I__6341 (
            .O(N__32093),
            .I(N__32090));
    LocalMux I__6340 (
            .O(N__32090),
            .I(N__32087));
    Span4Mux_h I__6339 (
            .O(N__32087),
            .I(N__32084));
    Odrv4 I__6338 (
            .O(N__32084),
            .I(\current_shift_inst.un38_control_input_cry_12_c_RNOZ0 ));
    InMux I__6337 (
            .O(N__32081),
            .I(N__32078));
    LocalMux I__6336 (
            .O(N__32078),
            .I(N__32075));
    Span4Mux_h I__6335 (
            .O(N__32075),
            .I(N__32072));
    Odrv4 I__6334 (
            .O(N__32072),
            .I(\current_shift_inst.un38_control_input_cry_15_c_RNOZ0 ));
    InMux I__6333 (
            .O(N__32069),
            .I(N__32066));
    LocalMux I__6332 (
            .O(N__32066),
            .I(N__32063));
    Span4Mux_h I__6331 (
            .O(N__32063),
            .I(N__32060));
    Odrv4 I__6330 (
            .O(N__32060),
            .I(\current_shift_inst.un38_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__6329 (
            .O(N__32057),
            .I(N__32051));
    InMux I__6328 (
            .O(N__32056),
            .I(N__32043));
    InMux I__6327 (
            .O(N__32055),
            .I(N__32043));
    InMux I__6326 (
            .O(N__32054),
            .I(N__32043));
    InMux I__6325 (
            .O(N__32051),
            .I(N__32038));
    InMux I__6324 (
            .O(N__32050),
            .I(N__32038));
    LocalMux I__6323 (
            .O(N__32043),
            .I(N__32035));
    LocalMux I__6322 (
            .O(N__32038),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__6321 (
            .O(N__32035),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__6320 (
            .O(N__32030),
            .I(N__32026));
    InMux I__6319 (
            .O(N__32029),
            .I(N__32016));
    InMux I__6318 (
            .O(N__32026),
            .I(N__32016));
    InMux I__6317 (
            .O(N__32025),
            .I(N__32016));
    InMux I__6316 (
            .O(N__32024),
            .I(N__32011));
    InMux I__6315 (
            .O(N__32023),
            .I(N__32011));
    LocalMux I__6314 (
            .O(N__32016),
            .I(N__32008));
    LocalMux I__6313 (
            .O(N__32011),
            .I(N__32004));
    Span4Mux_h I__6312 (
            .O(N__32008),
            .I(N__32001));
    InMux I__6311 (
            .O(N__32007),
            .I(N__31998));
    Span4Mux_v I__6310 (
            .O(N__32004),
            .I(N__31995));
    Span4Mux_v I__6309 (
            .O(N__32001),
            .I(N__31992));
    LocalMux I__6308 (
            .O(N__31998),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__6307 (
            .O(N__31995),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__6306 (
            .O(N__31992),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__6305 (
            .O(N__31985),
            .I(N__31982));
    LocalMux I__6304 (
            .O(N__31982),
            .I(N__31979));
    Span4Mux_v I__6303 (
            .O(N__31979),
            .I(N__31976));
    Span4Mux_h I__6302 (
            .O(N__31976),
            .I(N__31973));
    Odrv4 I__6301 (
            .O(N__31973),
            .I(\phase_controller_inst2.stoper_hc.N_45 ));
    InMux I__6300 (
            .O(N__31970),
            .I(N__31967));
    LocalMux I__6299 (
            .O(N__31967),
            .I(N__31964));
    Odrv4 I__6298 (
            .O(N__31964),
            .I(\phase_controller_inst1.stoper_tr.N_219 ));
    InMux I__6297 (
            .O(N__31961),
            .I(N__31958));
    LocalMux I__6296 (
            .O(N__31958),
            .I(N__31953));
    InMux I__6295 (
            .O(N__31957),
            .I(N__31950));
    InMux I__6294 (
            .O(N__31956),
            .I(N__31947));
    Span4Mux_v I__6293 (
            .O(N__31953),
            .I(N__31942));
    LocalMux I__6292 (
            .O(N__31950),
            .I(N__31942));
    LocalMux I__6291 (
            .O(N__31947),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    Odrv4 I__6290 (
            .O(N__31942),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    InMux I__6289 (
            .O(N__31937),
            .I(N__31933));
    InMux I__6288 (
            .O(N__31936),
            .I(N__31930));
    LocalMux I__6287 (
            .O(N__31933),
            .I(N__31926));
    LocalMux I__6286 (
            .O(N__31930),
            .I(N__31923));
    InMux I__6285 (
            .O(N__31929),
            .I(N__31920));
    Span4Mux_v I__6284 (
            .O(N__31926),
            .I(N__31915));
    Span4Mux_h I__6283 (
            .O(N__31923),
            .I(N__31915));
    LocalMux I__6282 (
            .O(N__31920),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    Odrv4 I__6281 (
            .O(N__31915),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    CascadeMux I__6280 (
            .O(N__31910),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    InMux I__6279 (
            .O(N__31907),
            .I(N__31904));
    LocalMux I__6278 (
            .O(N__31904),
            .I(N__31901));
    Span4Mux_h I__6277 (
            .O(N__31901),
            .I(N__31898));
    Odrv4 I__6276 (
            .O(N__31898),
            .I(\current_shift_inst.un38_control_input_cry_0_c_RNOZ0 ));
    InMux I__6275 (
            .O(N__31895),
            .I(N__31892));
    LocalMux I__6274 (
            .O(N__31892),
            .I(N__31889));
    Span4Mux_h I__6273 (
            .O(N__31889),
            .I(N__31886));
    Odrv4 I__6272 (
            .O(N__31886),
            .I(\current_shift_inst.un38_control_input_cry_6_c_RNOZ0 ));
    InMux I__6271 (
            .O(N__31883),
            .I(N__31880));
    LocalMux I__6270 (
            .O(N__31880),
            .I(N__31877));
    Span4Mux_h I__6269 (
            .O(N__31877),
            .I(N__31874));
    Odrv4 I__6268 (
            .O(N__31874),
            .I(\current_shift_inst.un38_control_input_cry_9_c_RNOZ0 ));
    CascadeMux I__6267 (
            .O(N__31871),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7_cascade_));
    CascadeMux I__6266 (
            .O(N__31868),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2_cascade_ ));
    InMux I__6265 (
            .O(N__31865),
            .I(N__31860));
    CascadeMux I__6264 (
            .O(N__31864),
            .I(N__31851));
    CascadeMux I__6263 (
            .O(N__31863),
            .I(N__31848));
    LocalMux I__6262 (
            .O(N__31860),
            .I(N__31844));
    InMux I__6261 (
            .O(N__31859),
            .I(N__31839));
    InMux I__6260 (
            .O(N__31858),
            .I(N__31839));
    InMux I__6259 (
            .O(N__31857),
            .I(N__31836));
    InMux I__6258 (
            .O(N__31856),
            .I(N__31830));
    InMux I__6257 (
            .O(N__31855),
            .I(N__31830));
    InMux I__6256 (
            .O(N__31854),
            .I(N__31827));
    InMux I__6255 (
            .O(N__31851),
            .I(N__31820));
    InMux I__6254 (
            .O(N__31848),
            .I(N__31820));
    InMux I__6253 (
            .O(N__31847),
            .I(N__31820));
    Span4Mux_v I__6252 (
            .O(N__31844),
            .I(N__31813));
    LocalMux I__6251 (
            .O(N__31839),
            .I(N__31810));
    LocalMux I__6250 (
            .O(N__31836),
            .I(N__31805));
    InMux I__6249 (
            .O(N__31835),
            .I(N__31796));
    LocalMux I__6248 (
            .O(N__31830),
            .I(N__31793));
    LocalMux I__6247 (
            .O(N__31827),
            .I(N__31788));
    LocalMux I__6246 (
            .O(N__31820),
            .I(N__31788));
    InMux I__6245 (
            .O(N__31819),
            .I(N__31779));
    InMux I__6244 (
            .O(N__31818),
            .I(N__31779));
    InMux I__6243 (
            .O(N__31817),
            .I(N__31779));
    InMux I__6242 (
            .O(N__31816),
            .I(N__31779));
    Sp12to4 I__6241 (
            .O(N__31813),
            .I(N__31768));
    Span4Mux_h I__6240 (
            .O(N__31810),
            .I(N__31765));
    InMux I__6239 (
            .O(N__31809),
            .I(N__31762));
    InMux I__6238 (
            .O(N__31808),
            .I(N__31759));
    Span12Mux_v I__6237 (
            .O(N__31805),
            .I(N__31756));
    InMux I__6236 (
            .O(N__31804),
            .I(N__31747));
    InMux I__6235 (
            .O(N__31803),
            .I(N__31747));
    InMux I__6234 (
            .O(N__31802),
            .I(N__31747));
    InMux I__6233 (
            .O(N__31801),
            .I(N__31747));
    InMux I__6232 (
            .O(N__31800),
            .I(N__31742));
    InMux I__6231 (
            .O(N__31799),
            .I(N__31742));
    LocalMux I__6230 (
            .O(N__31796),
            .I(N__31735));
    Span4Mux_v I__6229 (
            .O(N__31793),
            .I(N__31735));
    Span4Mux_v I__6228 (
            .O(N__31788),
            .I(N__31735));
    LocalMux I__6227 (
            .O(N__31779),
            .I(N__31732));
    InMux I__6226 (
            .O(N__31778),
            .I(N__31723));
    InMux I__6225 (
            .O(N__31777),
            .I(N__31723));
    InMux I__6224 (
            .O(N__31776),
            .I(N__31723));
    InMux I__6223 (
            .O(N__31775),
            .I(N__31723));
    InMux I__6222 (
            .O(N__31774),
            .I(N__31714));
    InMux I__6221 (
            .O(N__31773),
            .I(N__31714));
    InMux I__6220 (
            .O(N__31772),
            .I(N__31714));
    InMux I__6219 (
            .O(N__31771),
            .I(N__31714));
    Odrv12 I__6218 (
            .O(N__31768),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    Odrv4 I__6217 (
            .O(N__31765),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__6216 (
            .O(N__31762),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__6215 (
            .O(N__31759),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    Odrv12 I__6214 (
            .O(N__31756),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__6213 (
            .O(N__31747),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__6212 (
            .O(N__31742),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    Odrv4 I__6211 (
            .O(N__31735),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    Odrv4 I__6210 (
            .O(N__31732),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__6209 (
            .O(N__31723),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__6208 (
            .O(N__31714),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    InMux I__6207 (
            .O(N__31691),
            .I(N__31688));
    LocalMux I__6206 (
            .O(N__31688),
            .I(N__31684));
    CascadeMux I__6205 (
            .O(N__31687),
            .I(N__31680));
    Span4Mux_h I__6204 (
            .O(N__31684),
            .I(N__31676));
    InMux I__6203 (
            .O(N__31683),
            .I(N__31673));
    InMux I__6202 (
            .O(N__31680),
            .I(N__31670));
    InMux I__6201 (
            .O(N__31679),
            .I(N__31667));
    Odrv4 I__6200 (
            .O(N__31676),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6));
    LocalMux I__6199 (
            .O(N__31673),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6));
    LocalMux I__6198 (
            .O(N__31670),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6));
    LocalMux I__6197 (
            .O(N__31667),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6));
    CascadeMux I__6196 (
            .O(N__31658),
            .I(N__31654));
    CascadeMux I__6195 (
            .O(N__31657),
            .I(N__31651));
    InMux I__6194 (
            .O(N__31654),
            .I(N__31646));
    InMux I__6193 (
            .O(N__31651),
            .I(N__31642));
    CascadeMux I__6192 (
            .O(N__31650),
            .I(N__31639));
    CascadeMux I__6191 (
            .O(N__31649),
            .I(N__31634));
    LocalMux I__6190 (
            .O(N__31646),
            .I(N__31631));
    InMux I__6189 (
            .O(N__31645),
            .I(N__31628));
    LocalMux I__6188 (
            .O(N__31642),
            .I(N__31625));
    InMux I__6187 (
            .O(N__31639),
            .I(N__31622));
    InMux I__6186 (
            .O(N__31638),
            .I(N__31614));
    InMux I__6185 (
            .O(N__31637),
            .I(N__31614));
    InMux I__6184 (
            .O(N__31634),
            .I(N__31614));
    Sp12to4 I__6183 (
            .O(N__31631),
            .I(N__31609));
    LocalMux I__6182 (
            .O(N__31628),
            .I(N__31609));
    Span4Mux_h I__6181 (
            .O(N__31625),
            .I(N__31603));
    LocalMux I__6180 (
            .O(N__31622),
            .I(N__31603));
    InMux I__6179 (
            .O(N__31621),
            .I(N__31600));
    LocalMux I__6178 (
            .O(N__31614),
            .I(N__31597));
    Span12Mux_v I__6177 (
            .O(N__31609),
            .I(N__31594));
    InMux I__6176 (
            .O(N__31608),
            .I(N__31591));
    Span4Mux_h I__6175 (
            .O(N__31603),
            .I(N__31584));
    LocalMux I__6174 (
            .O(N__31600),
            .I(N__31584));
    Span4Mux_h I__6173 (
            .O(N__31597),
            .I(N__31584));
    Odrv12 I__6172 (
            .O(N__31594),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    LocalMux I__6171 (
            .O(N__31591),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    Odrv4 I__6170 (
            .O(N__31584),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    InMux I__6169 (
            .O(N__31577),
            .I(N__31574));
    LocalMux I__6168 (
            .O(N__31574),
            .I(N__31571));
    Span4Mux_h I__6167 (
            .O(N__31571),
            .I(N__31567));
    InMux I__6166 (
            .O(N__31570),
            .I(N__31563));
    Span4Mux_v I__6165 (
            .O(N__31567),
            .I(N__31560));
    InMux I__6164 (
            .O(N__31566),
            .I(N__31557));
    LocalMux I__6163 (
            .O(N__31563),
            .I(N__31554));
    Odrv4 I__6162 (
            .O(N__31560),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ));
    LocalMux I__6161 (
            .O(N__31557),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ));
    Odrv4 I__6160 (
            .O(N__31554),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ));
    InMux I__6159 (
            .O(N__31547),
            .I(N__31544));
    LocalMux I__6158 (
            .O(N__31544),
            .I(N__31541));
    Span4Mux_v I__6157 (
            .O(N__31541),
            .I(N__31538));
    Odrv4 I__6156 (
            .O(N__31538),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6 ));
    CascadeMux I__6155 (
            .O(N__31535),
            .I(\phase_controller_inst1.stoper_tr.N_235_cascade_ ));
    CascadeMux I__6154 (
            .O(N__31532),
            .I(\phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3_cascade_ ));
    CEMux I__6153 (
            .O(N__31529),
            .I(N__31523));
    CEMux I__6152 (
            .O(N__31528),
            .I(N__31519));
    CEMux I__6151 (
            .O(N__31527),
            .I(N__31516));
    CEMux I__6150 (
            .O(N__31526),
            .I(N__31513));
    LocalMux I__6149 (
            .O(N__31523),
            .I(N__31510));
    CEMux I__6148 (
            .O(N__31522),
            .I(N__31507));
    LocalMux I__6147 (
            .O(N__31519),
            .I(N__31504));
    LocalMux I__6146 (
            .O(N__31516),
            .I(N__31501));
    LocalMux I__6145 (
            .O(N__31513),
            .I(N__31498));
    Span4Mux_v I__6144 (
            .O(N__31510),
            .I(N__31493));
    LocalMux I__6143 (
            .O(N__31507),
            .I(N__31493));
    Span4Mux_h I__6142 (
            .O(N__31504),
            .I(N__31488));
    Span4Mux_h I__6141 (
            .O(N__31501),
            .I(N__31488));
    Span4Mux_h I__6140 (
            .O(N__31498),
            .I(N__31483));
    Span4Mux_h I__6139 (
            .O(N__31493),
            .I(N__31483));
    Span4Mux_h I__6138 (
            .O(N__31488),
            .I(N__31480));
    Span4Mux_h I__6137 (
            .O(N__31483),
            .I(N__31477));
    Odrv4 I__6136 (
            .O(N__31480),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa_0 ));
    Odrv4 I__6135 (
            .O(N__31477),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa_0 ));
    InMux I__6134 (
            .O(N__31472),
            .I(N__31467));
    CascadeMux I__6133 (
            .O(N__31471),
            .I(N__31464));
    InMux I__6132 (
            .O(N__31470),
            .I(N__31459));
    LocalMux I__6131 (
            .O(N__31467),
            .I(N__31453));
    InMux I__6130 (
            .O(N__31464),
            .I(N__31448));
    InMux I__6129 (
            .O(N__31463),
            .I(N__31448));
    InMux I__6128 (
            .O(N__31462),
            .I(N__31445));
    LocalMux I__6127 (
            .O(N__31459),
            .I(N__31442));
    InMux I__6126 (
            .O(N__31458),
            .I(N__31439));
    InMux I__6125 (
            .O(N__31457),
            .I(N__31434));
    InMux I__6124 (
            .O(N__31456),
            .I(N__31434));
    Span4Mux_v I__6123 (
            .O(N__31453),
            .I(N__31431));
    LocalMux I__6122 (
            .O(N__31448),
            .I(N__31428));
    LocalMux I__6121 (
            .O(N__31445),
            .I(N__31423));
    Span4Mux_h I__6120 (
            .O(N__31442),
            .I(N__31423));
    LocalMux I__6119 (
            .O(N__31439),
            .I(N__31420));
    LocalMux I__6118 (
            .O(N__31434),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__6117 (
            .O(N__31431),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__6116 (
            .O(N__31428),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__6115 (
            .O(N__31423),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__6114 (
            .O(N__31420),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    SRMux I__6113 (
            .O(N__31409),
            .I(N__31404));
    SRMux I__6112 (
            .O(N__31408),
            .I(N__31401));
    SRMux I__6111 (
            .O(N__31407),
            .I(N__31397));
    LocalMux I__6110 (
            .O(N__31404),
            .I(N__31394));
    LocalMux I__6109 (
            .O(N__31401),
            .I(N__31391));
    SRMux I__6108 (
            .O(N__31400),
            .I(N__31388));
    LocalMux I__6107 (
            .O(N__31397),
            .I(N__31385));
    Span4Mux_v I__6106 (
            .O(N__31394),
            .I(N__31378));
    Span4Mux_v I__6105 (
            .O(N__31391),
            .I(N__31378));
    LocalMux I__6104 (
            .O(N__31388),
            .I(N__31378));
    Span4Mux_h I__6103 (
            .O(N__31385),
            .I(N__31375));
    Sp12to4 I__6102 (
            .O(N__31378),
            .I(N__31372));
    Span4Mux_h I__6101 (
            .O(N__31375),
            .I(N__31369));
    Odrv12 I__6100 (
            .O(N__31372),
            .I(\phase_controller_inst2.stoper_hc.un1_stoper_state12_1_0_i ));
    Odrv4 I__6099 (
            .O(N__31369),
            .I(\phase_controller_inst2.stoper_hc.un1_stoper_state12_1_0_i ));
    CascadeMux I__6098 (
            .O(N__31364),
            .I(\delay_measurement_inst.delay_tr_timer.N_358_cascade_ ));
    CascadeMux I__6097 (
            .O(N__31361),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ));
    CascadeMux I__6096 (
            .O(N__31358),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9_cascade_ ));
    InMux I__6095 (
            .O(N__31355),
            .I(N__31352));
    LocalMux I__6094 (
            .O(N__31352),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ));
    InMux I__6093 (
            .O(N__31349),
            .I(N__31345));
    InMux I__6092 (
            .O(N__31348),
            .I(N__31342));
    LocalMux I__6091 (
            .O(N__31345),
            .I(N__31338));
    LocalMux I__6090 (
            .O(N__31342),
            .I(N__31335));
    InMux I__6089 (
            .O(N__31341),
            .I(N__31332));
    Span4Mux_h I__6088 (
            .O(N__31338),
            .I(N__31329));
    Span4Mux_v I__6087 (
            .O(N__31335),
            .I(N__31326));
    LocalMux I__6086 (
            .O(N__31332),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    Odrv4 I__6085 (
            .O(N__31329),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    Odrv4 I__6084 (
            .O(N__31326),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    InMux I__6083 (
            .O(N__31319),
            .I(N__31316));
    LocalMux I__6082 (
            .O(N__31316),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ));
    CascadeMux I__6081 (
            .O(N__31313),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_ ));
    CascadeMux I__6080 (
            .O(N__31310),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ));
    CascadeMux I__6079 (
            .O(N__31307),
            .I(N__31304));
    InMux I__6078 (
            .O(N__31304),
            .I(N__31300));
    InMux I__6077 (
            .O(N__31303),
            .I(N__31297));
    LocalMux I__6076 (
            .O(N__31300),
            .I(N__31294));
    LocalMux I__6075 (
            .O(N__31297),
            .I(N__31288));
    Span4Mux_v I__6074 (
            .O(N__31294),
            .I(N__31288));
    InMux I__6073 (
            .O(N__31293),
            .I(N__31285));
    Odrv4 I__6072 (
            .O(N__31288),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    LocalMux I__6071 (
            .O(N__31285),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    InMux I__6070 (
            .O(N__31280),
            .I(N__31277));
    LocalMux I__6069 (
            .O(N__31277),
            .I(N__31274));
    Span4Mux_v I__6068 (
            .O(N__31274),
            .I(N__31271));
    Odrv4 I__6067 (
            .O(N__31271),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ));
    InMux I__6066 (
            .O(N__31268),
            .I(N__31264));
    InMux I__6065 (
            .O(N__31267),
            .I(N__31260));
    LocalMux I__6064 (
            .O(N__31264),
            .I(N__31257));
    InMux I__6063 (
            .O(N__31263),
            .I(N__31254));
    LocalMux I__6062 (
            .O(N__31260),
            .I(N__31250));
    Span4Mux_h I__6061 (
            .O(N__31257),
            .I(N__31245));
    LocalMux I__6060 (
            .O(N__31254),
            .I(N__31245));
    InMux I__6059 (
            .O(N__31253),
            .I(N__31242));
    Span4Mux_v I__6058 (
            .O(N__31250),
            .I(N__31234));
    Span4Mux_v I__6057 (
            .O(N__31245),
            .I(N__31234));
    LocalMux I__6056 (
            .O(N__31242),
            .I(N__31234));
    InMux I__6055 (
            .O(N__31241),
            .I(N__31231));
    Odrv4 I__6054 (
            .O(N__31234),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__6053 (
            .O(N__31231),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__6052 (
            .O(N__31226),
            .I(N__31222));
    InMux I__6051 (
            .O(N__31225),
            .I(N__31219));
    LocalMux I__6050 (
            .O(N__31222),
            .I(N__31216));
    LocalMux I__6049 (
            .O(N__31219),
            .I(N__31213));
    Span4Mux_v I__6048 (
            .O(N__31216),
            .I(N__31209));
    Span4Mux_h I__6047 (
            .O(N__31213),
            .I(N__31206));
    InMux I__6046 (
            .O(N__31212),
            .I(N__31203));
    Odrv4 I__6045 (
            .O(N__31209),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv4 I__6044 (
            .O(N__31206),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    LocalMux I__6043 (
            .O(N__31203),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__6042 (
            .O(N__31196),
            .I(N__31193));
    LocalMux I__6041 (
            .O(N__31193),
            .I(N__31190));
    Odrv4 I__6040 (
            .O(N__31190),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_9 ));
    InMux I__6039 (
            .O(N__31187),
            .I(N__31182));
    InMux I__6038 (
            .O(N__31186),
            .I(N__31179));
    InMux I__6037 (
            .O(N__31185),
            .I(N__31176));
    LocalMux I__6036 (
            .O(N__31182),
            .I(N__31173));
    LocalMux I__6035 (
            .O(N__31179),
            .I(N__31170));
    LocalMux I__6034 (
            .O(N__31176),
            .I(N__31163));
    Span4Mux_v I__6033 (
            .O(N__31173),
            .I(N__31163));
    Span4Mux_v I__6032 (
            .O(N__31170),
            .I(N__31163));
    Odrv4 I__6031 (
            .O(N__31163),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    InMux I__6030 (
            .O(N__31160),
            .I(N__31157));
    LocalMux I__6029 (
            .O(N__31157),
            .I(N__31154));
    Span4Mux_h I__6028 (
            .O(N__31154),
            .I(N__31151));
    Odrv4 I__6027 (
            .O(N__31151),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ));
    CascadeMux I__6026 (
            .O(N__31148),
            .I(N__31145));
    InMux I__6025 (
            .O(N__31145),
            .I(N__31142));
    LocalMux I__6024 (
            .O(N__31142),
            .I(N__31138));
    InMux I__6023 (
            .O(N__31141),
            .I(N__31134));
    Span4Mux_h I__6022 (
            .O(N__31138),
            .I(N__31131));
    InMux I__6021 (
            .O(N__31137),
            .I(N__31128));
    LocalMux I__6020 (
            .O(N__31134),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    Odrv4 I__6019 (
            .O(N__31131),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    LocalMux I__6018 (
            .O(N__31128),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    InMux I__6017 (
            .O(N__31121),
            .I(N__31118));
    LocalMux I__6016 (
            .O(N__31118),
            .I(N__31115));
    Odrv4 I__6015 (
            .O(N__31115),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ));
    InMux I__6014 (
            .O(N__31112),
            .I(N__31108));
    InMux I__6013 (
            .O(N__31111),
            .I(N__31105));
    LocalMux I__6012 (
            .O(N__31108),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    LocalMux I__6011 (
            .O(N__31105),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    CascadeMux I__6010 (
            .O(N__31100),
            .I(N__31097));
    InMux I__6009 (
            .O(N__31097),
            .I(N__31092));
    CascadeMux I__6008 (
            .O(N__31096),
            .I(N__31089));
    InMux I__6007 (
            .O(N__31095),
            .I(N__31086));
    LocalMux I__6006 (
            .O(N__31092),
            .I(N__31082));
    InMux I__6005 (
            .O(N__31089),
            .I(N__31079));
    LocalMux I__6004 (
            .O(N__31086),
            .I(N__31076));
    InMux I__6003 (
            .O(N__31085),
            .I(N__31073));
    Span4Mux_h I__6002 (
            .O(N__31082),
            .I(N__31070));
    LocalMux I__6001 (
            .O(N__31079),
            .I(N__31067));
    Span4Mux_v I__6000 (
            .O(N__31076),
            .I(N__31060));
    LocalMux I__5999 (
            .O(N__31073),
            .I(N__31060));
    Span4Mux_v I__5998 (
            .O(N__31070),
            .I(N__31060));
    Span4Mux_v I__5997 (
            .O(N__31067),
            .I(N__31056));
    Span4Mux_h I__5996 (
            .O(N__31060),
            .I(N__31053));
    InMux I__5995 (
            .O(N__31059),
            .I(N__31050));
    Odrv4 I__5994 (
            .O(N__31056),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__5993 (
            .O(N__31053),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__5992 (
            .O(N__31050),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    CascadeMux I__5991 (
            .O(N__31043),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13_cascade_ ));
    InMux I__5990 (
            .O(N__31040),
            .I(N__31037));
    LocalMux I__5989 (
            .O(N__31037),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ));
    InMux I__5988 (
            .O(N__31034),
            .I(N__31030));
    InMux I__5987 (
            .O(N__31033),
            .I(N__31027));
    LocalMux I__5986 (
            .O(N__31030),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    LocalMux I__5985 (
            .O(N__31027),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    CascadeMux I__5984 (
            .O(N__31022),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14_cascade_ ));
    InMux I__5983 (
            .O(N__31019),
            .I(N__31016));
    LocalMux I__5982 (
            .O(N__31016),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ));
    CascadeMux I__5981 (
            .O(N__31013),
            .I(N__31010));
    InMux I__5980 (
            .O(N__31010),
            .I(N__31006));
    CascadeMux I__5979 (
            .O(N__31009),
            .I(N__31003));
    LocalMux I__5978 (
            .O(N__31006),
            .I(N__30999));
    InMux I__5977 (
            .O(N__31003),
            .I(N__30996));
    InMux I__5976 (
            .O(N__31002),
            .I(N__30991));
    Span4Mux_h I__5975 (
            .O(N__30999),
            .I(N__30986));
    LocalMux I__5974 (
            .O(N__30996),
            .I(N__30986));
    InMux I__5973 (
            .O(N__30995),
            .I(N__30983));
    InMux I__5972 (
            .O(N__30994),
            .I(N__30980));
    LocalMux I__5971 (
            .O(N__30991),
            .I(N__30975));
    Span4Mux_v I__5970 (
            .O(N__30986),
            .I(N__30975));
    LocalMux I__5969 (
            .O(N__30983),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__5968 (
            .O(N__30980),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__5967 (
            .O(N__30975),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__5966 (
            .O(N__30968),
            .I(N__30963));
    InMux I__5965 (
            .O(N__30967),
            .I(N__30960));
    InMux I__5964 (
            .O(N__30966),
            .I(N__30957));
    LocalMux I__5963 (
            .O(N__30963),
            .I(N__30954));
    LocalMux I__5962 (
            .O(N__30960),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    LocalMux I__5961 (
            .O(N__30957),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv12 I__5960 (
            .O(N__30954),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    CascadeMux I__5959 (
            .O(N__30947),
            .I(N__30944));
    InMux I__5958 (
            .O(N__30944),
            .I(N__30941));
    LocalMux I__5957 (
            .O(N__30941),
            .I(N__30938));
    Span4Mux_h I__5956 (
            .O(N__30938),
            .I(N__30935));
    Span4Mux_v I__5955 (
            .O(N__30935),
            .I(N__30932));
    Odrv4 I__5954 (
            .O(N__30932),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ));
    InMux I__5953 (
            .O(N__30929),
            .I(N__30924));
    InMux I__5952 (
            .O(N__30928),
            .I(N__30921));
    InMux I__5951 (
            .O(N__30927),
            .I(N__30918));
    LocalMux I__5950 (
            .O(N__30924),
            .I(N__30915));
    LocalMux I__5949 (
            .O(N__30921),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    LocalMux I__5948 (
            .O(N__30918),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    Odrv4 I__5947 (
            .O(N__30915),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    InMux I__5946 (
            .O(N__30908),
            .I(N__30904));
    InMux I__5945 (
            .O(N__30907),
            .I(N__30901));
    LocalMux I__5944 (
            .O(N__30904),
            .I(N__30897));
    LocalMux I__5943 (
            .O(N__30901),
            .I(N__30894));
    InMux I__5942 (
            .O(N__30900),
            .I(N__30889));
    Span4Mux_v I__5941 (
            .O(N__30897),
            .I(N__30886));
    Span12Mux_h I__5940 (
            .O(N__30894),
            .I(N__30883));
    InMux I__5939 (
            .O(N__30893),
            .I(N__30880));
    InMux I__5938 (
            .O(N__30892),
            .I(N__30877));
    LocalMux I__5937 (
            .O(N__30889),
            .I(N__30872));
    Span4Mux_v I__5936 (
            .O(N__30886),
            .I(N__30872));
    Odrv12 I__5935 (
            .O(N__30883),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__5934 (
            .O(N__30880),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__5933 (
            .O(N__30877),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__5932 (
            .O(N__30872),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__5931 (
            .O(N__30863),
            .I(N__30860));
    LocalMux I__5930 (
            .O(N__30860),
            .I(N__30857));
    Span4Mux_h I__5929 (
            .O(N__30857),
            .I(N__30854));
    Odrv4 I__5928 (
            .O(N__30854),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ));
    CascadeMux I__5927 (
            .O(N__30851),
            .I(N__30848));
    InMux I__5926 (
            .O(N__30848),
            .I(N__30844));
    InMux I__5925 (
            .O(N__30847),
            .I(N__30841));
    LocalMux I__5924 (
            .O(N__30844),
            .I(N__30837));
    LocalMux I__5923 (
            .O(N__30841),
            .I(N__30834));
    InMux I__5922 (
            .O(N__30840),
            .I(N__30831));
    Span4Mux_v I__5921 (
            .O(N__30837),
            .I(N__30826));
    Span4Mux_v I__5920 (
            .O(N__30834),
            .I(N__30826));
    LocalMux I__5919 (
            .O(N__30831),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    Odrv4 I__5918 (
            .O(N__30826),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    InMux I__5917 (
            .O(N__30821),
            .I(N__30818));
    LocalMux I__5916 (
            .O(N__30818),
            .I(N__30815));
    Span4Mux_h I__5915 (
            .O(N__30815),
            .I(N__30812));
    Odrv4 I__5914 (
            .O(N__30812),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ));
    InMux I__5913 (
            .O(N__30809),
            .I(N__30805));
    InMux I__5912 (
            .O(N__30808),
            .I(N__30801));
    LocalMux I__5911 (
            .O(N__30805),
            .I(N__30798));
    InMux I__5910 (
            .O(N__30804),
            .I(N__30795));
    LocalMux I__5909 (
            .O(N__30801),
            .I(N__30792));
    Span12Mux_h I__5908 (
            .O(N__30798),
            .I(N__30787));
    LocalMux I__5907 (
            .O(N__30795),
            .I(N__30782));
    Span4Mux_h I__5906 (
            .O(N__30792),
            .I(N__30782));
    InMux I__5905 (
            .O(N__30791),
            .I(N__30777));
    InMux I__5904 (
            .O(N__30790),
            .I(N__30777));
    Odrv12 I__5903 (
            .O(N__30787),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__5902 (
            .O(N__30782),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__5901 (
            .O(N__30777),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__5900 (
            .O(N__30770),
            .I(N__30765));
    InMux I__5899 (
            .O(N__30769),
            .I(N__30762));
    InMux I__5898 (
            .O(N__30768),
            .I(N__30759));
    LocalMux I__5897 (
            .O(N__30765),
            .I(N__30756));
    LocalMux I__5896 (
            .O(N__30762),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    LocalMux I__5895 (
            .O(N__30759),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    Odrv4 I__5894 (
            .O(N__30756),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    InMux I__5893 (
            .O(N__30749),
            .I(N__30746));
    LocalMux I__5892 (
            .O(N__30746),
            .I(N__30743));
    Odrv4 I__5891 (
            .O(N__30743),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ));
    InMux I__5890 (
            .O(N__30740),
            .I(N__30735));
    InMux I__5889 (
            .O(N__30739),
            .I(N__30732));
    InMux I__5888 (
            .O(N__30738),
            .I(N__30729));
    LocalMux I__5887 (
            .O(N__30735),
            .I(N__30726));
    LocalMux I__5886 (
            .O(N__30732),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    LocalMux I__5885 (
            .O(N__30729),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    Odrv12 I__5884 (
            .O(N__30726),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    InMux I__5883 (
            .O(N__30719),
            .I(N__30716));
    LocalMux I__5882 (
            .O(N__30716),
            .I(N__30713));
    Span4Mux_h I__5881 (
            .O(N__30713),
            .I(N__30710));
    Odrv4 I__5880 (
            .O(N__30710),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ));
    InMux I__5879 (
            .O(N__30707),
            .I(N__30704));
    LocalMux I__5878 (
            .O(N__30704),
            .I(N__30699));
    InMux I__5877 (
            .O(N__30703),
            .I(N__30696));
    InMux I__5876 (
            .O(N__30702),
            .I(N__30693));
    Span4Mux_v I__5875 (
            .O(N__30699),
            .I(N__30690));
    LocalMux I__5874 (
            .O(N__30696),
            .I(N__30687));
    LocalMux I__5873 (
            .O(N__30693),
            .I(N__30682));
    Span4Mux_h I__5872 (
            .O(N__30690),
            .I(N__30679));
    Span4Mux_h I__5871 (
            .O(N__30687),
            .I(N__30676));
    InMux I__5870 (
            .O(N__30686),
            .I(N__30671));
    InMux I__5869 (
            .O(N__30685),
            .I(N__30671));
    Odrv4 I__5868 (
            .O(N__30682),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__5867 (
            .O(N__30679),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__5866 (
            .O(N__30676),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__5865 (
            .O(N__30671),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    CascadeMux I__5864 (
            .O(N__30662),
            .I(N__30659));
    InMux I__5863 (
            .O(N__30659),
            .I(N__30656));
    LocalMux I__5862 (
            .O(N__30656),
            .I(N__30653));
    Span4Mux_h I__5861 (
            .O(N__30653),
            .I(N__30650));
    Odrv4 I__5860 (
            .O(N__30650),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ));
    CascadeMux I__5859 (
            .O(N__30647),
            .I(N__30644));
    InMux I__5858 (
            .O(N__30644),
            .I(N__30640));
    InMux I__5857 (
            .O(N__30643),
            .I(N__30637));
    LocalMux I__5856 (
            .O(N__30640),
            .I(N__30634));
    LocalMux I__5855 (
            .O(N__30637),
            .I(N__30631));
    Span4Mux_v I__5854 (
            .O(N__30634),
            .I(N__30627));
    Span4Mux_h I__5853 (
            .O(N__30631),
            .I(N__30622));
    InMux I__5852 (
            .O(N__30630),
            .I(N__30619));
    Span4Mux_h I__5851 (
            .O(N__30627),
            .I(N__30616));
    InMux I__5850 (
            .O(N__30626),
            .I(N__30611));
    InMux I__5849 (
            .O(N__30625),
            .I(N__30611));
    Odrv4 I__5848 (
            .O(N__30622),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__5847 (
            .O(N__30619),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__5846 (
            .O(N__30616),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__5845 (
            .O(N__30611),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__5844 (
            .O(N__30602),
            .I(N__30599));
    LocalMux I__5843 (
            .O(N__30599),
            .I(N__30596));
    Span4Mux_h I__5842 (
            .O(N__30596),
            .I(N__30591));
    CascadeMux I__5841 (
            .O(N__30595),
            .I(N__30588));
    InMux I__5840 (
            .O(N__30594),
            .I(N__30585));
    Span4Mux_v I__5839 (
            .O(N__30591),
            .I(N__30582));
    InMux I__5838 (
            .O(N__30588),
            .I(N__30579));
    LocalMux I__5837 (
            .O(N__30585),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    Odrv4 I__5836 (
            .O(N__30582),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    LocalMux I__5835 (
            .O(N__30579),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    InMux I__5834 (
            .O(N__30572),
            .I(N__30569));
    LocalMux I__5833 (
            .O(N__30569),
            .I(N__30566));
    Span4Mux_v I__5832 (
            .O(N__30566),
            .I(N__30563));
    Odrv4 I__5831 (
            .O(N__30563),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ));
    InMux I__5830 (
            .O(N__30560),
            .I(N__30555));
    InMux I__5829 (
            .O(N__30559),
            .I(N__30552));
    InMux I__5828 (
            .O(N__30558),
            .I(N__30549));
    LocalMux I__5827 (
            .O(N__30555),
            .I(N__30546));
    LocalMux I__5826 (
            .O(N__30552),
            .I(N__30543));
    LocalMux I__5825 (
            .O(N__30549),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    Odrv4 I__5824 (
            .O(N__30546),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    Odrv12 I__5823 (
            .O(N__30543),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    CascadeMux I__5822 (
            .O(N__30536),
            .I(N__30533));
    InMux I__5821 (
            .O(N__30533),
            .I(N__30530));
    LocalMux I__5820 (
            .O(N__30530),
            .I(N__30525));
    InMux I__5819 (
            .O(N__30529),
            .I(N__30520));
    InMux I__5818 (
            .O(N__30528),
            .I(N__30517));
    Span4Mux_v I__5817 (
            .O(N__30525),
            .I(N__30514));
    CascadeMux I__5816 (
            .O(N__30524),
            .I(N__30511));
    CascadeMux I__5815 (
            .O(N__30523),
            .I(N__30508));
    LocalMux I__5814 (
            .O(N__30520),
            .I(N__30505));
    LocalMux I__5813 (
            .O(N__30517),
            .I(N__30502));
    Span4Mux_h I__5812 (
            .O(N__30514),
            .I(N__30499));
    InMux I__5811 (
            .O(N__30511),
            .I(N__30496));
    InMux I__5810 (
            .O(N__30508),
            .I(N__30493));
    Span4Mux_h I__5809 (
            .O(N__30505),
            .I(N__30490));
    Odrv12 I__5808 (
            .O(N__30502),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__5807 (
            .O(N__30499),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__5806 (
            .O(N__30496),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__5805 (
            .O(N__30493),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__5804 (
            .O(N__30490),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__5803 (
            .O(N__30479),
            .I(N__30476));
    InMux I__5802 (
            .O(N__30476),
            .I(N__30473));
    LocalMux I__5801 (
            .O(N__30473),
            .I(N__30470));
    Span4Mux_h I__5800 (
            .O(N__30470),
            .I(N__30467));
    Odrv4 I__5799 (
            .O(N__30467),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ));
    InMux I__5798 (
            .O(N__30464),
            .I(N__30459));
    InMux I__5797 (
            .O(N__30463),
            .I(N__30456));
    InMux I__5796 (
            .O(N__30462),
            .I(N__30453));
    LocalMux I__5795 (
            .O(N__30459),
            .I(N__30450));
    LocalMux I__5794 (
            .O(N__30456),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    LocalMux I__5793 (
            .O(N__30453),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    Odrv12 I__5792 (
            .O(N__30450),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    CascadeMux I__5791 (
            .O(N__30443),
            .I(N__30440));
    InMux I__5790 (
            .O(N__30440),
            .I(N__30436));
    InMux I__5789 (
            .O(N__30439),
            .I(N__30433));
    LocalMux I__5788 (
            .O(N__30436),
            .I(N__30429));
    LocalMux I__5787 (
            .O(N__30433),
            .I(N__30426));
    InMux I__5786 (
            .O(N__30432),
            .I(N__30423));
    Span4Mux_v I__5785 (
            .O(N__30429),
            .I(N__30418));
    Span4Mux_h I__5784 (
            .O(N__30426),
            .I(N__30413));
    LocalMux I__5783 (
            .O(N__30423),
            .I(N__30413));
    InMux I__5782 (
            .O(N__30422),
            .I(N__30410));
    InMux I__5781 (
            .O(N__30421),
            .I(N__30407));
    Span4Mux_h I__5780 (
            .O(N__30418),
            .I(N__30404));
    Span4Mux_h I__5779 (
            .O(N__30413),
            .I(N__30399));
    LocalMux I__5778 (
            .O(N__30410),
            .I(N__30399));
    LocalMux I__5777 (
            .O(N__30407),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__5776 (
            .O(N__30404),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__5775 (
            .O(N__30399),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__5774 (
            .O(N__30392),
            .I(N__30389));
    LocalMux I__5773 (
            .O(N__30389),
            .I(N__30386));
    Odrv4 I__5772 (
            .O(N__30386),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ));
    InMux I__5771 (
            .O(N__30383),
            .I(N__30379));
    InMux I__5770 (
            .O(N__30382),
            .I(N__30376));
    LocalMux I__5769 (
            .O(N__30379),
            .I(N__30373));
    LocalMux I__5768 (
            .O(N__30376),
            .I(N__30370));
    Span12Mux_h I__5767 (
            .O(N__30373),
            .I(N__30364));
    Span4Mux_h I__5766 (
            .O(N__30370),
            .I(N__30361));
    InMux I__5765 (
            .O(N__30369),
            .I(N__30358));
    InMux I__5764 (
            .O(N__30368),
            .I(N__30353));
    InMux I__5763 (
            .O(N__30367),
            .I(N__30353));
    Odrv12 I__5762 (
            .O(N__30364),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__5761 (
            .O(N__30361),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__5760 (
            .O(N__30358),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__5759 (
            .O(N__30353),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__5758 (
            .O(N__30344),
            .I(N__30341));
    InMux I__5757 (
            .O(N__30341),
            .I(N__30338));
    LocalMux I__5756 (
            .O(N__30338),
            .I(N__30335));
    Span4Mux_v I__5755 (
            .O(N__30335),
            .I(N__30331));
    InMux I__5754 (
            .O(N__30334),
            .I(N__30327));
    Span4Mux_v I__5753 (
            .O(N__30331),
            .I(N__30324));
    InMux I__5752 (
            .O(N__30330),
            .I(N__30321));
    LocalMux I__5751 (
            .O(N__30327),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv4 I__5750 (
            .O(N__30324),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    LocalMux I__5749 (
            .O(N__30321),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__5748 (
            .O(N__30314),
            .I(N__30311));
    LocalMux I__5747 (
            .O(N__30311),
            .I(N__30308));
    Span4Mux_v I__5746 (
            .O(N__30308),
            .I(N__30305));
    Odrv4 I__5745 (
            .O(N__30305),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_8 ));
    InMux I__5744 (
            .O(N__30302),
            .I(N__30298));
    InMux I__5743 (
            .O(N__30301),
            .I(N__30295));
    LocalMux I__5742 (
            .O(N__30298),
            .I(N__30291));
    LocalMux I__5741 (
            .O(N__30295),
            .I(N__30288));
    InMux I__5740 (
            .O(N__30294),
            .I(N__30283));
    Span12Mux_v I__5739 (
            .O(N__30291),
            .I(N__30280));
    Span4Mux_v I__5738 (
            .O(N__30288),
            .I(N__30277));
    InMux I__5737 (
            .O(N__30287),
            .I(N__30272));
    InMux I__5736 (
            .O(N__30286),
            .I(N__30272));
    LocalMux I__5735 (
            .O(N__30283),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv12 I__5734 (
            .O(N__30280),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__5733 (
            .O(N__30277),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__5732 (
            .O(N__30272),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__5731 (
            .O(N__30263),
            .I(N__30260));
    LocalMux I__5730 (
            .O(N__30260),
            .I(N__30257));
    Span4Mux_h I__5729 (
            .O(N__30257),
            .I(N__30254));
    Odrv4 I__5728 (
            .O(N__30254),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ));
    InMux I__5727 (
            .O(N__30251),
            .I(N__30246));
    InMux I__5726 (
            .O(N__30250),
            .I(N__30243));
    InMux I__5725 (
            .O(N__30249),
            .I(N__30240));
    LocalMux I__5724 (
            .O(N__30246),
            .I(N__30237));
    LocalMux I__5723 (
            .O(N__30243),
            .I(N__30234));
    LocalMux I__5722 (
            .O(N__30240),
            .I(N__30231));
    Span4Mux_h I__5721 (
            .O(N__30237),
            .I(N__30228));
    Span4Mux_v I__5720 (
            .O(N__30234),
            .I(N__30223));
    Span4Mux_v I__5719 (
            .O(N__30231),
            .I(N__30223));
    Odrv4 I__5718 (
            .O(N__30228),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv4 I__5717 (
            .O(N__30223),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__5716 (
            .O(N__30218),
            .I(N__30215));
    LocalMux I__5715 (
            .O(N__30215),
            .I(N__30212));
    Span4Mux_h I__5714 (
            .O(N__30212),
            .I(N__30209));
    Odrv4 I__5713 (
            .O(N__30209),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_11 ));
    CascadeMux I__5712 (
            .O(N__30206),
            .I(N__30203));
    InMux I__5711 (
            .O(N__30203),
            .I(N__30198));
    InMux I__5710 (
            .O(N__30202),
            .I(N__30195));
    InMux I__5709 (
            .O(N__30201),
            .I(N__30192));
    LocalMux I__5708 (
            .O(N__30198),
            .I(N__30187));
    LocalMux I__5707 (
            .O(N__30195),
            .I(N__30187));
    LocalMux I__5706 (
            .O(N__30192),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv12 I__5705 (
            .O(N__30187),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__5704 (
            .O(N__30182),
            .I(bfn_13_27_0_));
    CascadeMux I__5703 (
            .O(N__30179),
            .I(N__30176));
    InMux I__5702 (
            .O(N__30176),
            .I(N__30172));
    InMux I__5701 (
            .O(N__30175),
            .I(N__30169));
    LocalMux I__5700 (
            .O(N__30172),
            .I(N__30163));
    LocalMux I__5699 (
            .O(N__30169),
            .I(N__30163));
    InMux I__5698 (
            .O(N__30168),
            .I(N__30160));
    Span4Mux_v I__5697 (
            .O(N__30163),
            .I(N__30157));
    LocalMux I__5696 (
            .O(N__30160),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__5695 (
            .O(N__30157),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__5694 (
            .O(N__30152),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__5693 (
            .O(N__30149),
            .I(N__30143));
    InMux I__5692 (
            .O(N__30148),
            .I(N__30143));
    LocalMux I__5691 (
            .O(N__30143),
            .I(N__30139));
    InMux I__5690 (
            .O(N__30142),
            .I(N__30136));
    Span4Mux_v I__5689 (
            .O(N__30139),
            .I(N__30133));
    LocalMux I__5688 (
            .O(N__30136),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__5687 (
            .O(N__30133),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__5686 (
            .O(N__30128),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__5685 (
            .O(N__30125),
            .I(N__30118));
    InMux I__5684 (
            .O(N__30124),
            .I(N__30118));
    InMux I__5683 (
            .O(N__30123),
            .I(N__30115));
    LocalMux I__5682 (
            .O(N__30118),
            .I(N__30112));
    LocalMux I__5681 (
            .O(N__30115),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv12 I__5680 (
            .O(N__30112),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__5679 (
            .O(N__30107),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    CascadeMux I__5678 (
            .O(N__30104),
            .I(N__30101));
    InMux I__5677 (
            .O(N__30101),
            .I(N__30098));
    LocalMux I__5676 (
            .O(N__30098),
            .I(N__30094));
    InMux I__5675 (
            .O(N__30097),
            .I(N__30091));
    Span4Mux_v I__5674 (
            .O(N__30094),
            .I(N__30088));
    LocalMux I__5673 (
            .O(N__30091),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__5672 (
            .O(N__30088),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__5671 (
            .O(N__30083),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__5670 (
            .O(N__30080),
            .I(N__30060));
    InMux I__5669 (
            .O(N__30079),
            .I(N__30060));
    InMux I__5668 (
            .O(N__30078),
            .I(N__30060));
    InMux I__5667 (
            .O(N__30077),
            .I(N__30060));
    InMux I__5666 (
            .O(N__30076),
            .I(N__30033));
    InMux I__5665 (
            .O(N__30075),
            .I(N__30033));
    InMux I__5664 (
            .O(N__30074),
            .I(N__30033));
    InMux I__5663 (
            .O(N__30073),
            .I(N__30033));
    InMux I__5662 (
            .O(N__30072),
            .I(N__30024));
    InMux I__5661 (
            .O(N__30071),
            .I(N__30024));
    InMux I__5660 (
            .O(N__30070),
            .I(N__30024));
    InMux I__5659 (
            .O(N__30069),
            .I(N__30024));
    LocalMux I__5658 (
            .O(N__30060),
            .I(N__30021));
    InMux I__5657 (
            .O(N__30059),
            .I(N__30016));
    InMux I__5656 (
            .O(N__30058),
            .I(N__30016));
    InMux I__5655 (
            .O(N__30057),
            .I(N__30007));
    InMux I__5654 (
            .O(N__30056),
            .I(N__30007));
    InMux I__5653 (
            .O(N__30055),
            .I(N__30007));
    InMux I__5652 (
            .O(N__30054),
            .I(N__30007));
    InMux I__5651 (
            .O(N__30053),
            .I(N__29998));
    InMux I__5650 (
            .O(N__30052),
            .I(N__29998));
    InMux I__5649 (
            .O(N__30051),
            .I(N__29998));
    InMux I__5648 (
            .O(N__30050),
            .I(N__29998));
    InMux I__5647 (
            .O(N__30049),
            .I(N__29989));
    InMux I__5646 (
            .O(N__30048),
            .I(N__29989));
    InMux I__5645 (
            .O(N__30047),
            .I(N__29989));
    InMux I__5644 (
            .O(N__30046),
            .I(N__29989));
    InMux I__5643 (
            .O(N__30045),
            .I(N__29980));
    InMux I__5642 (
            .O(N__30044),
            .I(N__29980));
    InMux I__5641 (
            .O(N__30043),
            .I(N__29980));
    InMux I__5640 (
            .O(N__30042),
            .I(N__29980));
    LocalMux I__5639 (
            .O(N__30033),
            .I(N__29975));
    LocalMux I__5638 (
            .O(N__30024),
            .I(N__29975));
    Odrv4 I__5637 (
            .O(N__30021),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__5636 (
            .O(N__30016),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__5635 (
            .O(N__30007),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__5634 (
            .O(N__29998),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__5633 (
            .O(N__29989),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__5632 (
            .O(N__29980),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__5631 (
            .O(N__29975),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__5630 (
            .O(N__29960),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CascadeMux I__5629 (
            .O(N__29957),
            .I(N__29954));
    InMux I__5628 (
            .O(N__29954),
            .I(N__29951));
    LocalMux I__5627 (
            .O(N__29951),
            .I(N__29947));
    InMux I__5626 (
            .O(N__29950),
            .I(N__29944));
    Span4Mux_v I__5625 (
            .O(N__29947),
            .I(N__29941));
    LocalMux I__5624 (
            .O(N__29944),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__5623 (
            .O(N__29941),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__5622 (
            .O(N__29936),
            .I(N__29933));
    LocalMux I__5621 (
            .O(N__29933),
            .I(N__29927));
    CEMux I__5620 (
            .O(N__29932),
            .I(N__29924));
    CEMux I__5619 (
            .O(N__29931),
            .I(N__29921));
    CEMux I__5618 (
            .O(N__29930),
            .I(N__29918));
    Span4Mux_h I__5617 (
            .O(N__29927),
            .I(N__29915));
    LocalMux I__5616 (
            .O(N__29924),
            .I(N__29910));
    LocalMux I__5615 (
            .O(N__29921),
            .I(N__29910));
    LocalMux I__5614 (
            .O(N__29918),
            .I(N__29907));
    Odrv4 I__5613 (
            .O(N__29915),
            .I(\current_shift_inst.timer_s1.N_167_i ));
    Odrv4 I__5612 (
            .O(N__29910),
            .I(\current_shift_inst.timer_s1.N_167_i ));
    Odrv4 I__5611 (
            .O(N__29907),
            .I(\current_shift_inst.timer_s1.N_167_i ));
    InMux I__5610 (
            .O(N__29900),
            .I(N__29894));
    InMux I__5609 (
            .O(N__29899),
            .I(N__29894));
    LocalMux I__5608 (
            .O(N__29894),
            .I(N__29890));
    InMux I__5607 (
            .O(N__29893),
            .I(N__29887));
    Span4Mux_v I__5606 (
            .O(N__29890),
            .I(N__29884));
    LocalMux I__5605 (
            .O(N__29887),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__5604 (
            .O(N__29884),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__5603 (
            .O(N__29879),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__5602 (
            .O(N__29876),
            .I(N__29873));
    InMux I__5601 (
            .O(N__29873),
            .I(N__29869));
    InMux I__5600 (
            .O(N__29872),
            .I(N__29866));
    LocalMux I__5599 (
            .O(N__29869),
            .I(N__29862));
    LocalMux I__5598 (
            .O(N__29866),
            .I(N__29859));
    InMux I__5597 (
            .O(N__29865),
            .I(N__29856));
    Span4Mux_v I__5596 (
            .O(N__29862),
            .I(N__29851));
    Span4Mux_v I__5595 (
            .O(N__29859),
            .I(N__29851));
    LocalMux I__5594 (
            .O(N__29856),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__5593 (
            .O(N__29851),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__5592 (
            .O(N__29846),
            .I(bfn_13_26_0_));
    CascadeMux I__5591 (
            .O(N__29843),
            .I(N__29839));
    CascadeMux I__5590 (
            .O(N__29842),
            .I(N__29836));
    InMux I__5589 (
            .O(N__29839),
            .I(N__29833));
    InMux I__5588 (
            .O(N__29836),
            .I(N__29830));
    LocalMux I__5587 (
            .O(N__29833),
            .I(N__29826));
    LocalMux I__5586 (
            .O(N__29830),
            .I(N__29823));
    InMux I__5585 (
            .O(N__29829),
            .I(N__29820));
    Span4Mux_v I__5584 (
            .O(N__29826),
            .I(N__29815));
    Span4Mux_v I__5583 (
            .O(N__29823),
            .I(N__29815));
    LocalMux I__5582 (
            .O(N__29820),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__5581 (
            .O(N__29815),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__5580 (
            .O(N__29810),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__5579 (
            .O(N__29807),
            .I(N__29801));
    InMux I__5578 (
            .O(N__29806),
            .I(N__29801));
    LocalMux I__5577 (
            .O(N__29801),
            .I(N__29797));
    InMux I__5576 (
            .O(N__29800),
            .I(N__29794));
    Span4Mux_v I__5575 (
            .O(N__29797),
            .I(N__29791));
    LocalMux I__5574 (
            .O(N__29794),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__5573 (
            .O(N__29791),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__5572 (
            .O(N__29786),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__5571 (
            .O(N__29783),
            .I(N__29776));
    InMux I__5570 (
            .O(N__29782),
            .I(N__29776));
    InMux I__5569 (
            .O(N__29781),
            .I(N__29773));
    LocalMux I__5568 (
            .O(N__29776),
            .I(N__29770));
    LocalMux I__5567 (
            .O(N__29773),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv12 I__5566 (
            .O(N__29770),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__5565 (
            .O(N__29765),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__5564 (
            .O(N__29762),
            .I(N__29758));
    CascadeMux I__5563 (
            .O(N__29761),
            .I(N__29755));
    InMux I__5562 (
            .O(N__29758),
            .I(N__29750));
    InMux I__5561 (
            .O(N__29755),
            .I(N__29750));
    LocalMux I__5560 (
            .O(N__29750),
            .I(N__29746));
    InMux I__5559 (
            .O(N__29749),
            .I(N__29743));
    Span4Mux_v I__5558 (
            .O(N__29746),
            .I(N__29740));
    LocalMux I__5557 (
            .O(N__29743),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__5556 (
            .O(N__29740),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__5555 (
            .O(N__29735),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__5554 (
            .O(N__29732),
            .I(N__29728));
    CascadeMux I__5553 (
            .O(N__29731),
            .I(N__29725));
    InMux I__5552 (
            .O(N__29728),
            .I(N__29720));
    InMux I__5551 (
            .O(N__29725),
            .I(N__29720));
    LocalMux I__5550 (
            .O(N__29720),
            .I(N__29716));
    InMux I__5549 (
            .O(N__29719),
            .I(N__29713));
    Span4Mux_v I__5548 (
            .O(N__29716),
            .I(N__29710));
    LocalMux I__5547 (
            .O(N__29713),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__5546 (
            .O(N__29710),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__5545 (
            .O(N__29705),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__5544 (
            .O(N__29702),
            .I(N__29699));
    InMux I__5543 (
            .O(N__29699),
            .I(N__29694));
    InMux I__5542 (
            .O(N__29698),
            .I(N__29691));
    InMux I__5541 (
            .O(N__29697),
            .I(N__29688));
    LocalMux I__5540 (
            .O(N__29694),
            .I(N__29683));
    LocalMux I__5539 (
            .O(N__29691),
            .I(N__29683));
    LocalMux I__5538 (
            .O(N__29688),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv12 I__5537 (
            .O(N__29683),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__5536 (
            .O(N__29678),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    CascadeMux I__5535 (
            .O(N__29675),
            .I(N__29672));
    InMux I__5534 (
            .O(N__29672),
            .I(N__29668));
    InMux I__5533 (
            .O(N__29671),
            .I(N__29665));
    LocalMux I__5532 (
            .O(N__29668),
            .I(N__29659));
    LocalMux I__5531 (
            .O(N__29665),
            .I(N__29659));
    InMux I__5530 (
            .O(N__29664),
            .I(N__29656));
    Span4Mux_v I__5529 (
            .O(N__29659),
            .I(N__29653));
    LocalMux I__5528 (
            .O(N__29656),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__5527 (
            .O(N__29653),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__5526 (
            .O(N__29648),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__5525 (
            .O(N__29645),
            .I(N__29639));
    InMux I__5524 (
            .O(N__29644),
            .I(N__29639));
    LocalMux I__5523 (
            .O(N__29639),
            .I(N__29635));
    InMux I__5522 (
            .O(N__29638),
            .I(N__29632));
    Span4Mux_v I__5521 (
            .O(N__29635),
            .I(N__29629));
    LocalMux I__5520 (
            .O(N__29632),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__5519 (
            .O(N__29629),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__5518 (
            .O(N__29624),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__5517 (
            .O(N__29621),
            .I(N__29618));
    InMux I__5516 (
            .O(N__29618),
            .I(N__29615));
    LocalMux I__5515 (
            .O(N__29615),
            .I(N__29610));
    InMux I__5514 (
            .O(N__29614),
            .I(N__29607));
    InMux I__5513 (
            .O(N__29613),
            .I(N__29604));
    Span4Mux_v I__5512 (
            .O(N__29610),
            .I(N__29601));
    LocalMux I__5511 (
            .O(N__29607),
            .I(N__29598));
    LocalMux I__5510 (
            .O(N__29604),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__5509 (
            .O(N__29601),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv12 I__5508 (
            .O(N__29598),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__5507 (
            .O(N__29591),
            .I(bfn_13_25_0_));
    CascadeMux I__5506 (
            .O(N__29588),
            .I(N__29585));
    InMux I__5505 (
            .O(N__29585),
            .I(N__29581));
    CascadeMux I__5504 (
            .O(N__29584),
            .I(N__29578));
    LocalMux I__5503 (
            .O(N__29581),
            .I(N__29574));
    InMux I__5502 (
            .O(N__29578),
            .I(N__29571));
    InMux I__5501 (
            .O(N__29577),
            .I(N__29568));
    Span4Mux_v I__5500 (
            .O(N__29574),
            .I(N__29565));
    LocalMux I__5499 (
            .O(N__29571),
            .I(N__29562));
    LocalMux I__5498 (
            .O(N__29568),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__5497 (
            .O(N__29565),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv12 I__5496 (
            .O(N__29562),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__5495 (
            .O(N__29555),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__5494 (
            .O(N__29552),
            .I(N__29546));
    InMux I__5493 (
            .O(N__29551),
            .I(N__29546));
    LocalMux I__5492 (
            .O(N__29546),
            .I(N__29542));
    InMux I__5491 (
            .O(N__29545),
            .I(N__29539));
    Span4Mux_v I__5490 (
            .O(N__29542),
            .I(N__29536));
    LocalMux I__5489 (
            .O(N__29539),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__5488 (
            .O(N__29536),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__5487 (
            .O(N__29531),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__5486 (
            .O(N__29528),
            .I(N__29521));
    InMux I__5485 (
            .O(N__29527),
            .I(N__29521));
    InMux I__5484 (
            .O(N__29526),
            .I(N__29518));
    LocalMux I__5483 (
            .O(N__29521),
            .I(N__29515));
    LocalMux I__5482 (
            .O(N__29518),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv12 I__5481 (
            .O(N__29515),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__5480 (
            .O(N__29510),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    CascadeMux I__5479 (
            .O(N__29507),
            .I(N__29503));
    CascadeMux I__5478 (
            .O(N__29506),
            .I(N__29500));
    InMux I__5477 (
            .O(N__29503),
            .I(N__29495));
    InMux I__5476 (
            .O(N__29500),
            .I(N__29495));
    LocalMux I__5475 (
            .O(N__29495),
            .I(N__29491));
    InMux I__5474 (
            .O(N__29494),
            .I(N__29488));
    Span4Mux_v I__5473 (
            .O(N__29491),
            .I(N__29485));
    LocalMux I__5472 (
            .O(N__29488),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__5471 (
            .O(N__29485),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__5470 (
            .O(N__29480),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__5469 (
            .O(N__29477),
            .I(N__29473));
    CascadeMux I__5468 (
            .O(N__29476),
            .I(N__29470));
    InMux I__5467 (
            .O(N__29473),
            .I(N__29465));
    InMux I__5466 (
            .O(N__29470),
            .I(N__29465));
    LocalMux I__5465 (
            .O(N__29465),
            .I(N__29461));
    InMux I__5464 (
            .O(N__29464),
            .I(N__29458));
    Span4Mux_v I__5463 (
            .O(N__29461),
            .I(N__29455));
    LocalMux I__5462 (
            .O(N__29458),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__5461 (
            .O(N__29455),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__5460 (
            .O(N__29450),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__5459 (
            .O(N__29447),
            .I(N__29444));
    InMux I__5458 (
            .O(N__29444),
            .I(N__29440));
    InMux I__5457 (
            .O(N__29443),
            .I(N__29437));
    LocalMux I__5456 (
            .O(N__29440),
            .I(N__29431));
    LocalMux I__5455 (
            .O(N__29437),
            .I(N__29431));
    InMux I__5454 (
            .O(N__29436),
            .I(N__29428));
    Span4Mux_v I__5453 (
            .O(N__29431),
            .I(N__29425));
    LocalMux I__5452 (
            .O(N__29428),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__5451 (
            .O(N__29425),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__5450 (
            .O(N__29420),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__5449 (
            .O(N__29417),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__5448 (
            .O(N__29414),
            .I(N__29407));
    InMux I__5447 (
            .O(N__29413),
            .I(N__29407));
    InMux I__5446 (
            .O(N__29412),
            .I(N__29404));
    LocalMux I__5445 (
            .O(N__29407),
            .I(N__29400));
    LocalMux I__5444 (
            .O(N__29404),
            .I(N__29397));
    InMux I__5443 (
            .O(N__29403),
            .I(N__29394));
    Span4Mux_v I__5442 (
            .O(N__29400),
            .I(N__29391));
    Odrv12 I__5441 (
            .O(N__29397),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__5440 (
            .O(N__29394),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__5439 (
            .O(N__29391),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__5438 (
            .O(N__29384),
            .I(N__29381));
    LocalMux I__5437 (
            .O(N__29381),
            .I(N__29378));
    Odrv12 I__5436 (
            .O(N__29378),
            .I(s2_phy_c));
    InMux I__5435 (
            .O(N__29375),
            .I(bfn_13_24_0_));
    InMux I__5434 (
            .O(N__29372),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__5433 (
            .O(N__29369),
            .I(N__29362));
    InMux I__5432 (
            .O(N__29368),
            .I(N__29362));
    InMux I__5431 (
            .O(N__29367),
            .I(N__29359));
    LocalMux I__5430 (
            .O(N__29362),
            .I(N__29356));
    LocalMux I__5429 (
            .O(N__29359),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv12 I__5428 (
            .O(N__29356),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__5427 (
            .O(N__29351),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    CascadeMux I__5426 (
            .O(N__29348),
            .I(N__29344));
    InMux I__5425 (
            .O(N__29347),
            .I(N__29340));
    InMux I__5424 (
            .O(N__29344),
            .I(N__29337));
    InMux I__5423 (
            .O(N__29343),
            .I(N__29334));
    LocalMux I__5422 (
            .O(N__29340),
            .I(N__29327));
    LocalMux I__5421 (
            .O(N__29337),
            .I(N__29327));
    LocalMux I__5420 (
            .O(N__29334),
            .I(N__29327));
    Odrv12 I__5419 (
            .O(N__29327),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__5418 (
            .O(N__29324),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__5417 (
            .O(N__29321),
            .I(N__29317));
    InMux I__5416 (
            .O(N__29320),
            .I(N__29314));
    InMux I__5415 (
            .O(N__29317),
            .I(N__29311));
    LocalMux I__5414 (
            .O(N__29314),
            .I(N__29305));
    LocalMux I__5413 (
            .O(N__29311),
            .I(N__29305));
    InMux I__5412 (
            .O(N__29310),
            .I(N__29302));
    Span4Mux_v I__5411 (
            .O(N__29305),
            .I(N__29299));
    LocalMux I__5410 (
            .O(N__29302),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__5409 (
            .O(N__29299),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__5408 (
            .O(N__29294),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__5407 (
            .O(N__29291),
            .I(N__29288));
    InMux I__5406 (
            .O(N__29288),
            .I(N__29284));
    InMux I__5405 (
            .O(N__29287),
            .I(N__29281));
    LocalMux I__5404 (
            .O(N__29284),
            .I(N__29275));
    LocalMux I__5403 (
            .O(N__29281),
            .I(N__29275));
    InMux I__5402 (
            .O(N__29280),
            .I(N__29272));
    Span4Mux_v I__5401 (
            .O(N__29275),
            .I(N__29269));
    LocalMux I__5400 (
            .O(N__29272),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__5399 (
            .O(N__29269),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__5398 (
            .O(N__29264),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    CascadeMux I__5397 (
            .O(N__29261),
            .I(N__29257));
    CascadeMux I__5396 (
            .O(N__29260),
            .I(N__29254));
    InMux I__5395 (
            .O(N__29257),
            .I(N__29249));
    InMux I__5394 (
            .O(N__29254),
            .I(N__29249));
    LocalMux I__5393 (
            .O(N__29249),
            .I(N__29245));
    InMux I__5392 (
            .O(N__29248),
            .I(N__29242));
    Span4Mux_v I__5391 (
            .O(N__29245),
            .I(N__29239));
    LocalMux I__5390 (
            .O(N__29242),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__5389 (
            .O(N__29239),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__5388 (
            .O(N__29234),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__5387 (
            .O(N__29231),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__5386 (
            .O(N__29228),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__5385 (
            .O(N__29225),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__5384 (
            .O(N__29222),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__5383 (
            .O(N__29219),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__5382 (
            .O(N__29216),
            .I(bfn_13_22_0_));
    InMux I__5381 (
            .O(N__29213),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__5380 (
            .O(N__29210),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__5379 (
            .O(N__29207),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__5378 (
            .O(N__29204),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__5377 (
            .O(N__29201),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__5376 (
            .O(N__29198),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__5375 (
            .O(N__29195),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__5374 (
            .O(N__29192),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__5373 (
            .O(N__29189),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__5372 (
            .O(N__29186),
            .I(bfn_13_21_0_));
    InMux I__5371 (
            .O(N__29183),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__5370 (
            .O(N__29180),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__5369 (
            .O(N__29177),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__5368 (
            .O(N__29174),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__5367 (
            .O(N__29171),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__5366 (
            .O(N__29168),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__5365 (
            .O(N__29165),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__5364 (
            .O(N__29162),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__5363 (
            .O(N__29159),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__5362 (
            .O(N__29156),
            .I(bfn_13_20_0_));
    InMux I__5361 (
            .O(N__29153),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__5360 (
            .O(N__29150),
            .I(N__29147));
    LocalMux I__5359 (
            .O(N__29147),
            .I(\current_shift_inst.un38_control_input_cry_1_c_RNOZ0 ));
    InMux I__5358 (
            .O(N__29144),
            .I(N__29140));
    InMux I__5357 (
            .O(N__29143),
            .I(N__29137));
    LocalMux I__5356 (
            .O(N__29140),
            .I(N__29132));
    LocalMux I__5355 (
            .O(N__29137),
            .I(N__29129));
    InMux I__5354 (
            .O(N__29136),
            .I(N__29126));
    InMux I__5353 (
            .O(N__29135),
            .I(N__29123));
    Span12Mux_v I__5352 (
            .O(N__29132),
            .I(N__29120));
    Span12Mux_v I__5351 (
            .O(N__29129),
            .I(N__29117));
    LocalMux I__5350 (
            .O(N__29126),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__5349 (
            .O(N__29123),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv12 I__5348 (
            .O(N__29120),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv12 I__5347 (
            .O(N__29117),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__5346 (
            .O(N__29108),
            .I(N__29105));
    LocalMux I__5345 (
            .O(N__29105),
            .I(N__29101));
    InMux I__5344 (
            .O(N__29104),
            .I(N__29098));
    Span4Mux_v I__5343 (
            .O(N__29101),
            .I(N__29094));
    LocalMux I__5342 (
            .O(N__29098),
            .I(N__29091));
    InMux I__5341 (
            .O(N__29097),
            .I(N__29088));
    Span4Mux_h I__5340 (
            .O(N__29094),
            .I(N__29083));
    Span4Mux_v I__5339 (
            .O(N__29091),
            .I(N__29083));
    LocalMux I__5338 (
            .O(N__29088),
            .I(N__29080));
    Span4Mux_v I__5337 (
            .O(N__29083),
            .I(N__29077));
    Span12Mux_v I__5336 (
            .O(N__29080),
            .I(N__29074));
    Span4Mux_v I__5335 (
            .O(N__29077),
            .I(N__29071));
    Odrv12 I__5334 (
            .O(N__29074),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__5333 (
            .O(N__29071),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__5332 (
            .O(N__29066),
            .I(N__29062));
    InMux I__5331 (
            .O(N__29065),
            .I(N__29059));
    LocalMux I__5330 (
            .O(N__29062),
            .I(N__29056));
    LocalMux I__5329 (
            .O(N__29059),
            .I(N__29051));
    Span4Mux_v I__5328 (
            .O(N__29056),
            .I(N__29048));
    InMux I__5327 (
            .O(N__29055),
            .I(N__29043));
    InMux I__5326 (
            .O(N__29054),
            .I(N__29043));
    Span4Mux_v I__5325 (
            .O(N__29051),
            .I(N__29040));
    Odrv4 I__5324 (
            .O(N__29048),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__5323 (
            .O(N__29043),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__5322 (
            .O(N__29040),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__5321 (
            .O(N__29033),
            .I(N__29021));
    InMux I__5320 (
            .O(N__29032),
            .I(N__29021));
    InMux I__5319 (
            .O(N__29031),
            .I(N__29021));
    InMux I__5318 (
            .O(N__29030),
            .I(N__29021));
    LocalMux I__5317 (
            .O(N__29021),
            .I(N__28996));
    InMux I__5316 (
            .O(N__29020),
            .I(N__28987));
    InMux I__5315 (
            .O(N__29019),
            .I(N__28987));
    InMux I__5314 (
            .O(N__29018),
            .I(N__28987));
    InMux I__5313 (
            .O(N__29017),
            .I(N__28987));
    InMux I__5312 (
            .O(N__29016),
            .I(N__28978));
    InMux I__5311 (
            .O(N__29015),
            .I(N__28978));
    InMux I__5310 (
            .O(N__29014),
            .I(N__28978));
    InMux I__5309 (
            .O(N__29013),
            .I(N__28978));
    InMux I__5308 (
            .O(N__29012),
            .I(N__28969));
    InMux I__5307 (
            .O(N__29011),
            .I(N__28969));
    InMux I__5306 (
            .O(N__29010),
            .I(N__28960));
    InMux I__5305 (
            .O(N__29009),
            .I(N__28960));
    InMux I__5304 (
            .O(N__29008),
            .I(N__28960));
    InMux I__5303 (
            .O(N__29007),
            .I(N__28960));
    InMux I__5302 (
            .O(N__29006),
            .I(N__28951));
    InMux I__5301 (
            .O(N__29005),
            .I(N__28951));
    InMux I__5300 (
            .O(N__29004),
            .I(N__28951));
    InMux I__5299 (
            .O(N__29003),
            .I(N__28951));
    InMux I__5298 (
            .O(N__29002),
            .I(N__28942));
    InMux I__5297 (
            .O(N__29001),
            .I(N__28942));
    InMux I__5296 (
            .O(N__29000),
            .I(N__28942));
    InMux I__5295 (
            .O(N__28999),
            .I(N__28942));
    Span4Mux_v I__5294 (
            .O(N__28996),
            .I(N__28935));
    LocalMux I__5293 (
            .O(N__28987),
            .I(N__28935));
    LocalMux I__5292 (
            .O(N__28978),
            .I(N__28935));
    InMux I__5291 (
            .O(N__28977),
            .I(N__28926));
    InMux I__5290 (
            .O(N__28976),
            .I(N__28926));
    InMux I__5289 (
            .O(N__28975),
            .I(N__28926));
    InMux I__5288 (
            .O(N__28974),
            .I(N__28926));
    LocalMux I__5287 (
            .O(N__28969),
            .I(N__28921));
    LocalMux I__5286 (
            .O(N__28960),
            .I(N__28921));
    LocalMux I__5285 (
            .O(N__28951),
            .I(N__28918));
    LocalMux I__5284 (
            .O(N__28942),
            .I(N__28913));
    Span4Mux_v I__5283 (
            .O(N__28935),
            .I(N__28913));
    LocalMux I__5282 (
            .O(N__28926),
            .I(N__28910));
    Span4Mux_v I__5281 (
            .O(N__28921),
            .I(N__28901));
    Span4Mux_v I__5280 (
            .O(N__28918),
            .I(N__28901));
    Span4Mux_h I__5279 (
            .O(N__28913),
            .I(N__28901));
    Span4Mux_h I__5278 (
            .O(N__28910),
            .I(N__28901));
    Span4Mux_h I__5277 (
            .O(N__28901),
            .I(N__28898));
    Odrv4 I__5276 (
            .O(N__28898),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    CascadeMux I__5275 (
            .O(N__28895),
            .I(N__28891));
    InMux I__5274 (
            .O(N__28894),
            .I(N__28887));
    InMux I__5273 (
            .O(N__28891),
            .I(N__28884));
    InMux I__5272 (
            .O(N__28890),
            .I(N__28881));
    LocalMux I__5271 (
            .O(N__28887),
            .I(N__28878));
    LocalMux I__5270 (
            .O(N__28884),
            .I(N__28875));
    LocalMux I__5269 (
            .O(N__28881),
            .I(N__28872));
    Span4Mux_h I__5268 (
            .O(N__28878),
            .I(N__28867));
    Span4Mux_v I__5267 (
            .O(N__28875),
            .I(N__28867));
    Span4Mux_v I__5266 (
            .O(N__28872),
            .I(N__28864));
    Odrv4 I__5265 (
            .O(N__28867),
            .I(il_max_comp1_D2));
    Odrv4 I__5264 (
            .O(N__28864),
            .I(il_max_comp1_D2));
    InMux I__5263 (
            .O(N__28859),
            .I(N__28853));
    InMux I__5262 (
            .O(N__28858),
            .I(N__28845));
    InMux I__5261 (
            .O(N__28857),
            .I(N__28845));
    InMux I__5260 (
            .O(N__28856),
            .I(N__28845));
    LocalMux I__5259 (
            .O(N__28853),
            .I(N__28842));
    InMux I__5258 (
            .O(N__28852),
            .I(N__28839));
    LocalMux I__5257 (
            .O(N__28845),
            .I(N__28835));
    Span4Mux_v I__5256 (
            .O(N__28842),
            .I(N__28830));
    LocalMux I__5255 (
            .O(N__28839),
            .I(N__28830));
    InMux I__5254 (
            .O(N__28838),
            .I(N__28827));
    Span4Mux_h I__5253 (
            .O(N__28835),
            .I(N__28824));
    Span4Mux_h I__5252 (
            .O(N__28830),
            .I(N__28821));
    LocalMux I__5251 (
            .O(N__28827),
            .I(state_3));
    Odrv4 I__5250 (
            .O(N__28824),
            .I(state_3));
    Odrv4 I__5249 (
            .O(N__28821),
            .I(state_3));
    CascadeMux I__5248 (
            .O(N__28814),
            .I(N__28810));
    CascadeMux I__5247 (
            .O(N__28813),
            .I(N__28805));
    InMux I__5246 (
            .O(N__28810),
            .I(N__28801));
    InMux I__5245 (
            .O(N__28809),
            .I(N__28798));
    InMux I__5244 (
            .O(N__28808),
            .I(N__28794));
    InMux I__5243 (
            .O(N__28805),
            .I(N__28789));
    InMux I__5242 (
            .O(N__28804),
            .I(N__28789));
    LocalMux I__5241 (
            .O(N__28801),
            .I(N__28786));
    LocalMux I__5240 (
            .O(N__28798),
            .I(N__28783));
    InMux I__5239 (
            .O(N__28797),
            .I(N__28780));
    LocalMux I__5238 (
            .O(N__28794),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__5237 (
            .O(N__28789),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__5236 (
            .O(N__28786),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__5235 (
            .O(N__28783),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__5234 (
            .O(N__28780),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__5233 (
            .O(N__28769),
            .I(N__28766));
    InMux I__5232 (
            .O(N__28766),
            .I(N__28763));
    LocalMux I__5231 (
            .O(N__28763),
            .I(N__28758));
    InMux I__5230 (
            .O(N__28762),
            .I(N__28755));
    InMux I__5229 (
            .O(N__28761),
            .I(N__28752));
    Span4Mux_v I__5228 (
            .O(N__28758),
            .I(N__28749));
    LocalMux I__5227 (
            .O(N__28755),
            .I(N__28744));
    LocalMux I__5226 (
            .O(N__28752),
            .I(N__28744));
    Span4Mux_h I__5225 (
            .O(N__28749),
            .I(N__28741));
    Span4Mux_v I__5224 (
            .O(N__28744),
            .I(N__28738));
    Odrv4 I__5223 (
            .O(N__28741),
            .I(il_min_comp1_D2));
    Odrv4 I__5222 (
            .O(N__28738),
            .I(il_min_comp1_D2));
    InMux I__5221 (
            .O(N__28733),
            .I(N__28729));
    InMux I__5220 (
            .O(N__28732),
            .I(N__28726));
    LocalMux I__5219 (
            .O(N__28729),
            .I(N__28720));
    LocalMux I__5218 (
            .O(N__28726),
            .I(N__28720));
    InMux I__5217 (
            .O(N__28725),
            .I(N__28717));
    Span4Mux_v I__5216 (
            .O(N__28720),
            .I(N__28714));
    LocalMux I__5215 (
            .O(N__28717),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv4 I__5214 (
            .O(N__28714),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__5213 (
            .O(N__28709),
            .I(N__28706));
    LocalMux I__5212 (
            .O(N__28706),
            .I(N__28702));
    InMux I__5211 (
            .O(N__28705),
            .I(N__28698));
    Span4Mux_h I__5210 (
            .O(N__28702),
            .I(N__28695));
    InMux I__5209 (
            .O(N__28701),
            .I(N__28692));
    LocalMux I__5208 (
            .O(N__28698),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__5207 (
            .O(N__28695),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__5206 (
            .O(N__28692),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__5205 (
            .O(N__28685),
            .I(N__28682));
    LocalMux I__5204 (
            .O(N__28682),
            .I(N__28679));
    Odrv12 I__5203 (
            .O(N__28679),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ));
    InMux I__5202 (
            .O(N__28676),
            .I(N__28673));
    LocalMux I__5201 (
            .O(N__28673),
            .I(N__28670));
    Span4Mux_h I__5200 (
            .O(N__28670),
            .I(N__28667));
    Odrv4 I__5199 (
            .O(N__28667),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ));
    InMux I__5198 (
            .O(N__28664),
            .I(N__28658));
    InMux I__5197 (
            .O(N__28663),
            .I(N__28655));
    InMux I__5196 (
            .O(N__28662),
            .I(N__28652));
    InMux I__5195 (
            .O(N__28661),
            .I(N__28649));
    LocalMux I__5194 (
            .O(N__28658),
            .I(N__28646));
    LocalMux I__5193 (
            .O(N__28655),
            .I(N__28641));
    LocalMux I__5192 (
            .O(N__28652),
            .I(N__28641));
    LocalMux I__5191 (
            .O(N__28649),
            .I(N__28637));
    Span12Mux_h I__5190 (
            .O(N__28646),
            .I(N__28632));
    Span12Mux_v I__5189 (
            .O(N__28641),
            .I(N__28632));
    InMux I__5188 (
            .O(N__28640),
            .I(N__28629));
    Odrv4 I__5187 (
            .O(N__28637),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv12 I__5186 (
            .O(N__28632),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__5185 (
            .O(N__28629),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__5184 (
            .O(N__28622),
            .I(N__28619));
    LocalMux I__5183 (
            .O(N__28619),
            .I(N__28616));
    Span4Mux_v I__5182 (
            .O(N__28616),
            .I(N__28613));
    Odrv4 I__5181 (
            .O(N__28613),
            .I(\current_shift_inst.un38_control_input_cry_19_c_RNOZ0 ));
    InMux I__5180 (
            .O(N__28610),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ));
    InMux I__5179 (
            .O(N__28607),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ));
    InMux I__5178 (
            .O(N__28604),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ));
    InMux I__5177 (
            .O(N__28601),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_31 ));
    CascadeMux I__5176 (
            .O(N__28598),
            .I(N__28593));
    CascadeMux I__5175 (
            .O(N__28597),
            .I(N__28590));
    InMux I__5174 (
            .O(N__28596),
            .I(N__28580));
    InMux I__5173 (
            .O(N__28593),
            .I(N__28580));
    InMux I__5172 (
            .O(N__28590),
            .I(N__28580));
    InMux I__5171 (
            .O(N__28589),
            .I(N__28580));
    LocalMux I__5170 (
            .O(N__28580),
            .I(N__28575));
    InMux I__5169 (
            .O(N__28579),
            .I(N__28572));
    InMux I__5168 (
            .O(N__28578),
            .I(N__28569));
    Span4Mux_h I__5167 (
            .O(N__28575),
            .I(N__28566));
    LocalMux I__5166 (
            .O(N__28572),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__5165 (
            .O(N__28569),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__5164 (
            .O(N__28566),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__5163 (
            .O(N__28559),
            .I(N__28556));
    LocalMux I__5162 (
            .O(N__28556),
            .I(N__28549));
    InMux I__5161 (
            .O(N__28555),
            .I(N__28540));
    InMux I__5160 (
            .O(N__28554),
            .I(N__28540));
    InMux I__5159 (
            .O(N__28553),
            .I(N__28540));
    InMux I__5158 (
            .O(N__28552),
            .I(N__28540));
    Span4Mux_h I__5157 (
            .O(N__28549),
            .I(N__28537));
    LocalMux I__5156 (
            .O(N__28540),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__5155 (
            .O(N__28537),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__5154 (
            .O(N__28532),
            .I(N__28529));
    LocalMux I__5153 (
            .O(N__28529),
            .I(N__28526));
    Span4Mux_v I__5152 (
            .O(N__28526),
            .I(N__28523));
    Odrv4 I__5151 (
            .O(N__28523),
            .I(\phase_controller_inst1.stoper_tr.N_45 ));
    InMux I__5150 (
            .O(N__28520),
            .I(N__28516));
    InMux I__5149 (
            .O(N__28519),
            .I(N__28513));
    LocalMux I__5148 (
            .O(N__28516),
            .I(N__28510));
    LocalMux I__5147 (
            .O(N__28513),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    Odrv12 I__5146 (
            .O(N__28510),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    InMux I__5145 (
            .O(N__28505),
            .I(N__28502));
    LocalMux I__5144 (
            .O(N__28502),
            .I(N__28499));
    Odrv12 I__5143 (
            .O(N__28499),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ));
    InMux I__5142 (
            .O(N__28496),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ));
    InMux I__5141 (
            .O(N__28493),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ));
    InMux I__5140 (
            .O(N__28490),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ));
    InMux I__5139 (
            .O(N__28487),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ));
    InMux I__5138 (
            .O(N__28484),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ));
    InMux I__5137 (
            .O(N__28481),
            .I(bfn_13_14_0_));
    CascadeMux I__5136 (
            .O(N__28478),
            .I(N__28475));
    InMux I__5135 (
            .O(N__28475),
            .I(N__28472));
    LocalMux I__5134 (
            .O(N__28472),
            .I(N__28469));
    Span4Mux_v I__5133 (
            .O(N__28469),
            .I(N__28466));
    Odrv4 I__5132 (
            .O(N__28466),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ));
    InMux I__5131 (
            .O(N__28463),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ));
    InMux I__5130 (
            .O(N__28460),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ));
    InMux I__5129 (
            .O(N__28457),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ));
    InMux I__5128 (
            .O(N__28454),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ));
    InMux I__5127 (
            .O(N__28451),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ));
    InMux I__5126 (
            .O(N__28448),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ));
    InMux I__5125 (
            .O(N__28445),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ));
    InMux I__5124 (
            .O(N__28442),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ));
    InMux I__5123 (
            .O(N__28439),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ));
    InMux I__5122 (
            .O(N__28436),
            .I(bfn_13_13_0_));
    InMux I__5121 (
            .O(N__28433),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ));
    InMux I__5120 (
            .O(N__28430),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ));
    InMux I__5119 (
            .O(N__28427),
            .I(N__28424));
    LocalMux I__5118 (
            .O(N__28424),
            .I(N__28420));
    InMux I__5117 (
            .O(N__28423),
            .I(N__28417));
    Span4Mux_h I__5116 (
            .O(N__28420),
            .I(N__28414));
    LocalMux I__5115 (
            .O(N__28417),
            .I(N__28411));
    Odrv4 I__5114 (
            .O(N__28414),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv4 I__5113 (
            .O(N__28411),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__5112 (
            .O(N__28406),
            .I(N__28403));
    LocalMux I__5111 (
            .O(N__28403),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ));
    InMux I__5110 (
            .O(N__28400),
            .I(N__28397));
    LocalMux I__5109 (
            .O(N__28397),
            .I(N__28394));
    Span4Mux_h I__5108 (
            .O(N__28394),
            .I(N__28390));
    InMux I__5107 (
            .O(N__28393),
            .I(N__28387));
    Odrv4 I__5106 (
            .O(N__28390),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    LocalMux I__5105 (
            .O(N__28387),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__5104 (
            .O(N__28382),
            .I(N__28379));
    LocalMux I__5103 (
            .O(N__28379),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ));
    InMux I__5102 (
            .O(N__28376),
            .I(N__28373));
    LocalMux I__5101 (
            .O(N__28373),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ));
    CascadeMux I__5100 (
            .O(N__28370),
            .I(N__28367));
    InMux I__5099 (
            .O(N__28367),
            .I(N__28364));
    LocalMux I__5098 (
            .O(N__28364),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_4 ));
    InMux I__5097 (
            .O(N__28361),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ));
    InMux I__5096 (
            .O(N__28358),
            .I(N__28355));
    LocalMux I__5095 (
            .O(N__28355),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ));
    CascadeMux I__5094 (
            .O(N__28352),
            .I(N__28349));
    InMux I__5093 (
            .O(N__28349),
            .I(N__28346));
    LocalMux I__5092 (
            .O(N__28346),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_5 ));
    InMux I__5091 (
            .O(N__28343),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ));
    InMux I__5090 (
            .O(N__28340),
            .I(N__28337));
    LocalMux I__5089 (
            .O(N__28337),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ));
    InMux I__5088 (
            .O(N__28334),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ));
    InMux I__5087 (
            .O(N__28331),
            .I(N__28328));
    LocalMux I__5086 (
            .O(N__28328),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ));
    InMux I__5085 (
            .O(N__28325),
            .I(N__28322));
    LocalMux I__5084 (
            .O(N__28322),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_7 ));
    InMux I__5083 (
            .O(N__28319),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ));
    InMux I__5082 (
            .O(N__28316),
            .I(N__28313));
    LocalMux I__5081 (
            .O(N__28313),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ));
    InMux I__5080 (
            .O(N__28310),
            .I(bfn_13_12_0_));
    InMux I__5079 (
            .O(N__28307),
            .I(N__28304));
    LocalMux I__5078 (
            .O(N__28304),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ));
    InMux I__5077 (
            .O(N__28301),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ));
    InMux I__5076 (
            .O(N__28298),
            .I(N__28295));
    LocalMux I__5075 (
            .O(N__28295),
            .I(N__28292));
    Span4Mux_h I__5074 (
            .O(N__28292),
            .I(N__28287));
    InMux I__5073 (
            .O(N__28291),
            .I(N__28282));
    InMux I__5072 (
            .O(N__28290),
            .I(N__28282));
    Odrv4 I__5071 (
            .O(N__28287),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    LocalMux I__5070 (
            .O(N__28282),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__5069 (
            .O(N__28277),
            .I(N__28274));
    LocalMux I__5068 (
            .O(N__28274),
            .I(N__28271));
    Span4Mux_h I__5067 (
            .O(N__28271),
            .I(N__28266));
    InMux I__5066 (
            .O(N__28270),
            .I(N__28261));
    InMux I__5065 (
            .O(N__28269),
            .I(N__28261));
    Odrv4 I__5064 (
            .O(N__28266),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    LocalMux I__5063 (
            .O(N__28261),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__5062 (
            .O(N__28256),
            .I(N__28253));
    LocalMux I__5061 (
            .O(N__28253),
            .I(N__28249));
    InMux I__5060 (
            .O(N__28252),
            .I(N__28246));
    Span4Mux_h I__5059 (
            .O(N__28249),
            .I(N__28241));
    LocalMux I__5058 (
            .O(N__28246),
            .I(N__28241));
    Odrv4 I__5057 (
            .O(N__28241),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__5056 (
            .O(N__28238),
            .I(N__28235));
    LocalMux I__5055 (
            .O(N__28235),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ));
    InMux I__5054 (
            .O(N__28232),
            .I(N__28228));
    InMux I__5053 (
            .O(N__28231),
            .I(N__28225));
    LocalMux I__5052 (
            .O(N__28228),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    LocalMux I__5051 (
            .O(N__28225),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__5050 (
            .O(N__28220),
            .I(N__28217));
    LocalMux I__5049 (
            .O(N__28217),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ));
    InMux I__5048 (
            .O(N__28214),
            .I(N__28211));
    LocalMux I__5047 (
            .O(N__28211),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ));
    InMux I__5046 (
            .O(N__28208),
            .I(N__28205));
    LocalMux I__5045 (
            .O(N__28205),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__5044 (
            .O(N__28202),
            .I(N__28199));
    LocalMux I__5043 (
            .O(N__28199),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    CascadeMux I__5042 (
            .O(N__28196),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19_cascade_ ));
    CascadeMux I__5041 (
            .O(N__28193),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ));
    InMux I__5040 (
            .O(N__28190),
            .I(N__28187));
    LocalMux I__5039 (
            .O(N__28187),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ));
    InMux I__5038 (
            .O(N__28184),
            .I(N__28181));
    LocalMux I__5037 (
            .O(N__28181),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16 ));
    InMux I__5036 (
            .O(N__28178),
            .I(N__28175));
    LocalMux I__5035 (
            .O(N__28175),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ));
    InMux I__5034 (
            .O(N__28172),
            .I(N__28169));
    LocalMux I__5033 (
            .O(N__28169),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    InMux I__5032 (
            .O(N__28166),
            .I(N__28162));
    InMux I__5031 (
            .O(N__28165),
            .I(N__28159));
    LocalMux I__5030 (
            .O(N__28162),
            .I(\current_shift_inst.PI_CTRL.N_74_21 ));
    LocalMux I__5029 (
            .O(N__28159),
            .I(\current_shift_inst.PI_CTRL.N_74_21 ));
    InMux I__5028 (
            .O(N__28154),
            .I(N__28151));
    LocalMux I__5027 (
            .O(N__28151),
            .I(N__28148));
    Span4Mux_h I__5026 (
            .O(N__28148),
            .I(N__28144));
    InMux I__5025 (
            .O(N__28147),
            .I(N__28141));
    Odrv4 I__5024 (
            .O(N__28144),
            .I(\current_shift_inst.PI_CTRL.N_72 ));
    LocalMux I__5023 (
            .O(N__28141),
            .I(\current_shift_inst.PI_CTRL.N_72 ));
    InMux I__5022 (
            .O(N__28136),
            .I(N__28133));
    LocalMux I__5021 (
            .O(N__28133),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    InMux I__5020 (
            .O(N__28130),
            .I(N__28120));
    InMux I__5019 (
            .O(N__28129),
            .I(N__28120));
    InMux I__5018 (
            .O(N__28128),
            .I(N__28120));
    InMux I__5017 (
            .O(N__28127),
            .I(N__28117));
    LocalMux I__5016 (
            .O(N__28120),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__5015 (
            .O(N__28117),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__5014 (
            .O(N__28112),
            .I(N__28106));
    InMux I__5013 (
            .O(N__28111),
            .I(N__28099));
    InMux I__5012 (
            .O(N__28110),
            .I(N__28099));
    InMux I__5011 (
            .O(N__28109),
            .I(N__28099));
    LocalMux I__5010 (
            .O(N__28106),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__5009 (
            .O(N__28099),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    CascadeMux I__5008 (
            .O(N__28094),
            .I(N__28091));
    InMux I__5007 (
            .O(N__28091),
            .I(N__28083));
    InMux I__5006 (
            .O(N__28090),
            .I(N__28083));
    InMux I__5005 (
            .O(N__28089),
            .I(N__28078));
    InMux I__5004 (
            .O(N__28088),
            .I(N__28078));
    LocalMux I__5003 (
            .O(N__28083),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__5002 (
            .O(N__28078),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    IoInMux I__5001 (
            .O(N__28073),
            .I(N__28070));
    LocalMux I__5000 (
            .O(N__28070),
            .I(N__28067));
    IoSpan4Mux I__4999 (
            .O(N__28067),
            .I(N__28064));
    Span4Mux_s0_v I__4998 (
            .O(N__28064),
            .I(N__28061));
    Odrv4 I__4997 (
            .O(N__28061),
            .I(\pll_inst.red_c_i ));
    CascadeMux I__4996 (
            .O(N__28058),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18_cascade_ ));
    InMux I__4995 (
            .O(N__28055),
            .I(N__28052));
    LocalMux I__4994 (
            .O(N__28052),
            .I(\current_shift_inst.PI_CTRL.N_62 ));
    CascadeMux I__4993 (
            .O(N__28049),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_ ));
    InMux I__4992 (
            .O(N__28046),
            .I(N__28040));
    InMux I__4991 (
            .O(N__28045),
            .I(N__28040));
    LocalMux I__4990 (
            .O(N__28040),
            .I(\current_shift_inst.un38_control_input_axb_30 ));
    InMux I__4989 (
            .O(N__28037),
            .I(N__28033));
    InMux I__4988 (
            .O(N__28036),
            .I(N__28030));
    LocalMux I__4987 (
            .O(N__28033),
            .I(N__28027));
    LocalMux I__4986 (
            .O(N__28030),
            .I(N__28024));
    Odrv4 I__4985 (
            .O(N__28027),
            .I(\phase_controller_inst2.time_passed_RNI9M3O ));
    Odrv4 I__4984 (
            .O(N__28024),
            .I(\phase_controller_inst2.time_passed_RNI9M3O ));
    InMux I__4983 (
            .O(N__28019),
            .I(N__28016));
    LocalMux I__4982 (
            .O(N__28016),
            .I(N__28012));
    InMux I__4981 (
            .O(N__28015),
            .I(N__28006));
    Span4Mux_h I__4980 (
            .O(N__28012),
            .I(N__28003));
    InMux I__4979 (
            .O(N__28011),
            .I(N__28000));
    InMux I__4978 (
            .O(N__28010),
            .I(N__27995));
    InMux I__4977 (
            .O(N__28009),
            .I(N__27995));
    LocalMux I__4976 (
            .O(N__28006),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    Odrv4 I__4975 (
            .O(N__28003),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__4974 (
            .O(N__28000),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__4973 (
            .O(N__27995),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    IoInMux I__4972 (
            .O(N__27986),
            .I(N__27983));
    LocalMux I__4971 (
            .O(N__27983),
            .I(N__27980));
    Span4Mux_s3_v I__4970 (
            .O(N__27980),
            .I(N__27977));
    Span4Mux_h I__4969 (
            .O(N__27977),
            .I(N__27974));
    Span4Mux_v I__4968 (
            .O(N__27974),
            .I(N__27970));
    InMux I__4967 (
            .O(N__27973),
            .I(N__27967));
    Odrv4 I__4966 (
            .O(N__27970),
            .I(T01_c));
    LocalMux I__4965 (
            .O(N__27967),
            .I(T01_c));
    IoInMux I__4964 (
            .O(N__27962),
            .I(N__27959));
    LocalMux I__4963 (
            .O(N__27959),
            .I(N__27956));
    Span4Mux_s1_v I__4962 (
            .O(N__27956),
            .I(N__27953));
    Span4Mux_v I__4961 (
            .O(N__27953),
            .I(N__27948));
    InMux I__4960 (
            .O(N__27952),
            .I(N__27943));
    InMux I__4959 (
            .O(N__27951),
            .I(N__27943));
    Odrv4 I__4958 (
            .O(N__27948),
            .I(s1_phy_c));
    LocalMux I__4957 (
            .O(N__27943),
            .I(s1_phy_c));
    CascadeMux I__4956 (
            .O(N__27938),
            .I(N__27933));
    InMux I__4955 (
            .O(N__27937),
            .I(N__27930));
    InMux I__4954 (
            .O(N__27936),
            .I(N__27926));
    InMux I__4953 (
            .O(N__27933),
            .I(N__27923));
    LocalMux I__4952 (
            .O(N__27930),
            .I(N__27920));
    InMux I__4951 (
            .O(N__27929),
            .I(N__27917));
    LocalMux I__4950 (
            .O(N__27926),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__4949 (
            .O(N__27923),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    Odrv4 I__4948 (
            .O(N__27920),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__4947 (
            .O(N__27917),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__4946 (
            .O(N__27908),
            .I(N__27902));
    InMux I__4945 (
            .O(N__27907),
            .I(N__27899));
    InMux I__4944 (
            .O(N__27906),
            .I(N__27896));
    CascadeMux I__4943 (
            .O(N__27905),
            .I(N__27892));
    LocalMux I__4942 (
            .O(N__27902),
            .I(N__27888));
    LocalMux I__4941 (
            .O(N__27899),
            .I(N__27885));
    LocalMux I__4940 (
            .O(N__27896),
            .I(N__27882));
    InMux I__4939 (
            .O(N__27895),
            .I(N__27879));
    InMux I__4938 (
            .O(N__27892),
            .I(N__27876));
    InMux I__4937 (
            .O(N__27891),
            .I(N__27873));
    Span4Mux_h I__4936 (
            .O(N__27888),
            .I(N__27868));
    Span4Mux_v I__4935 (
            .O(N__27885),
            .I(N__27868));
    Span4Mux_h I__4934 (
            .O(N__27882),
            .I(N__27863));
    LocalMux I__4933 (
            .O(N__27879),
            .I(N__27863));
    LocalMux I__4932 (
            .O(N__27876),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__4931 (
            .O(N__27873),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__4930 (
            .O(N__27868),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__4929 (
            .O(N__27863),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    IoInMux I__4928 (
            .O(N__27854),
            .I(N__27851));
    LocalMux I__4927 (
            .O(N__27851),
            .I(N__27848));
    Span4Mux_s2_v I__4926 (
            .O(N__27848),
            .I(N__27845));
    Span4Mux_h I__4925 (
            .O(N__27845),
            .I(N__27841));
    InMux I__4924 (
            .O(N__27844),
            .I(N__27838));
    Odrv4 I__4923 (
            .O(N__27841),
            .I(T45_c));
    LocalMux I__4922 (
            .O(N__27838),
            .I(T45_c));
    IoInMux I__4921 (
            .O(N__27833),
            .I(N__27830));
    LocalMux I__4920 (
            .O(N__27830),
            .I(N__27827));
    Span4Mux_s1_v I__4919 (
            .O(N__27827),
            .I(N__27824));
    Odrv4 I__4918 (
            .O(N__27824),
            .I(\current_shift_inst.timer_s1.N_166_i ));
    InMux I__4917 (
            .O(N__27821),
            .I(N__27818));
    LocalMux I__4916 (
            .O(N__27818),
            .I(\current_shift_inst.control_input_1_axb_3 ));
    InMux I__4915 (
            .O(N__27815),
            .I(bfn_12_21_0_));
    InMux I__4914 (
            .O(N__27812),
            .I(N__27809));
    LocalMux I__4913 (
            .O(N__27809),
            .I(\current_shift_inst.control_input_1_axb_4 ));
    InMux I__4912 (
            .O(N__27806),
            .I(\current_shift_inst.un38_control_input_cry_23 ));
    InMux I__4911 (
            .O(N__27803),
            .I(N__27800));
    LocalMux I__4910 (
            .O(N__27800),
            .I(\current_shift_inst.control_input_1_axb_5 ));
    InMux I__4909 (
            .O(N__27797),
            .I(\current_shift_inst.un38_control_input_cry_24 ));
    InMux I__4908 (
            .O(N__27794),
            .I(N__27791));
    LocalMux I__4907 (
            .O(N__27791),
            .I(\current_shift_inst.control_input_1_axb_6 ));
    InMux I__4906 (
            .O(N__27788),
            .I(\current_shift_inst.un38_control_input_cry_25 ));
    InMux I__4905 (
            .O(N__27785),
            .I(N__27782));
    LocalMux I__4904 (
            .O(N__27782),
            .I(N__27779));
    Span4Mux_v I__4903 (
            .O(N__27779),
            .I(N__27776));
    Odrv4 I__4902 (
            .O(N__27776),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__4901 (
            .O(N__27773),
            .I(N__27770));
    LocalMux I__4900 (
            .O(N__27770),
            .I(\current_shift_inst.control_input_1_axb_7 ));
    InMux I__4899 (
            .O(N__27767),
            .I(\current_shift_inst.un38_control_input_cry_26 ));
    InMux I__4898 (
            .O(N__27764),
            .I(N__27761));
    LocalMux I__4897 (
            .O(N__27761),
            .I(\current_shift_inst.control_input_1_axb_8 ));
    InMux I__4896 (
            .O(N__27758),
            .I(\current_shift_inst.un38_control_input_cry_27 ));
    InMux I__4895 (
            .O(N__27755),
            .I(N__27752));
    LocalMux I__4894 (
            .O(N__27752),
            .I(\current_shift_inst.control_input_1_axb_9 ));
    InMux I__4893 (
            .O(N__27749),
            .I(\current_shift_inst.un38_control_input_cry_28 ));
    InMux I__4892 (
            .O(N__27746),
            .I(\current_shift_inst.un38_control_input_cry_29 ));
    CascadeMux I__4891 (
            .O(N__27743),
            .I(N__27740));
    InMux I__4890 (
            .O(N__27740),
            .I(N__27736));
    InMux I__4889 (
            .O(N__27739),
            .I(N__27733));
    LocalMux I__4888 (
            .O(N__27736),
            .I(\current_shift_inst.un38_control_input_cry_29_THRU_CO ));
    LocalMux I__4887 (
            .O(N__27733),
            .I(\current_shift_inst.un38_control_input_cry_29_THRU_CO ));
    InMux I__4886 (
            .O(N__27728),
            .I(N__27725));
    LocalMux I__4885 (
            .O(N__27725),
            .I(\current_shift_inst.control_input_1_axb_0 ));
    InMux I__4884 (
            .O(N__27722),
            .I(\current_shift_inst.un38_control_input_cry_19 ));
    InMux I__4883 (
            .O(N__27719),
            .I(N__27716));
    LocalMux I__4882 (
            .O(N__27716),
            .I(\current_shift_inst.control_input_1_axb_1 ));
    InMux I__4881 (
            .O(N__27713),
            .I(\current_shift_inst.un38_control_input_cry_20 ));
    InMux I__4880 (
            .O(N__27710),
            .I(N__27707));
    LocalMux I__4879 (
            .O(N__27707),
            .I(\current_shift_inst.control_input_1_axb_2 ));
    InMux I__4878 (
            .O(N__27704),
            .I(\current_shift_inst.un38_control_input_cry_21 ));
    InMux I__4877 (
            .O(N__27701),
            .I(N__27698));
    LocalMux I__4876 (
            .O(N__27698),
            .I(N__27695));
    Odrv12 I__4875 (
            .O(N__27695),
            .I(\current_shift_inst.un38_control_input_cry_7_c_RNOZ0 ));
    InMux I__4874 (
            .O(N__27692),
            .I(N__27689));
    LocalMux I__4873 (
            .O(N__27689),
            .I(\current_shift_inst.un38_control_input_cry_3_c_RNOZ0 ));
    InMux I__4872 (
            .O(N__27686),
            .I(N__27683));
    LocalMux I__4871 (
            .O(N__27683),
            .I(\current_shift_inst.un38_control_input_cry_4_c_RNOZ0 ));
    InMux I__4870 (
            .O(N__27680),
            .I(N__27676));
    InMux I__4869 (
            .O(N__27679),
            .I(N__27673));
    LocalMux I__4868 (
            .O(N__27676),
            .I(N__27670));
    LocalMux I__4867 (
            .O(N__27673),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__4866 (
            .O(N__27670),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__4865 (
            .O(N__27665),
            .I(N__27662));
    LocalMux I__4864 (
            .O(N__27662),
            .I(N__27659));
    Span4Mux_h I__4863 (
            .O(N__27659),
            .I(N__27656));
    Odrv4 I__4862 (
            .O(N__27656),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__4861 (
            .O(N__27653),
            .I(N__27650));
    InMux I__4860 (
            .O(N__27650),
            .I(N__27647));
    LocalMux I__4859 (
            .O(N__27647),
            .I(N__27644));
    Odrv4 I__4858 (
            .O(N__27644),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__4857 (
            .O(N__27641),
            .I(N__27638));
    LocalMux I__4856 (
            .O(N__27638),
            .I(N__27635));
    Span4Mux_h I__4855 (
            .O(N__27635),
            .I(N__27632));
    Odrv4 I__4854 (
            .O(N__27632),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    InMux I__4853 (
            .O(N__27629),
            .I(N__27625));
    InMux I__4852 (
            .O(N__27628),
            .I(N__27622));
    LocalMux I__4851 (
            .O(N__27625),
            .I(N__27619));
    LocalMux I__4850 (
            .O(N__27622),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__4849 (
            .O(N__27619),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__4848 (
            .O(N__27614),
            .I(N__27611));
    InMux I__4847 (
            .O(N__27611),
            .I(N__27608));
    LocalMux I__4846 (
            .O(N__27608),
            .I(N__27605));
    Odrv4 I__4845 (
            .O(N__27605),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__4844 (
            .O(N__27602),
            .I(N__27598));
    InMux I__4843 (
            .O(N__27601),
            .I(N__27595));
    LocalMux I__4842 (
            .O(N__27598),
            .I(N__27592));
    LocalMux I__4841 (
            .O(N__27595),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__4840 (
            .O(N__27592),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__4839 (
            .O(N__27587),
            .I(N__27584));
    LocalMux I__4838 (
            .O(N__27584),
            .I(N__27581));
    Span4Mux_v I__4837 (
            .O(N__27581),
            .I(N__27578));
    Odrv4 I__4836 (
            .O(N__27578),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__4835 (
            .O(N__27575),
            .I(N__27572));
    InMux I__4834 (
            .O(N__27572),
            .I(N__27569));
    LocalMux I__4833 (
            .O(N__27569),
            .I(N__27566));
    Odrv4 I__4832 (
            .O(N__27566),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ));
    InMux I__4831 (
            .O(N__27563),
            .I(N__27559));
    InMux I__4830 (
            .O(N__27562),
            .I(N__27556));
    LocalMux I__4829 (
            .O(N__27559),
            .I(N__27553));
    LocalMux I__4828 (
            .O(N__27556),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__4827 (
            .O(N__27553),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__4826 (
            .O(N__27548),
            .I(N__27545));
    LocalMux I__4825 (
            .O(N__27545),
            .I(N__27542));
    Span4Mux_h I__4824 (
            .O(N__27542),
            .I(N__27539));
    Odrv4 I__4823 (
            .O(N__27539),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__4822 (
            .O(N__27536),
            .I(N__27533));
    InMux I__4821 (
            .O(N__27533),
            .I(N__27530));
    LocalMux I__4820 (
            .O(N__27530),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ));
    InMux I__4819 (
            .O(N__27527),
            .I(N__27523));
    InMux I__4818 (
            .O(N__27526),
            .I(N__27520));
    LocalMux I__4817 (
            .O(N__27523),
            .I(N__27517));
    LocalMux I__4816 (
            .O(N__27520),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__4815 (
            .O(N__27517),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__4814 (
            .O(N__27512),
            .I(N__27509));
    LocalMux I__4813 (
            .O(N__27509),
            .I(N__27506));
    Span4Mux_v I__4812 (
            .O(N__27506),
            .I(N__27503));
    Odrv4 I__4811 (
            .O(N__27503),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__4810 (
            .O(N__27500),
            .I(N__27497));
    InMux I__4809 (
            .O(N__27497),
            .I(N__27494));
    LocalMux I__4808 (
            .O(N__27494),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ));
    InMux I__4807 (
            .O(N__27491),
            .I(N__27488));
    LocalMux I__4806 (
            .O(N__27488),
            .I(N__27485));
    Span4Mux_v I__4805 (
            .O(N__27485),
            .I(N__27482));
    Odrv4 I__4804 (
            .O(N__27482),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__4803 (
            .O(N__27479),
            .I(N__27475));
    InMux I__4802 (
            .O(N__27478),
            .I(N__27472));
    LocalMux I__4801 (
            .O(N__27475),
            .I(N__27469));
    LocalMux I__4800 (
            .O(N__27472),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__4799 (
            .O(N__27469),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__4798 (
            .O(N__27464),
            .I(N__27461));
    InMux I__4797 (
            .O(N__27461),
            .I(N__27458));
    LocalMux I__4796 (
            .O(N__27458),
            .I(N__27455));
    Odrv4 I__4795 (
            .O(N__27455),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ));
    InMux I__4794 (
            .O(N__27452),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__4793 (
            .O(N__27449),
            .I(N__27446));
    LocalMux I__4792 (
            .O(N__27446),
            .I(N__27442));
    InMux I__4791 (
            .O(N__27445),
            .I(N__27439));
    Span4Mux_h I__4790 (
            .O(N__27442),
            .I(N__27436));
    LocalMux I__4789 (
            .O(N__27439),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__4788 (
            .O(N__27436),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__4787 (
            .O(N__27431),
            .I(N__27428));
    LocalMux I__4786 (
            .O(N__27428),
            .I(N__27425));
    Span4Mux_v I__4785 (
            .O(N__27425),
            .I(N__27422));
    Odrv4 I__4784 (
            .O(N__27422),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__4783 (
            .O(N__27419),
            .I(N__27416));
    InMux I__4782 (
            .O(N__27416),
            .I(N__27413));
    LocalMux I__4781 (
            .O(N__27413),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__4780 (
            .O(N__27410),
            .I(N__27407));
    LocalMux I__4779 (
            .O(N__27407),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    InMux I__4778 (
            .O(N__27404),
            .I(N__27400));
    InMux I__4777 (
            .O(N__27403),
            .I(N__27397));
    LocalMux I__4776 (
            .O(N__27400),
            .I(N__27394));
    LocalMux I__4775 (
            .O(N__27397),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__4774 (
            .O(N__27394),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__4773 (
            .O(N__27389),
            .I(N__27386));
    InMux I__4772 (
            .O(N__27386),
            .I(N__27383));
    LocalMux I__4771 (
            .O(N__27383),
            .I(N__27380));
    Odrv12 I__4770 (
            .O(N__27380),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__4769 (
            .O(N__27377),
            .I(N__27373));
    InMux I__4768 (
            .O(N__27376),
            .I(N__27370));
    LocalMux I__4767 (
            .O(N__27373),
            .I(N__27367));
    LocalMux I__4766 (
            .O(N__27370),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__4765 (
            .O(N__27367),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__4764 (
            .O(N__27362),
            .I(N__27359));
    LocalMux I__4763 (
            .O(N__27359),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__4762 (
            .O(N__27356),
            .I(N__27353));
    InMux I__4761 (
            .O(N__27353),
            .I(N__27350));
    LocalMux I__4760 (
            .O(N__27350),
            .I(N__27347));
    Odrv4 I__4759 (
            .O(N__27347),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__4758 (
            .O(N__27344),
            .I(N__27341));
    LocalMux I__4757 (
            .O(N__27341),
            .I(N__27338));
    Span12Mux_h I__4756 (
            .O(N__27338),
            .I(N__27335));
    Odrv12 I__4755 (
            .O(N__27335),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    InMux I__4754 (
            .O(N__27332),
            .I(N__27329));
    LocalMux I__4753 (
            .O(N__27329),
            .I(N__27326));
    Span4Mux_h I__4752 (
            .O(N__27326),
            .I(N__27322));
    InMux I__4751 (
            .O(N__27325),
            .I(N__27319));
    Span4Mux_h I__4750 (
            .O(N__27322),
            .I(N__27316));
    LocalMux I__4749 (
            .O(N__27319),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__4748 (
            .O(N__27316),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__4747 (
            .O(N__27311),
            .I(N__27308));
    InMux I__4746 (
            .O(N__27308),
            .I(N__27305));
    LocalMux I__4745 (
            .O(N__27305),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__4744 (
            .O(N__27302),
            .I(N__27299));
    LocalMux I__4743 (
            .O(N__27299),
            .I(N__27296));
    Span4Mux_h I__4742 (
            .O(N__27296),
            .I(N__27293));
    Odrv4 I__4741 (
            .O(N__27293),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    InMux I__4740 (
            .O(N__27290),
            .I(N__27286));
    InMux I__4739 (
            .O(N__27289),
            .I(N__27283));
    LocalMux I__4738 (
            .O(N__27286),
            .I(N__27280));
    LocalMux I__4737 (
            .O(N__27283),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__4736 (
            .O(N__27280),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__4735 (
            .O(N__27275),
            .I(N__27272));
    InMux I__4734 (
            .O(N__27272),
            .I(N__27269));
    LocalMux I__4733 (
            .O(N__27269),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__4732 (
            .O(N__27266),
            .I(N__27263));
    LocalMux I__4731 (
            .O(N__27263),
            .I(N__27259));
    InMux I__4730 (
            .O(N__27262),
            .I(N__27256));
    Span4Mux_v I__4729 (
            .O(N__27259),
            .I(N__27253));
    LocalMux I__4728 (
            .O(N__27256),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__4727 (
            .O(N__27253),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__4726 (
            .O(N__27248),
            .I(N__27245));
    LocalMux I__4725 (
            .O(N__27245),
            .I(N__27242));
    Span4Mux_h I__4724 (
            .O(N__27242),
            .I(N__27239));
    Odrv4 I__4723 (
            .O(N__27239),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__4722 (
            .O(N__27236),
            .I(N__27233));
    InMux I__4721 (
            .O(N__27233),
            .I(N__27230));
    LocalMux I__4720 (
            .O(N__27230),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    InMux I__4719 (
            .O(N__27227),
            .I(N__27224));
    LocalMux I__4718 (
            .O(N__27224),
            .I(N__27221));
    Span4Mux_h I__4717 (
            .O(N__27221),
            .I(N__27218));
    Span4Mux_h I__4716 (
            .O(N__27218),
            .I(N__27215));
    Odrv4 I__4715 (
            .O(N__27215),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    InMux I__4714 (
            .O(N__27212),
            .I(N__27208));
    InMux I__4713 (
            .O(N__27211),
            .I(N__27205));
    LocalMux I__4712 (
            .O(N__27208),
            .I(N__27202));
    LocalMux I__4711 (
            .O(N__27205),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__4710 (
            .O(N__27202),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__4709 (
            .O(N__27197),
            .I(N__27194));
    InMux I__4708 (
            .O(N__27194),
            .I(N__27191));
    LocalMux I__4707 (
            .O(N__27191),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__4706 (
            .O(N__27188),
            .I(N__27184));
    InMux I__4705 (
            .O(N__27187),
            .I(N__27181));
    LocalMux I__4704 (
            .O(N__27184),
            .I(N__27178));
    LocalMux I__4703 (
            .O(N__27181),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__4702 (
            .O(N__27178),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__4701 (
            .O(N__27173),
            .I(N__27170));
    LocalMux I__4700 (
            .O(N__27170),
            .I(N__27167));
    Span4Mux_v I__4699 (
            .O(N__27167),
            .I(N__27164));
    Span4Mux_h I__4698 (
            .O(N__27164),
            .I(N__27161));
    Odrv4 I__4697 (
            .O(N__27161),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__4696 (
            .O(N__27158),
            .I(N__27155));
    InMux I__4695 (
            .O(N__27155),
            .I(N__27152));
    LocalMux I__4694 (
            .O(N__27152),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__4693 (
            .O(N__27149),
            .I(N__27146));
    LocalMux I__4692 (
            .O(N__27146),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__4691 (
            .O(N__27143),
            .I(N__27140));
    InMux I__4690 (
            .O(N__27140),
            .I(N__27137));
    LocalMux I__4689 (
            .O(N__27137),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__4688 (
            .O(N__27134),
            .I(N__27131));
    InMux I__4687 (
            .O(N__27131),
            .I(N__27128));
    LocalMux I__4686 (
            .O(N__27128),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    InMux I__4685 (
            .O(N__27125),
            .I(N__27121));
    InMux I__4684 (
            .O(N__27124),
            .I(N__27118));
    LocalMux I__4683 (
            .O(N__27121),
            .I(N__27115));
    LocalMux I__4682 (
            .O(N__27118),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__4681 (
            .O(N__27115),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__4680 (
            .O(N__27110),
            .I(N__27107));
    LocalMux I__4679 (
            .O(N__27107),
            .I(N__27104));
    Odrv4 I__4678 (
            .O(N__27104),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__4677 (
            .O(N__27101),
            .I(N__27097));
    InMux I__4676 (
            .O(N__27100),
            .I(N__27094));
    InMux I__4675 (
            .O(N__27097),
            .I(N__27091));
    LocalMux I__4674 (
            .O(N__27094),
            .I(N__27088));
    LocalMux I__4673 (
            .O(N__27091),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__4672 (
            .O(N__27088),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__4671 (
            .O(N__27083),
            .I(N__27080));
    InMux I__4670 (
            .O(N__27080),
            .I(N__27077));
    LocalMux I__4669 (
            .O(N__27077),
            .I(N__27074));
    Span4Mux_h I__4668 (
            .O(N__27074),
            .I(N__27071));
    Odrv4 I__4667 (
            .O(N__27071),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    InMux I__4666 (
            .O(N__27068),
            .I(N__27065));
    LocalMux I__4665 (
            .O(N__27065),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__4664 (
            .O(N__27062),
            .I(N__27059));
    LocalMux I__4663 (
            .O(N__27059),
            .I(N__27056));
    Span4Mux_h I__4662 (
            .O(N__27056),
            .I(N__27053));
    Odrv4 I__4661 (
            .O(N__27053),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    InMux I__4660 (
            .O(N__27050),
            .I(N__27046));
    InMux I__4659 (
            .O(N__27049),
            .I(N__27043));
    LocalMux I__4658 (
            .O(N__27046),
            .I(N__27040));
    LocalMux I__4657 (
            .O(N__27043),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__4656 (
            .O(N__27040),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__4655 (
            .O(N__27035),
            .I(N__27032));
    InMux I__4654 (
            .O(N__27032),
            .I(N__27029));
    LocalMux I__4653 (
            .O(N__27029),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__4652 (
            .O(N__27026),
            .I(N__27022));
    InMux I__4651 (
            .O(N__27025),
            .I(N__27019));
    LocalMux I__4650 (
            .O(N__27022),
            .I(N__27016));
    LocalMux I__4649 (
            .O(N__27019),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__4648 (
            .O(N__27016),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__4647 (
            .O(N__27011),
            .I(N__27008));
    LocalMux I__4646 (
            .O(N__27008),
            .I(N__27005));
    Span4Mux_h I__4645 (
            .O(N__27005),
            .I(N__27002));
    Odrv4 I__4644 (
            .O(N__27002),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__4643 (
            .O(N__26999),
            .I(N__26996));
    InMux I__4642 (
            .O(N__26996),
            .I(N__26993));
    LocalMux I__4641 (
            .O(N__26993),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__4640 (
            .O(N__26990),
            .I(N__26987));
    LocalMux I__4639 (
            .O(N__26987),
            .I(N__26984));
    Span4Mux_v I__4638 (
            .O(N__26984),
            .I(N__26981));
    Span4Mux_v I__4637 (
            .O(N__26981),
            .I(N__26978));
    Odrv4 I__4636 (
            .O(N__26978),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    InMux I__4635 (
            .O(N__26975),
            .I(N__26972));
    LocalMux I__4634 (
            .O(N__26972),
            .I(N__26969));
    Odrv4 I__4633 (
            .O(N__26969),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__4632 (
            .O(N__26966),
            .I(N__26963));
    LocalMux I__4631 (
            .O(N__26963),
            .I(N__26960));
    Span4Mux_v I__4630 (
            .O(N__26960),
            .I(N__26957));
    Span4Mux_v I__4629 (
            .O(N__26957),
            .I(N__26954));
    Odrv4 I__4628 (
            .O(N__26954),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    InMux I__4627 (
            .O(N__26951),
            .I(N__26948));
    LocalMux I__4626 (
            .O(N__26948),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__4625 (
            .O(N__26945),
            .I(N__26942));
    LocalMux I__4624 (
            .O(N__26942),
            .I(N__26939));
    Span4Mux_v I__4623 (
            .O(N__26939),
            .I(N__26936));
    Odrv4 I__4622 (
            .O(N__26936),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    InMux I__4621 (
            .O(N__26933),
            .I(N__26930));
    LocalMux I__4620 (
            .O(N__26930),
            .I(N__26927));
    Odrv4 I__4619 (
            .O(N__26927),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__4618 (
            .O(N__26924),
            .I(N__26921));
    LocalMux I__4617 (
            .O(N__26921),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHEZ0 ));
    InMux I__4616 (
            .O(N__26918),
            .I(N__26915));
    LocalMux I__4615 (
            .O(N__26915),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__4614 (
            .O(N__26912),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__4613 (
            .O(N__26909),
            .I(N__26906));
    LocalMux I__4612 (
            .O(N__26906),
            .I(N__26903));
    Span4Mux_h I__4611 (
            .O(N__26903),
            .I(N__26898));
    InMux I__4610 (
            .O(N__26902),
            .I(N__26893));
    InMux I__4609 (
            .O(N__26901),
            .I(N__26893));
    Odrv4 I__4608 (
            .O(N__26898),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    LocalMux I__4607 (
            .O(N__26893),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__4606 (
            .O(N__26888),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__4605 (
            .O(N__26885),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__4604 (
            .O(N__26882),
            .I(N__26879));
    LocalMux I__4603 (
            .O(N__26879),
            .I(N__26876));
    Span12Mux_v I__4602 (
            .O(N__26876),
            .I(N__26873));
    Odrv12 I__4601 (
            .O(N__26873),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__4600 (
            .O(N__26870),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__4599 (
            .O(N__26867),
            .I(bfn_12_12_0_));
    InMux I__4598 (
            .O(N__26864),
            .I(N__26861));
    LocalMux I__4597 (
            .O(N__26861),
            .I(N__26858));
    Span4Mux_v I__4596 (
            .O(N__26858),
            .I(N__26855));
    Span4Mux_v I__4595 (
            .O(N__26855),
            .I(N__26852));
    Odrv4 I__4594 (
            .O(N__26852),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__4593 (
            .O(N__26849),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__4592 (
            .O(N__26846),
            .I(N__26843));
    LocalMux I__4591 (
            .O(N__26843),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__4590 (
            .O(N__26840),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__4589 (
            .O(N__26837),
            .I(N__26834));
    LocalMux I__4588 (
            .O(N__26834),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__4587 (
            .O(N__26831),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__4586 (
            .O(N__26828),
            .I(N__26825));
    LocalMux I__4585 (
            .O(N__26825),
            .I(N__26821));
    InMux I__4584 (
            .O(N__26824),
            .I(N__26818));
    Span4Mux_h I__4583 (
            .O(N__26821),
            .I(N__26815));
    LocalMux I__4582 (
            .O(N__26818),
            .I(N__26812));
    Sp12to4 I__4581 (
            .O(N__26815),
            .I(N__26807));
    Span12Mux_v I__4580 (
            .O(N__26812),
            .I(N__26807));
    Odrv12 I__4579 (
            .O(N__26807),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    InMux I__4578 (
            .O(N__26804),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__4577 (
            .O(N__26801),
            .I(N__26798));
    LocalMux I__4576 (
            .O(N__26798),
            .I(N__26794));
    InMux I__4575 (
            .O(N__26797),
            .I(N__26791));
    Span4Mux_v I__4574 (
            .O(N__26794),
            .I(N__26788));
    LocalMux I__4573 (
            .O(N__26791),
            .I(N__26785));
    Span4Mux_v I__4572 (
            .O(N__26788),
            .I(N__26782));
    Odrv12 I__4571 (
            .O(N__26785),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    Odrv4 I__4570 (
            .O(N__26782),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    InMux I__4569 (
            .O(N__26777),
            .I(N__26774));
    LocalMux I__4568 (
            .O(N__26774),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__4567 (
            .O(N__26771),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__4566 (
            .O(N__26768),
            .I(N__26765));
    LocalMux I__4565 (
            .O(N__26765),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__4564 (
            .O(N__26762),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__4563 (
            .O(N__26759),
            .I(N__26756));
    LocalMux I__4562 (
            .O(N__26756),
            .I(N__26753));
    Span4Mux_v I__4561 (
            .O(N__26753),
            .I(N__26750));
    Odrv4 I__4560 (
            .O(N__26750),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__4559 (
            .O(N__26747),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    CascadeMux I__4558 (
            .O(N__26744),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_ ));
    InMux I__4557 (
            .O(N__26741),
            .I(N__26738));
    LocalMux I__4556 (
            .O(N__26738),
            .I(N__26735));
    Odrv4 I__4555 (
            .O(N__26735),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ));
    CascadeMux I__4554 (
            .O(N__26732),
            .I(\current_shift_inst.PI_CTRL.N_74_16_cascade_ ));
    InMux I__4553 (
            .O(N__26729),
            .I(N__26726));
    LocalMux I__4552 (
            .O(N__26726),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    InMux I__4551 (
            .O(N__26723),
            .I(N__26720));
    LocalMux I__4550 (
            .O(N__26720),
            .I(N__26716));
    InMux I__4549 (
            .O(N__26719),
            .I(N__26713));
    Span4Mux_s1_v I__4548 (
            .O(N__26716),
            .I(N__26708));
    LocalMux I__4547 (
            .O(N__26713),
            .I(N__26708));
    Span4Mux_v I__4546 (
            .O(N__26708),
            .I(N__26705));
    Span4Mux_h I__4545 (
            .O(N__26705),
            .I(N__26702));
    Sp12to4 I__4544 (
            .O(N__26702),
            .I(N__26697));
    InMux I__4543 (
            .O(N__26701),
            .I(N__26694));
    InMux I__4542 (
            .O(N__26700),
            .I(N__26691));
    Span12Mux_v I__4541 (
            .O(N__26697),
            .I(N__26688));
    LocalMux I__4540 (
            .O(N__26694),
            .I(N__26683));
    LocalMux I__4539 (
            .O(N__26691),
            .I(N__26683));
    Span12Mux_v I__4538 (
            .O(N__26688),
            .I(N__26680));
    Span12Mux_h I__4537 (
            .O(N__26683),
            .I(N__26677));
    Span12Mux_h I__4536 (
            .O(N__26680),
            .I(N__26674));
    Span12Mux_v I__4535 (
            .O(N__26677),
            .I(N__26671));
    Odrv12 I__4534 (
            .O(N__26674),
            .I(start_stop_c));
    Odrv12 I__4533 (
            .O(N__26671),
            .I(start_stop_c));
    InMux I__4532 (
            .O(N__26666),
            .I(N__26660));
    InMux I__4531 (
            .O(N__26665),
            .I(N__26657));
    InMux I__4530 (
            .O(N__26664),
            .I(N__26652));
    InMux I__4529 (
            .O(N__26663),
            .I(N__26652));
    LocalMux I__4528 (
            .O(N__26660),
            .I(N__26647));
    LocalMux I__4527 (
            .O(N__26657),
            .I(N__26642));
    LocalMux I__4526 (
            .O(N__26652),
            .I(N__26642));
    InMux I__4525 (
            .O(N__26651),
            .I(N__26639));
    InMux I__4524 (
            .O(N__26650),
            .I(N__26636));
    Odrv12 I__4523 (
            .O(N__26647),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__4522 (
            .O(N__26642),
            .I(phase_controller_inst1_state_4));
    LocalMux I__4521 (
            .O(N__26639),
            .I(phase_controller_inst1_state_4));
    LocalMux I__4520 (
            .O(N__26636),
            .I(phase_controller_inst1_state_4));
    InMux I__4519 (
            .O(N__26627),
            .I(N__26624));
    LocalMux I__4518 (
            .O(N__26624),
            .I(N__26619));
    InMux I__4517 (
            .O(N__26623),
            .I(N__26614));
    InMux I__4516 (
            .O(N__26622),
            .I(N__26614));
    Span4Mux_h I__4515 (
            .O(N__26619),
            .I(N__26611));
    LocalMux I__4514 (
            .O(N__26614),
            .I(N__26608));
    Odrv4 I__4513 (
            .O(N__26611),
            .I(il_min_comp2_D2));
    Odrv12 I__4512 (
            .O(N__26608),
            .I(il_min_comp2_D2));
    InMux I__4511 (
            .O(N__26603),
            .I(N__26599));
    InMux I__4510 (
            .O(N__26602),
            .I(N__26596));
    LocalMux I__4509 (
            .O(N__26599),
            .I(N__26593));
    LocalMux I__4508 (
            .O(N__26596),
            .I(N__26587));
    Span4Mux_s2_v I__4507 (
            .O(N__26593),
            .I(N__26584));
    CascadeMux I__4506 (
            .O(N__26592),
            .I(N__26581));
    InMux I__4505 (
            .O(N__26591),
            .I(N__26577));
    InMux I__4504 (
            .O(N__26590),
            .I(N__26574));
    Span4Mux_h I__4503 (
            .O(N__26587),
            .I(N__26569));
    Span4Mux_v I__4502 (
            .O(N__26584),
            .I(N__26569));
    InMux I__4501 (
            .O(N__26581),
            .I(N__26564));
    InMux I__4500 (
            .O(N__26580),
            .I(N__26564));
    LocalMux I__4499 (
            .O(N__26577),
            .I(N__26559));
    LocalMux I__4498 (
            .O(N__26574),
            .I(N__26559));
    Span4Mux_v I__4497 (
            .O(N__26569),
            .I(N__26556));
    LocalMux I__4496 (
            .O(N__26564),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__4495 (
            .O(N__26559),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__4494 (
            .O(N__26556),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    IoInMux I__4493 (
            .O(N__26549),
            .I(N__26546));
    LocalMux I__4492 (
            .O(N__26546),
            .I(N__26543));
    Span4Mux_s2_v I__4491 (
            .O(N__26543),
            .I(N__26540));
    Span4Mux_h I__4490 (
            .O(N__26540),
            .I(N__26537));
    Span4Mux_v I__4489 (
            .O(N__26537),
            .I(N__26533));
    InMux I__4488 (
            .O(N__26536),
            .I(N__26530));
    Odrv4 I__4487 (
            .O(N__26533),
            .I(T23_c));
    LocalMux I__4486 (
            .O(N__26530),
            .I(T23_c));
    InMux I__4485 (
            .O(N__26525),
            .I(N__26522));
    LocalMux I__4484 (
            .O(N__26522),
            .I(N__26519));
    Span4Mux_v I__4483 (
            .O(N__26519),
            .I(N__26516));
    Span4Mux_v I__4482 (
            .O(N__26516),
            .I(N__26513));
    Odrv4 I__4481 (
            .O(N__26513),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    InMux I__4480 (
            .O(N__26510),
            .I(\current_shift_inst.control_input_1_cry_3 ));
    InMux I__4479 (
            .O(N__26507),
            .I(\current_shift_inst.control_input_1_cry_4 ));
    InMux I__4478 (
            .O(N__26504),
            .I(\current_shift_inst.control_input_1_cry_5 ));
    InMux I__4477 (
            .O(N__26501),
            .I(N__26498));
    LocalMux I__4476 (
            .O(N__26498),
            .I(N__26495));
    Odrv12 I__4475 (
            .O(N__26495),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    InMux I__4474 (
            .O(N__26492),
            .I(\current_shift_inst.control_input_1_cry_6 ));
    InMux I__4473 (
            .O(N__26489),
            .I(bfn_11_22_0_));
    InMux I__4472 (
            .O(N__26486),
            .I(\current_shift_inst.control_input_1_cry_8 ));
    InMux I__4471 (
            .O(N__26483),
            .I(N__26480));
    LocalMux I__4470 (
            .O(N__26480),
            .I(N__26477));
    Span12Mux_v I__4469 (
            .O(N__26477),
            .I(N__26474));
    Odrv12 I__4468 (
            .O(N__26474),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    InMux I__4467 (
            .O(N__26471),
            .I(\current_shift_inst.control_input_1_cry_9 ));
    InMux I__4466 (
            .O(N__26468),
            .I(\current_shift_inst.control_input_1_cry_10 ));
    InMux I__4465 (
            .O(N__26465),
            .I(N__26462));
    LocalMux I__4464 (
            .O(N__26462),
            .I(\current_shift_inst.control_input_1_axb_10 ));
    InMux I__4463 (
            .O(N__26459),
            .I(N__26456));
    LocalMux I__4462 (
            .O(N__26456),
            .I(N__26453));
    Odrv4 I__4461 (
            .O(N__26453),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    CascadeMux I__4460 (
            .O(N__26450),
            .I(\phase_controller_inst2.start_timer_hc_RNOZ0Z_0_cascade_ ));
    InMux I__4459 (
            .O(N__26447),
            .I(N__26441));
    InMux I__4458 (
            .O(N__26446),
            .I(N__26434));
    InMux I__4457 (
            .O(N__26445),
            .I(N__26434));
    InMux I__4456 (
            .O(N__26444),
            .I(N__26434));
    LocalMux I__4455 (
            .O(N__26441),
            .I(\phase_controller_inst2.hc_time_passed ));
    LocalMux I__4454 (
            .O(N__26434),
            .I(\phase_controller_inst2.hc_time_passed ));
    CascadeMux I__4453 (
            .O(N__26429),
            .I(\phase_controller_inst2.start_timer_tr_0_sqmuxa_cascade_ ));
    InMux I__4452 (
            .O(N__26426),
            .I(\current_shift_inst.control_input_1_cry_0 ));
    InMux I__4451 (
            .O(N__26423),
            .I(N__26420));
    LocalMux I__4450 (
            .O(N__26420),
            .I(N__26417));
    Odrv12 I__4449 (
            .O(N__26417),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    InMux I__4448 (
            .O(N__26414),
            .I(\current_shift_inst.control_input_1_cry_1 ));
    InMux I__4447 (
            .O(N__26411),
            .I(N__26408));
    LocalMux I__4446 (
            .O(N__26408),
            .I(N__26405));
    Odrv4 I__4445 (
            .O(N__26405),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    InMux I__4444 (
            .O(N__26402),
            .I(\current_shift_inst.control_input_1_cry_2 ));
    InMux I__4443 (
            .O(N__26399),
            .I(N__26391));
    CascadeMux I__4442 (
            .O(N__26398),
            .I(N__26386));
    InMux I__4441 (
            .O(N__26397),
            .I(N__26383));
    CascadeMux I__4440 (
            .O(N__26396),
            .I(N__26378));
    CascadeMux I__4439 (
            .O(N__26395),
            .I(N__26375));
    CascadeMux I__4438 (
            .O(N__26394),
            .I(N__26370));
    LocalMux I__4437 (
            .O(N__26391),
            .I(N__26367));
    InMux I__4436 (
            .O(N__26390),
            .I(N__26364));
    InMux I__4435 (
            .O(N__26389),
            .I(N__26361));
    InMux I__4434 (
            .O(N__26386),
            .I(N__26358));
    LocalMux I__4433 (
            .O(N__26383),
            .I(N__26355));
    CascadeMux I__4432 (
            .O(N__26382),
            .I(N__26352));
    CascadeMux I__4431 (
            .O(N__26381),
            .I(N__26349));
    InMux I__4430 (
            .O(N__26378),
            .I(N__26345));
    InMux I__4429 (
            .O(N__26375),
            .I(N__26342));
    CascadeMux I__4428 (
            .O(N__26374),
            .I(N__26335));
    CascadeMux I__4427 (
            .O(N__26373),
            .I(N__26328));
    InMux I__4426 (
            .O(N__26370),
            .I(N__26325));
    Span4Mux_h I__4425 (
            .O(N__26367),
            .I(N__26322));
    LocalMux I__4424 (
            .O(N__26364),
            .I(N__26317));
    LocalMux I__4423 (
            .O(N__26361),
            .I(N__26317));
    LocalMux I__4422 (
            .O(N__26358),
            .I(N__26314));
    Span4Mux_h I__4421 (
            .O(N__26355),
            .I(N__26311));
    InMux I__4420 (
            .O(N__26352),
            .I(N__26304));
    InMux I__4419 (
            .O(N__26349),
            .I(N__26304));
    InMux I__4418 (
            .O(N__26348),
            .I(N__26304));
    LocalMux I__4417 (
            .O(N__26345),
            .I(N__26299));
    LocalMux I__4416 (
            .O(N__26342),
            .I(N__26299));
    InMux I__4415 (
            .O(N__26341),
            .I(N__26290));
    InMux I__4414 (
            .O(N__26340),
            .I(N__26290));
    InMux I__4413 (
            .O(N__26339),
            .I(N__26290));
    InMux I__4412 (
            .O(N__26338),
            .I(N__26290));
    InMux I__4411 (
            .O(N__26335),
            .I(N__26283));
    InMux I__4410 (
            .O(N__26334),
            .I(N__26283));
    InMux I__4409 (
            .O(N__26333),
            .I(N__26283));
    InMux I__4408 (
            .O(N__26332),
            .I(N__26276));
    InMux I__4407 (
            .O(N__26331),
            .I(N__26276));
    InMux I__4406 (
            .O(N__26328),
            .I(N__26276));
    LocalMux I__4405 (
            .O(N__26325),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    Odrv4 I__4404 (
            .O(N__26322),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    Odrv12 I__4403 (
            .O(N__26317),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    Odrv4 I__4402 (
            .O(N__26314),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    Odrv4 I__4401 (
            .O(N__26311),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__4400 (
            .O(N__26304),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    Odrv4 I__4399 (
            .O(N__26299),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__4398 (
            .O(N__26290),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__4397 (
            .O(N__26283),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__4396 (
            .O(N__26276),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    CascadeMux I__4395 (
            .O(N__26255),
            .I(N__26252));
    InMux I__4394 (
            .O(N__26252),
            .I(N__26249));
    LocalMux I__4393 (
            .O(N__26249),
            .I(N__26245));
    InMux I__4392 (
            .O(N__26248),
            .I(N__26241));
    Span4Mux_v I__4391 (
            .O(N__26245),
            .I(N__26238));
    InMux I__4390 (
            .O(N__26244),
            .I(N__26235));
    LocalMux I__4389 (
            .O(N__26241),
            .I(N__26232));
    Odrv4 I__4388 (
            .O(N__26238),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__4387 (
            .O(N__26235),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    Odrv4 I__4386 (
            .O(N__26232),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__4385 (
            .O(N__26225),
            .I(N__26221));
    InMux I__4384 (
            .O(N__26224),
            .I(N__26218));
    LocalMux I__4383 (
            .O(N__26221),
            .I(elapsed_time_ns_1_RNI81DJ11_0_2));
    LocalMux I__4382 (
            .O(N__26218),
            .I(elapsed_time_ns_1_RNI81DJ11_0_2));
    CascadeMux I__4381 (
            .O(N__26213),
            .I(elapsed_time_ns_1_RNI81DJ11_0_2_cascade_));
    InMux I__4380 (
            .O(N__26210),
            .I(N__26206));
    InMux I__4379 (
            .O(N__26209),
            .I(N__26201));
    LocalMux I__4378 (
            .O(N__26206),
            .I(N__26197));
    InMux I__4377 (
            .O(N__26205),
            .I(N__26194));
    InMux I__4376 (
            .O(N__26204),
            .I(N__26191));
    LocalMux I__4375 (
            .O(N__26201),
            .I(N__26188));
    InMux I__4374 (
            .O(N__26200),
            .I(N__26185));
    Span4Mux_v I__4373 (
            .O(N__26197),
            .I(N__26180));
    LocalMux I__4372 (
            .O(N__26194),
            .I(N__26180));
    LocalMux I__4371 (
            .O(N__26191),
            .I(elapsed_time_ns_1_RNIQURR91_0_3));
    Odrv4 I__4370 (
            .O(N__26188),
            .I(elapsed_time_ns_1_RNIQURR91_0_3));
    LocalMux I__4369 (
            .O(N__26185),
            .I(elapsed_time_ns_1_RNIQURR91_0_3));
    Odrv4 I__4368 (
            .O(N__26180),
            .I(elapsed_time_ns_1_RNIQURR91_0_3));
    InMux I__4367 (
            .O(N__26171),
            .I(N__26168));
    LocalMux I__4366 (
            .O(N__26168),
            .I(\phase_controller_inst1.stoper_hc.N_283 ));
    CascadeMux I__4365 (
            .O(N__26165),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_ ));
    InMux I__4364 (
            .O(N__26162),
            .I(N__26159));
    LocalMux I__4363 (
            .O(N__26159),
            .I(N__26155));
    InMux I__4362 (
            .O(N__26158),
            .I(N__26152));
    Odrv4 I__4361 (
            .O(N__26155),
            .I(\phase_controller_inst1.N_56 ));
    LocalMux I__4360 (
            .O(N__26152),
            .I(\phase_controller_inst1.N_56 ));
    CascadeMux I__4359 (
            .O(N__26147),
            .I(N__26144));
    InMux I__4358 (
            .O(N__26144),
            .I(N__26138));
    InMux I__4357 (
            .O(N__26143),
            .I(N__26138));
    LocalMux I__4356 (
            .O(N__26138),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__4355 (
            .O(N__26135),
            .I(N__26132));
    LocalMux I__4354 (
            .O(N__26132),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    CascadeMux I__4353 (
            .O(N__26129),
            .I(N__26126));
    InMux I__4352 (
            .O(N__26126),
            .I(N__26122));
    CascadeMux I__4351 (
            .O(N__26125),
            .I(N__26117));
    LocalMux I__4350 (
            .O(N__26122),
            .I(N__26114));
    CascadeMux I__4349 (
            .O(N__26121),
            .I(N__26111));
    InMux I__4348 (
            .O(N__26120),
            .I(N__26108));
    InMux I__4347 (
            .O(N__26117),
            .I(N__26105));
    Span4Mux_h I__4346 (
            .O(N__26114),
            .I(N__26102));
    InMux I__4345 (
            .O(N__26111),
            .I(N__26099));
    LocalMux I__4344 (
            .O(N__26108),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    LocalMux I__4343 (
            .O(N__26105),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    Odrv4 I__4342 (
            .O(N__26102),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    LocalMux I__4341 (
            .O(N__26099),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    InMux I__4340 (
            .O(N__26090),
            .I(N__26087));
    LocalMux I__4339 (
            .O(N__26087),
            .I(N__26084));
    Span4Mux_h I__4338 (
            .O(N__26084),
            .I(N__26081));
    Odrv4 I__4337 (
            .O(N__26081),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__4336 (
            .O(N__26078),
            .I(N__26073));
    CascadeMux I__4335 (
            .O(N__26077),
            .I(N__26069));
    InMux I__4334 (
            .O(N__26076),
            .I(N__26066));
    InMux I__4333 (
            .O(N__26073),
            .I(N__26063));
    InMux I__4332 (
            .O(N__26072),
            .I(N__26058));
    InMux I__4331 (
            .O(N__26069),
            .I(N__26058));
    LocalMux I__4330 (
            .O(N__26066),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    LocalMux I__4329 (
            .O(N__26063),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    LocalMux I__4328 (
            .O(N__26058),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    InMux I__4327 (
            .O(N__26051),
            .I(N__26048));
    LocalMux I__4326 (
            .O(N__26048),
            .I(N__26045));
    Span4Mux_v I__4325 (
            .O(N__26045),
            .I(N__26042));
    Odrv4 I__4324 (
            .O(N__26042),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    InMux I__4323 (
            .O(N__26039),
            .I(N__26026));
    InMux I__4322 (
            .O(N__26038),
            .I(N__26023));
    CascadeMux I__4321 (
            .O(N__26037),
            .I(N__26019));
    CascadeMux I__4320 (
            .O(N__26036),
            .I(N__26016));
    CascadeMux I__4319 (
            .O(N__26035),
            .I(N__26012));
    CascadeMux I__4318 (
            .O(N__26034),
            .I(N__26005));
    CascadeMux I__4317 (
            .O(N__26033),
            .I(N__26000));
    InMux I__4316 (
            .O(N__26032),
            .I(N__25987));
    InMux I__4315 (
            .O(N__26031),
            .I(N__25987));
    InMux I__4314 (
            .O(N__26030),
            .I(N__25987));
    InMux I__4313 (
            .O(N__26029),
            .I(N__25987));
    LocalMux I__4312 (
            .O(N__26026),
            .I(N__25982));
    LocalMux I__4311 (
            .O(N__26023),
            .I(N__25982));
    CascadeMux I__4310 (
            .O(N__26022),
            .I(N__25978));
    InMux I__4309 (
            .O(N__26019),
            .I(N__25961));
    InMux I__4308 (
            .O(N__26016),
            .I(N__25961));
    InMux I__4307 (
            .O(N__26015),
            .I(N__25961));
    InMux I__4306 (
            .O(N__26012),
            .I(N__25961));
    InMux I__4305 (
            .O(N__26011),
            .I(N__25961));
    InMux I__4304 (
            .O(N__26010),
            .I(N__25961));
    InMux I__4303 (
            .O(N__26009),
            .I(N__25961));
    InMux I__4302 (
            .O(N__26008),
            .I(N__25961));
    InMux I__4301 (
            .O(N__26005),
            .I(N__25944));
    InMux I__4300 (
            .O(N__26004),
            .I(N__25944));
    InMux I__4299 (
            .O(N__26003),
            .I(N__25944));
    InMux I__4298 (
            .O(N__26000),
            .I(N__25944));
    InMux I__4297 (
            .O(N__25999),
            .I(N__25944));
    InMux I__4296 (
            .O(N__25998),
            .I(N__25944));
    InMux I__4295 (
            .O(N__25997),
            .I(N__25944));
    InMux I__4294 (
            .O(N__25996),
            .I(N__25944));
    LocalMux I__4293 (
            .O(N__25987),
            .I(N__25941));
    Span4Mux_v I__4292 (
            .O(N__25982),
            .I(N__25926));
    InMux I__4291 (
            .O(N__25981),
            .I(N__25921));
    InMux I__4290 (
            .O(N__25978),
            .I(N__25921));
    LocalMux I__4289 (
            .O(N__25961),
            .I(N__25918));
    LocalMux I__4288 (
            .O(N__25944),
            .I(N__25915));
    Span4Mux_h I__4287 (
            .O(N__25941),
            .I(N__25912));
    InMux I__4286 (
            .O(N__25940),
            .I(N__25906));
    InMux I__4285 (
            .O(N__25939),
            .I(N__25906));
    InMux I__4284 (
            .O(N__25938),
            .I(N__25893));
    InMux I__4283 (
            .O(N__25937),
            .I(N__25893));
    InMux I__4282 (
            .O(N__25936),
            .I(N__25893));
    InMux I__4281 (
            .O(N__25935),
            .I(N__25893));
    InMux I__4280 (
            .O(N__25934),
            .I(N__25893));
    InMux I__4279 (
            .O(N__25933),
            .I(N__25893));
    InMux I__4278 (
            .O(N__25932),
            .I(N__25884));
    InMux I__4277 (
            .O(N__25931),
            .I(N__25884));
    InMux I__4276 (
            .O(N__25930),
            .I(N__25884));
    InMux I__4275 (
            .O(N__25929),
            .I(N__25884));
    Span4Mux_h I__4274 (
            .O(N__25926),
            .I(N__25881));
    LocalMux I__4273 (
            .O(N__25921),
            .I(N__25876));
    Span4Mux_v I__4272 (
            .O(N__25918),
            .I(N__25876));
    Span4Mux_h I__4271 (
            .O(N__25915),
            .I(N__25873));
    Span4Mux_h I__4270 (
            .O(N__25912),
            .I(N__25870));
    InMux I__4269 (
            .O(N__25911),
            .I(N__25867));
    LocalMux I__4268 (
            .O(N__25906),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    LocalMux I__4267 (
            .O(N__25893),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    LocalMux I__4266 (
            .O(N__25884),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    Odrv4 I__4265 (
            .O(N__25881),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    Odrv4 I__4264 (
            .O(N__25876),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    Odrv4 I__4263 (
            .O(N__25873),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    Odrv4 I__4262 (
            .O(N__25870),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    LocalMux I__4261 (
            .O(N__25867),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    InMux I__4260 (
            .O(N__25850),
            .I(N__25847));
    LocalMux I__4259 (
            .O(N__25847),
            .I(N__25842));
    InMux I__4258 (
            .O(N__25846),
            .I(N__25839));
    InMux I__4257 (
            .O(N__25845),
            .I(N__25836));
    Odrv4 I__4256 (
            .O(N__25842),
            .I(elapsed_time_ns_1_RNIDP2KD1_0_1));
    LocalMux I__4255 (
            .O(N__25839),
            .I(elapsed_time_ns_1_RNIDP2KD1_0_1));
    LocalMux I__4254 (
            .O(N__25836),
            .I(elapsed_time_ns_1_RNIDP2KD1_0_1));
    InMux I__4253 (
            .O(N__25829),
            .I(N__25825));
    InMux I__4252 (
            .O(N__25828),
            .I(N__25822));
    LocalMux I__4251 (
            .O(N__25825),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_0_1Z0Z_1 ));
    LocalMux I__4250 (
            .O(N__25822),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_0_1Z0Z_1 ));
    InMux I__4249 (
            .O(N__25817),
            .I(N__25814));
    LocalMux I__4248 (
            .O(N__25814),
            .I(N__25811));
    Span4Mux_h I__4247 (
            .O(N__25811),
            .I(N__25808));
    Odrv4 I__4246 (
            .O(N__25808),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__4245 (
            .O(N__25805),
            .I(N__25801));
    CascadeMux I__4244 (
            .O(N__25804),
            .I(N__25793));
    LocalMux I__4243 (
            .O(N__25801),
            .I(N__25782));
    InMux I__4242 (
            .O(N__25800),
            .I(N__25777));
    InMux I__4241 (
            .O(N__25799),
            .I(N__25777));
    InMux I__4240 (
            .O(N__25798),
            .I(N__25766));
    InMux I__4239 (
            .O(N__25797),
            .I(N__25766));
    InMux I__4238 (
            .O(N__25796),
            .I(N__25766));
    InMux I__4237 (
            .O(N__25793),
            .I(N__25766));
    InMux I__4236 (
            .O(N__25792),
            .I(N__25766));
    InMux I__4235 (
            .O(N__25791),
            .I(N__25761));
    InMux I__4234 (
            .O(N__25790),
            .I(N__25761));
    InMux I__4233 (
            .O(N__25789),
            .I(N__25752));
    InMux I__4232 (
            .O(N__25788),
            .I(N__25752));
    InMux I__4231 (
            .O(N__25787),
            .I(N__25752));
    InMux I__4230 (
            .O(N__25786),
            .I(N__25752));
    InMux I__4229 (
            .O(N__25785),
            .I(N__25749));
    Span4Mux_h I__4228 (
            .O(N__25782),
            .I(N__25746));
    LocalMux I__4227 (
            .O(N__25777),
            .I(\phase_controller_inst1.stoper_hc.N_325 ));
    LocalMux I__4226 (
            .O(N__25766),
            .I(\phase_controller_inst1.stoper_hc.N_325 ));
    LocalMux I__4225 (
            .O(N__25761),
            .I(\phase_controller_inst1.stoper_hc.N_325 ));
    LocalMux I__4224 (
            .O(N__25752),
            .I(\phase_controller_inst1.stoper_hc.N_325 ));
    LocalMux I__4223 (
            .O(N__25749),
            .I(\phase_controller_inst1.stoper_hc.N_325 ));
    Odrv4 I__4222 (
            .O(N__25746),
            .I(\phase_controller_inst1.stoper_hc.N_325 ));
    CascadeMux I__4221 (
            .O(N__25733),
            .I(N__25725));
    CascadeMux I__4220 (
            .O(N__25732),
            .I(N__25722));
    CascadeMux I__4219 (
            .O(N__25731),
            .I(N__25716));
    InMux I__4218 (
            .O(N__25730),
            .I(N__25711));
    InMux I__4217 (
            .O(N__25729),
            .I(N__25706));
    InMux I__4216 (
            .O(N__25728),
            .I(N__25706));
    InMux I__4215 (
            .O(N__25725),
            .I(N__25703));
    InMux I__4214 (
            .O(N__25722),
            .I(N__25700));
    InMux I__4213 (
            .O(N__25721),
            .I(N__25689));
    InMux I__4212 (
            .O(N__25720),
            .I(N__25689));
    InMux I__4211 (
            .O(N__25719),
            .I(N__25689));
    InMux I__4210 (
            .O(N__25716),
            .I(N__25689));
    InMux I__4209 (
            .O(N__25715),
            .I(N__25689));
    InMux I__4208 (
            .O(N__25714),
            .I(N__25686));
    LocalMux I__4207 (
            .O(N__25711),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__4206 (
            .O(N__25706),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__4205 (
            .O(N__25703),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__4204 (
            .O(N__25700),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__4203 (
            .O(N__25689),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__4202 (
            .O(N__25686),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    InMux I__4201 (
            .O(N__25673),
            .I(N__25669));
    InMux I__4200 (
            .O(N__25672),
            .I(N__25666));
    LocalMux I__4199 (
            .O(N__25669),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_0_0Z0Z_3 ));
    LocalMux I__4198 (
            .O(N__25666),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_0_0Z0Z_3 ));
    InMux I__4197 (
            .O(N__25661),
            .I(N__25658));
    LocalMux I__4196 (
            .O(N__25658),
            .I(N__25655));
    Span4Mux_v I__4195 (
            .O(N__25655),
            .I(N__25652));
    Odrv4 I__4194 (
            .O(N__25652),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    CEMux I__4193 (
            .O(N__25649),
            .I(N__25646));
    LocalMux I__4192 (
            .O(N__25646),
            .I(N__25643));
    Span4Mux_v I__4191 (
            .O(N__25643),
            .I(N__25638));
    CEMux I__4190 (
            .O(N__25642),
            .I(N__25635));
    CEMux I__4189 (
            .O(N__25641),
            .I(N__25632));
    Span4Mux_v I__4188 (
            .O(N__25638),
            .I(N__25629));
    LocalMux I__4187 (
            .O(N__25635),
            .I(N__25626));
    LocalMux I__4186 (
            .O(N__25632),
            .I(N__25623));
    Span4Mux_h I__4185 (
            .O(N__25629),
            .I(N__25618));
    Span4Mux_v I__4184 (
            .O(N__25626),
            .I(N__25618));
    Span12Mux_s10_h I__4183 (
            .O(N__25623),
            .I(N__25615));
    Span4Mux_h I__4182 (
            .O(N__25618),
            .I(N__25612));
    Odrv12 I__4181 (
            .O(N__25615),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa_0 ));
    Odrv4 I__4180 (
            .O(N__25612),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa_0 ));
    CEMux I__4179 (
            .O(N__25607),
            .I(N__25603));
    CEMux I__4178 (
            .O(N__25606),
            .I(N__25600));
    LocalMux I__4177 (
            .O(N__25603),
            .I(N__25597));
    LocalMux I__4176 (
            .O(N__25600),
            .I(N__25592));
    Span4Mux_v I__4175 (
            .O(N__25597),
            .I(N__25589));
    CEMux I__4174 (
            .O(N__25596),
            .I(N__25586));
    CEMux I__4173 (
            .O(N__25595),
            .I(N__25583));
    Span4Mux_v I__4172 (
            .O(N__25592),
            .I(N__25576));
    Span4Mux_h I__4171 (
            .O(N__25589),
            .I(N__25576));
    LocalMux I__4170 (
            .O(N__25586),
            .I(N__25576));
    LocalMux I__4169 (
            .O(N__25583),
            .I(N__25573));
    Span4Mux_h I__4168 (
            .O(N__25576),
            .I(N__25570));
    Span4Mux_h I__4167 (
            .O(N__25573),
            .I(N__25567));
    Odrv4 I__4166 (
            .O(N__25570),
            .I(\delay_measurement_inst.delay_hc_timer.N_433_i ));
    Odrv4 I__4165 (
            .O(N__25567),
            .I(\delay_measurement_inst.delay_hc_timer.N_433_i ));
    CascadeMux I__4164 (
            .O(N__25562),
            .I(N__25559));
    InMux I__4163 (
            .O(N__25559),
            .I(N__25556));
    LocalMux I__4162 (
            .O(N__25556),
            .I(N__25553));
    Span4Mux_v I__4161 (
            .O(N__25553),
            .I(N__25550));
    Odrv4 I__4160 (
            .O(N__25550),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    CascadeMux I__4159 (
            .O(N__25547),
            .I(N__25544));
    InMux I__4158 (
            .O(N__25544),
            .I(N__25541));
    LocalMux I__4157 (
            .O(N__25541),
            .I(N__25538));
    Span4Mux_h I__4156 (
            .O(N__25538),
            .I(N__25533));
    InMux I__4155 (
            .O(N__25537),
            .I(N__25528));
    InMux I__4154 (
            .O(N__25536),
            .I(N__25528));
    Odrv4 I__4153 (
            .O(N__25533),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    LocalMux I__4152 (
            .O(N__25528),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__4151 (
            .O(N__25523),
            .I(N__25520));
    LocalMux I__4150 (
            .O(N__25520),
            .I(N__25516));
    InMux I__4149 (
            .O(N__25519),
            .I(N__25512));
    Span4Mux_h I__4148 (
            .O(N__25516),
            .I(N__25509));
    InMux I__4147 (
            .O(N__25515),
            .I(N__25506));
    LocalMux I__4146 (
            .O(N__25512),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7));
    Odrv4 I__4145 (
            .O(N__25509),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7));
    LocalMux I__4144 (
            .O(N__25506),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7));
    CascadeMux I__4143 (
            .O(N__25499),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7_cascade_));
    CascadeMux I__4142 (
            .O(N__25496),
            .I(N__25493));
    InMux I__4141 (
            .O(N__25493),
            .I(N__25490));
    LocalMux I__4140 (
            .O(N__25490),
            .I(N__25487));
    Span4Mux_h I__4139 (
            .O(N__25487),
            .I(N__25483));
    InMux I__4138 (
            .O(N__25486),
            .I(N__25480));
    Odrv4 I__4137 (
            .O(N__25483),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__4136 (
            .O(N__25480),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    CascadeMux I__4135 (
            .O(N__25475),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ));
    InMux I__4134 (
            .O(N__25472),
            .I(N__25469));
    LocalMux I__4133 (
            .O(N__25469),
            .I(N__25465));
    InMux I__4132 (
            .O(N__25468),
            .I(N__25460));
    Span4Mux_h I__4131 (
            .O(N__25465),
            .I(N__25457));
    InMux I__4130 (
            .O(N__25464),
            .I(N__25454));
    InMux I__4129 (
            .O(N__25463),
            .I(N__25451));
    LocalMux I__4128 (
            .O(N__25460),
            .I(N__25445));
    Span4Mux_h I__4127 (
            .O(N__25457),
            .I(N__25442));
    LocalMux I__4126 (
            .O(N__25454),
            .I(N__25437));
    LocalMux I__4125 (
            .O(N__25451),
            .I(N__25437));
    InMux I__4124 (
            .O(N__25450),
            .I(N__25432));
    InMux I__4123 (
            .O(N__25449),
            .I(N__25432));
    InMux I__4122 (
            .O(N__25448),
            .I(N__25429));
    Odrv4 I__4121 (
            .O(N__25445),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    Odrv4 I__4120 (
            .O(N__25442),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    Odrv4 I__4119 (
            .O(N__25437),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    LocalMux I__4118 (
            .O(N__25432),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    LocalMux I__4117 (
            .O(N__25429),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    CascadeMux I__4116 (
            .O(N__25418),
            .I(elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_));
    InMux I__4115 (
            .O(N__25415),
            .I(N__25412));
    LocalMux I__4114 (
            .O(N__25412),
            .I(N__25409));
    Span4Mux_v I__4113 (
            .O(N__25409),
            .I(N__25406));
    Odrv4 I__4112 (
            .O(N__25406),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__4111 (
            .O(N__25403),
            .I(N__25399));
    InMux I__4110 (
            .O(N__25402),
            .I(N__25396));
    InMux I__4109 (
            .O(N__25399),
            .I(N__25393));
    LocalMux I__4108 (
            .O(N__25396),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_0Z0Z_2 ));
    LocalMux I__4107 (
            .O(N__25393),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_0Z0Z_2 ));
    InMux I__4106 (
            .O(N__25388),
            .I(N__25385));
    LocalMux I__4105 (
            .O(N__25385),
            .I(N__25382));
    Span4Mux_h I__4104 (
            .O(N__25382),
            .I(N__25379));
    Odrv4 I__4103 (
            .O(N__25379),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__4102 (
            .O(N__25376),
            .I(N__25373));
    InMux I__4101 (
            .O(N__25373),
            .I(N__25369));
    CascadeMux I__4100 (
            .O(N__25372),
            .I(N__25365));
    LocalMux I__4099 (
            .O(N__25369),
            .I(N__25362));
    InMux I__4098 (
            .O(N__25368),
            .I(N__25358));
    InMux I__4097 (
            .O(N__25365),
            .I(N__25355));
    Span4Mux_h I__4096 (
            .O(N__25362),
            .I(N__25352));
    InMux I__4095 (
            .O(N__25361),
            .I(N__25349));
    LocalMux I__4094 (
            .O(N__25358),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4));
    LocalMux I__4093 (
            .O(N__25355),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4));
    Odrv4 I__4092 (
            .O(N__25352),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4));
    LocalMux I__4091 (
            .O(N__25349),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4));
    InMux I__4090 (
            .O(N__25340),
            .I(N__25337));
    LocalMux I__4089 (
            .O(N__25337),
            .I(N__25334));
    Span4Mux_h I__4088 (
            .O(N__25334),
            .I(N__25331));
    Span4Mux_h I__4087 (
            .O(N__25331),
            .I(N__25328));
    Odrv4 I__4086 (
            .O(N__25328),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__4085 (
            .O(N__25325),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__4084 (
            .O(N__25322),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__4083 (
            .O(N__25319),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__4082 (
            .O(N__25316),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__4081 (
            .O(N__25313),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__4080 (
            .O(N__25310),
            .I(bfn_11_15_0_));
    InMux I__4079 (
            .O(N__25307),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__4078 (
            .O(N__25304),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__4077 (
            .O(N__25301),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__4076 (
            .O(N__25298),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__4075 (
            .O(N__25295),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__4074 (
            .O(N__25292),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__4073 (
            .O(N__25289),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__4072 (
            .O(N__25286),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__4071 (
            .O(N__25283),
            .I(bfn_11_14_0_));
    InMux I__4070 (
            .O(N__25280),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__4069 (
            .O(N__25277),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__4068 (
            .O(N__25274),
            .I(N__25271));
    LocalMux I__4067 (
            .O(N__25271),
            .I(N__25268));
    Odrv4 I__4066 (
            .O(N__25268),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    InMux I__4065 (
            .O(N__25265),
            .I(N__25262));
    LocalMux I__4064 (
            .O(N__25262),
            .I(N__25259));
    Odrv12 I__4063 (
            .O(N__25259),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__4062 (
            .O(N__25256),
            .I(N__25252));
    InMux I__4061 (
            .O(N__25255),
            .I(N__25249));
    LocalMux I__4060 (
            .O(N__25252),
            .I(N__25245));
    LocalMux I__4059 (
            .O(N__25249),
            .I(N__25241));
    CascadeMux I__4058 (
            .O(N__25248),
            .I(N__25236));
    Span4Mux_h I__4057 (
            .O(N__25245),
            .I(N__25231));
    InMux I__4056 (
            .O(N__25244),
            .I(N__25228));
    Span4Mux_v I__4055 (
            .O(N__25241),
            .I(N__25225));
    InMux I__4054 (
            .O(N__25240),
            .I(N__25214));
    InMux I__4053 (
            .O(N__25239),
            .I(N__25214));
    InMux I__4052 (
            .O(N__25236),
            .I(N__25214));
    InMux I__4051 (
            .O(N__25235),
            .I(N__25214));
    InMux I__4050 (
            .O(N__25234),
            .I(N__25214));
    Span4Mux_v I__4049 (
            .O(N__25231),
            .I(N__25211));
    LocalMux I__4048 (
            .O(N__25228),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__4047 (
            .O(N__25225),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__4046 (
            .O(N__25214),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__4045 (
            .O(N__25211),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    InMux I__4044 (
            .O(N__25202),
            .I(N__25196));
    InMux I__4043 (
            .O(N__25201),
            .I(N__25191));
    InMux I__4042 (
            .O(N__25200),
            .I(N__25188));
    InMux I__4041 (
            .O(N__25199),
            .I(N__25185));
    LocalMux I__4040 (
            .O(N__25196),
            .I(N__25182));
    InMux I__4039 (
            .O(N__25195),
            .I(N__25177));
    InMux I__4038 (
            .O(N__25194),
            .I(N__25177));
    LocalMux I__4037 (
            .O(N__25191),
            .I(N__25174));
    LocalMux I__4036 (
            .O(N__25188),
            .I(N__25171));
    LocalMux I__4035 (
            .O(N__25185),
            .I(N__25164));
    Span4Mux_h I__4034 (
            .O(N__25182),
            .I(N__25164));
    LocalMux I__4033 (
            .O(N__25177),
            .I(N__25164));
    Odrv4 I__4032 (
            .O(N__25174),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__4031 (
            .O(N__25171),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__4030 (
            .O(N__25164),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__4029 (
            .O(N__25157),
            .I(N__25154));
    InMux I__4028 (
            .O(N__25154),
            .I(N__25151));
    LocalMux I__4027 (
            .O(N__25151),
            .I(N__25147));
    InMux I__4026 (
            .O(N__25150),
            .I(N__25143));
    Span4Mux_h I__4025 (
            .O(N__25147),
            .I(N__25140));
    InMux I__4024 (
            .O(N__25146),
            .I(N__25137));
    LocalMux I__4023 (
            .O(N__25143),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__4022 (
            .O(N__25140),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__4021 (
            .O(N__25137),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    SRMux I__4020 (
            .O(N__25130),
            .I(N__25127));
    LocalMux I__4019 (
            .O(N__25127),
            .I(N__25122));
    SRMux I__4018 (
            .O(N__25126),
            .I(N__25119));
    SRMux I__4017 (
            .O(N__25125),
            .I(N__25115));
    Span4Mux_h I__4016 (
            .O(N__25122),
            .I(N__25110));
    LocalMux I__4015 (
            .O(N__25119),
            .I(N__25110));
    SRMux I__4014 (
            .O(N__25118),
            .I(N__25107));
    LocalMux I__4013 (
            .O(N__25115),
            .I(N__25104));
    Span4Mux_v I__4012 (
            .O(N__25110),
            .I(N__25101));
    LocalMux I__4011 (
            .O(N__25107),
            .I(N__25098));
    Span4Mux_h I__4010 (
            .O(N__25104),
            .I(N__25095));
    Span4Mux_h I__4009 (
            .O(N__25101),
            .I(N__25090));
    Span4Mux_v I__4008 (
            .O(N__25098),
            .I(N__25090));
    Sp12to4 I__4007 (
            .O(N__25095),
            .I(N__25087));
    Span4Mux_h I__4006 (
            .O(N__25090),
            .I(N__25084));
    Odrv12 I__4005 (
            .O(N__25087),
            .I(\phase_controller_inst1.stoper_hc.un1_stoper_state12_1_0_i ));
    Odrv4 I__4004 (
            .O(N__25084),
            .I(\phase_controller_inst1.stoper_hc.un1_stoper_state12_1_0_i ));
    InMux I__4003 (
            .O(N__25079),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ));
    IoInMux I__4002 (
            .O(N__25076),
            .I(N__25073));
    LocalMux I__4001 (
            .O(N__25073),
            .I(N__25070));
    Span4Mux_s3_v I__4000 (
            .O(N__25070),
            .I(N__25067));
    Sp12to4 I__3999 (
            .O(N__25067),
            .I(N__25064));
    Span12Mux_h I__3998 (
            .O(N__25064),
            .I(N__25060));
    InMux I__3997 (
            .O(N__25063),
            .I(N__25057));
    Odrv12 I__3996 (
            .O(N__25060),
            .I(T12_c));
    LocalMux I__3995 (
            .O(N__25057),
            .I(T12_c));
    InMux I__3994 (
            .O(N__25052),
            .I(N__25046));
    InMux I__3993 (
            .O(N__25051),
            .I(N__25046));
    LocalMux I__3992 (
            .O(N__25046),
            .I(state_ns_i_a3_1));
    ClkMux I__3991 (
            .O(N__25043),
            .I(N__25037));
    ClkMux I__3990 (
            .O(N__25042),
            .I(N__25037));
    GlobalMux I__3989 (
            .O(N__25037),
            .I(N__25034));
    gio2CtrlBuf I__3988 (
            .O(N__25034),
            .I(delay_hc_input_c_g));
    CascadeMux I__3987 (
            .O(N__25031),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__3986 (
            .O(N__25028),
            .I(N__25025));
    LocalMux I__3985 (
            .O(N__25025),
            .I(N__25022));
    Span4Mux_v I__3984 (
            .O(N__25022),
            .I(N__25019));
    Odrv4 I__3983 (
            .O(N__25019),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__3982 (
            .O(N__25016),
            .I(N__25013));
    InMux I__3981 (
            .O(N__25013),
            .I(N__25010));
    LocalMux I__3980 (
            .O(N__25010),
            .I(N__25007));
    Span4Mux_v I__3979 (
            .O(N__25007),
            .I(N__25004));
    Odrv4 I__3978 (
            .O(N__25004),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0 ));
    CascadeMux I__3977 (
            .O(N__25001),
            .I(\phase_controller_inst1.stoper_hc.N_45_cascade_ ));
    InMux I__3976 (
            .O(N__24998),
            .I(N__24991));
    InMux I__3975 (
            .O(N__24997),
            .I(N__24982));
    InMux I__3974 (
            .O(N__24996),
            .I(N__24982));
    InMux I__3973 (
            .O(N__24995),
            .I(N__24982));
    InMux I__3972 (
            .O(N__24994),
            .I(N__24982));
    LocalMux I__3971 (
            .O(N__24991),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__3970 (
            .O(N__24982),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__3969 (
            .O(N__24977),
            .I(N__24972));
    CascadeMux I__3968 (
            .O(N__24976),
            .I(N__24966));
    CascadeMux I__3967 (
            .O(N__24975),
            .I(N__24963));
    InMux I__3966 (
            .O(N__24972),
            .I(N__24954));
    InMux I__3965 (
            .O(N__24971),
            .I(N__24954));
    InMux I__3964 (
            .O(N__24970),
            .I(N__24954));
    InMux I__3963 (
            .O(N__24969),
            .I(N__24954));
    InMux I__3962 (
            .O(N__24966),
            .I(N__24951));
    InMux I__3961 (
            .O(N__24963),
            .I(N__24948));
    LocalMux I__3960 (
            .O(N__24954),
            .I(N__24945));
    LocalMux I__3959 (
            .O(N__24951),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__3958 (
            .O(N__24948),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__3957 (
            .O(N__24945),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    CascadeMux I__3956 (
            .O(N__24938),
            .I(N__24934));
    InMux I__3955 (
            .O(N__24937),
            .I(N__24931));
    InMux I__3954 (
            .O(N__24934),
            .I(N__24928));
    LocalMux I__3953 (
            .O(N__24931),
            .I(N__24922));
    LocalMux I__3952 (
            .O(N__24928),
            .I(N__24922));
    InMux I__3951 (
            .O(N__24927),
            .I(N__24919));
    Span4Mux_v I__3950 (
            .O(N__24922),
            .I(N__24914));
    LocalMux I__3949 (
            .O(N__24919),
            .I(N__24914));
    Span4Mux_h I__3948 (
            .O(N__24914),
            .I(N__24911));
    Odrv4 I__3947 (
            .O(N__24911),
            .I(il_max_comp2_D2));
    CascadeMux I__3946 (
            .O(N__24908),
            .I(\phase_controller_inst1.stoper_hc.N_325_cascade_ ));
    InMux I__3945 (
            .O(N__24905),
            .I(N__24902));
    LocalMux I__3944 (
            .O(N__24902),
            .I(N__24899));
    Span4Mux_h I__3943 (
            .O(N__24899),
            .I(N__24896));
    Odrv4 I__3942 (
            .O(N__24896),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2 ));
    CascadeMux I__3941 (
            .O(N__24893),
            .I(N__24888));
    InMux I__3940 (
            .O(N__24892),
            .I(N__24884));
    InMux I__3939 (
            .O(N__24891),
            .I(N__24878));
    InMux I__3938 (
            .O(N__24888),
            .I(N__24875));
    InMux I__3937 (
            .O(N__24887),
            .I(N__24872));
    LocalMux I__3936 (
            .O(N__24884),
            .I(N__24869));
    InMux I__3935 (
            .O(N__24883),
            .I(N__24865));
    InMux I__3934 (
            .O(N__24882),
            .I(N__24861));
    InMux I__3933 (
            .O(N__24881),
            .I(N__24858));
    LocalMux I__3932 (
            .O(N__24878),
            .I(N__24855));
    LocalMux I__3931 (
            .O(N__24875),
            .I(N__24850));
    LocalMux I__3930 (
            .O(N__24872),
            .I(N__24850));
    Span4Mux_v I__3929 (
            .O(N__24869),
            .I(N__24847));
    InMux I__3928 (
            .O(N__24868),
            .I(N__24844));
    LocalMux I__3927 (
            .O(N__24865),
            .I(N__24841));
    InMux I__3926 (
            .O(N__24864),
            .I(N__24838));
    LocalMux I__3925 (
            .O(N__24861),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    LocalMux I__3924 (
            .O(N__24858),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    Odrv4 I__3923 (
            .O(N__24855),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    Odrv4 I__3922 (
            .O(N__24850),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    Odrv4 I__3921 (
            .O(N__24847),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    LocalMux I__3920 (
            .O(N__24844),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    Odrv4 I__3919 (
            .O(N__24841),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    LocalMux I__3918 (
            .O(N__24838),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    CascadeMux I__3917 (
            .O(N__24821),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2_cascade_ ));
    CascadeMux I__3916 (
            .O(N__24818),
            .I(\phase_controller_inst1.stoper_hc.N_307_cascade_ ));
    CascadeMux I__3915 (
            .O(N__24815),
            .I(N__24812));
    InMux I__3914 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__3913 (
            .O(N__24809),
            .I(N__24806));
    Span4Mux_h I__3912 (
            .O(N__24806),
            .I(N__24801));
    InMux I__3911 (
            .O(N__24805),
            .I(N__24796));
    InMux I__3910 (
            .O(N__24804),
            .I(N__24796));
    Odrv4 I__3909 (
            .O(N__24801),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__3908 (
            .O(N__24796),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    CascadeMux I__3907 (
            .O(N__24791),
            .I(N__24788));
    InMux I__3906 (
            .O(N__24788),
            .I(N__24783));
    InMux I__3905 (
            .O(N__24787),
            .I(N__24778));
    InMux I__3904 (
            .O(N__24786),
            .I(N__24778));
    LocalMux I__3903 (
            .O(N__24783),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2 ));
    LocalMux I__3902 (
            .O(N__24778),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2 ));
    CascadeMux I__3901 (
            .O(N__24773),
            .I(N__24768));
    CascadeMux I__3900 (
            .O(N__24772),
            .I(N__24765));
    InMux I__3899 (
            .O(N__24771),
            .I(N__24762));
    InMux I__3898 (
            .O(N__24768),
            .I(N__24757));
    InMux I__3897 (
            .O(N__24765),
            .I(N__24757));
    LocalMux I__3896 (
            .O(N__24762),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_1Z0Z_2 ));
    LocalMux I__3895 (
            .O(N__24757),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_1Z0Z_2 ));
    CascadeMux I__3894 (
            .O(N__24752),
            .I(N__24745));
    InMux I__3893 (
            .O(N__24751),
            .I(N__24728));
    InMux I__3892 (
            .O(N__24750),
            .I(N__24728));
    InMux I__3891 (
            .O(N__24749),
            .I(N__24728));
    InMux I__3890 (
            .O(N__24748),
            .I(N__24728));
    InMux I__3889 (
            .O(N__24745),
            .I(N__24715));
    InMux I__3888 (
            .O(N__24744),
            .I(N__24715));
    InMux I__3887 (
            .O(N__24743),
            .I(N__24715));
    InMux I__3886 (
            .O(N__24742),
            .I(N__24715));
    InMux I__3885 (
            .O(N__24741),
            .I(N__24715));
    InMux I__3884 (
            .O(N__24740),
            .I(N__24710));
    InMux I__3883 (
            .O(N__24739),
            .I(N__24710));
    InMux I__3882 (
            .O(N__24738),
            .I(N__24705));
    InMux I__3881 (
            .O(N__24737),
            .I(N__24705));
    LocalMux I__3880 (
            .O(N__24728),
            .I(N__24702));
    CascadeMux I__3879 (
            .O(N__24727),
            .I(N__24696));
    CascadeMux I__3878 (
            .O(N__24726),
            .I(N__24693));
    LocalMux I__3877 (
            .O(N__24715),
            .I(N__24681));
    LocalMux I__3876 (
            .O(N__24710),
            .I(N__24681));
    LocalMux I__3875 (
            .O(N__24705),
            .I(N__24681));
    Span4Mux_v I__3874 (
            .O(N__24702),
            .I(N__24678));
    InMux I__3873 (
            .O(N__24701),
            .I(N__24675));
    CascadeMux I__3872 (
            .O(N__24700),
            .I(N__24671));
    InMux I__3871 (
            .O(N__24699),
            .I(N__24651));
    InMux I__3870 (
            .O(N__24696),
            .I(N__24651));
    InMux I__3869 (
            .O(N__24693),
            .I(N__24651));
    InMux I__3868 (
            .O(N__24692),
            .I(N__24651));
    InMux I__3867 (
            .O(N__24691),
            .I(N__24651));
    InMux I__3866 (
            .O(N__24690),
            .I(N__24651));
    InMux I__3865 (
            .O(N__24689),
            .I(N__24651));
    InMux I__3864 (
            .O(N__24688),
            .I(N__24651));
    Span4Mux_v I__3863 (
            .O(N__24681),
            .I(N__24646));
    Span4Mux_h I__3862 (
            .O(N__24678),
            .I(N__24646));
    LocalMux I__3861 (
            .O(N__24675),
            .I(N__24643));
    InMux I__3860 (
            .O(N__24674),
            .I(N__24638));
    InMux I__3859 (
            .O(N__24671),
            .I(N__24638));
    InMux I__3858 (
            .O(N__24670),
            .I(N__24631));
    InMux I__3857 (
            .O(N__24669),
            .I(N__24631));
    InMux I__3856 (
            .O(N__24668),
            .I(N__24631));
    LocalMux I__3855 (
            .O(N__24651),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15 ));
    Odrv4 I__3854 (
            .O(N__24646),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15 ));
    Odrv4 I__3853 (
            .O(N__24643),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15 ));
    LocalMux I__3852 (
            .O(N__24638),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15 ));
    LocalMux I__3851 (
            .O(N__24631),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15 ));
    InMux I__3850 (
            .O(N__24620),
            .I(N__24617));
    LocalMux I__3849 (
            .O(N__24617),
            .I(N__24614));
    Span4Mux_v I__3848 (
            .O(N__24614),
            .I(N__24611));
    Span4Mux_h I__3847 (
            .O(N__24611),
            .I(N__24608));
    Odrv4 I__3846 (
            .O(N__24608),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__3845 (
            .O(N__24605),
            .I(N__24601));
    InMux I__3844 (
            .O(N__24604),
            .I(N__24598));
    LocalMux I__3843 (
            .O(N__24601),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__3842 (
            .O(N__24598),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__3841 (
            .O(N__24593),
            .I(N__24590));
    InMux I__3840 (
            .O(N__24590),
            .I(N__24587));
    LocalMux I__3839 (
            .O(N__24587),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__3838 (
            .O(N__24584),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__3837 (
            .O(N__24581),
            .I(N__24578));
    LocalMux I__3836 (
            .O(N__24578),
            .I(N__24575));
    Odrv4 I__3835 (
            .O(N__24575),
            .I(il_max_comp1_D1));
    InMux I__3834 (
            .O(N__24572),
            .I(N__24568));
    InMux I__3833 (
            .O(N__24571),
            .I(N__24565));
    LocalMux I__3832 (
            .O(N__24568),
            .I(N__24561));
    LocalMux I__3831 (
            .O(N__24565),
            .I(N__24558));
    InMux I__3830 (
            .O(N__24564),
            .I(N__24555));
    Span12Mux_h I__3829 (
            .O(N__24561),
            .I(N__24552));
    Span4Mux_h I__3828 (
            .O(N__24558),
            .I(N__24547));
    LocalMux I__3827 (
            .O(N__24555),
            .I(N__24547));
    Odrv12 I__3826 (
            .O(N__24552),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    Odrv4 I__3825 (
            .O(N__24547),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__3824 (
            .O(N__24542),
            .I(N__24539));
    LocalMux I__3823 (
            .O(N__24539),
            .I(N__24536));
    Span4Mux_v I__3822 (
            .O(N__24536),
            .I(N__24533));
    Odrv4 I__3821 (
            .O(N__24533),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ));
    InMux I__3820 (
            .O(N__24530),
            .I(N__24527));
    LocalMux I__3819 (
            .O(N__24527),
            .I(N__24519));
    InMux I__3818 (
            .O(N__24526),
            .I(N__24516));
    InMux I__3817 (
            .O(N__24525),
            .I(N__24511));
    InMux I__3816 (
            .O(N__24524),
            .I(N__24511));
    InMux I__3815 (
            .O(N__24523),
            .I(N__24506));
    InMux I__3814 (
            .O(N__24522),
            .I(N__24506));
    Span4Mux_h I__3813 (
            .O(N__24519),
            .I(N__24503));
    LocalMux I__3812 (
            .O(N__24516),
            .I(N__24500));
    LocalMux I__3811 (
            .O(N__24511),
            .I(N__24495));
    LocalMux I__3810 (
            .O(N__24506),
            .I(N__24495));
    Span4Mux_v I__3809 (
            .O(N__24503),
            .I(N__24492));
    Span4Mux_v I__3808 (
            .O(N__24500),
            .I(N__24487));
    Span4Mux_v I__3807 (
            .O(N__24495),
            .I(N__24487));
    Odrv4 I__3806 (
            .O(N__24492),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__3805 (
            .O(N__24487),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__3804 (
            .O(N__24482),
            .I(N__24475));
    InMux I__3803 (
            .O(N__24481),
            .I(N__24475));
    InMux I__3802 (
            .O(N__24480),
            .I(N__24471));
    LocalMux I__3801 (
            .O(N__24475),
            .I(N__24468));
    InMux I__3800 (
            .O(N__24474),
            .I(N__24465));
    LocalMux I__3799 (
            .O(N__24471),
            .I(N__24461));
    Span4Mux_h I__3798 (
            .O(N__24468),
            .I(N__24458));
    LocalMux I__3797 (
            .O(N__24465),
            .I(N__24455));
    InMux I__3796 (
            .O(N__24464),
            .I(N__24452));
    Odrv12 I__3795 (
            .O(N__24461),
            .I(elapsed_time_ns_1_RNI62CED1_0_19));
    Odrv4 I__3794 (
            .O(N__24458),
            .I(elapsed_time_ns_1_RNI62CED1_0_19));
    Odrv4 I__3793 (
            .O(N__24455),
            .I(elapsed_time_ns_1_RNI62CED1_0_19));
    LocalMux I__3792 (
            .O(N__24452),
            .I(elapsed_time_ns_1_RNI62CED1_0_19));
    CascadeMux I__3791 (
            .O(N__24443),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_));
    InMux I__3790 (
            .O(N__24440),
            .I(N__24435));
    CascadeMux I__3789 (
            .O(N__24439),
            .I(N__24432));
    InMux I__3788 (
            .O(N__24438),
            .I(N__24429));
    LocalMux I__3787 (
            .O(N__24435),
            .I(N__24426));
    InMux I__3786 (
            .O(N__24432),
            .I(N__24423));
    LocalMux I__3785 (
            .O(N__24429),
            .I(N__24418));
    Span4Mux_h I__3784 (
            .O(N__24426),
            .I(N__24418));
    LocalMux I__3783 (
            .O(N__24423),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_a5_1_1_9 ));
    Odrv4 I__3782 (
            .O(N__24418),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_a5_1_1_9 ));
    InMux I__3781 (
            .O(N__24413),
            .I(N__24410));
    LocalMux I__3780 (
            .O(N__24410),
            .I(N__24405));
    InMux I__3779 (
            .O(N__24409),
            .I(N__24401));
    InMux I__3778 (
            .O(N__24408),
            .I(N__24398));
    Span4Mux_h I__3777 (
            .O(N__24405),
            .I(N__24395));
    InMux I__3776 (
            .O(N__24404),
            .I(N__24392));
    LocalMux I__3775 (
            .O(N__24401),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9 ));
    LocalMux I__3774 (
            .O(N__24398),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9 ));
    Odrv4 I__3773 (
            .O(N__24395),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9 ));
    LocalMux I__3772 (
            .O(N__24392),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9 ));
    InMux I__3771 (
            .O(N__24383),
            .I(N__24380));
    LocalMux I__3770 (
            .O(N__24380),
            .I(N__24377));
    Odrv12 I__3769 (
            .O(N__24377),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1Z0Z_6 ));
    InMux I__3768 (
            .O(N__24374),
            .I(N__24370));
    InMux I__3767 (
            .O(N__24373),
            .I(N__24367));
    LocalMux I__3766 (
            .O(N__24370),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__3765 (
            .O(N__24367),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__3764 (
            .O(N__24362),
            .I(N__24359));
    LocalMux I__3763 (
            .O(N__24359),
            .I(N__24356));
    Span4Mux_v I__3762 (
            .O(N__24356),
            .I(N__24353));
    Odrv4 I__3761 (
            .O(N__24353),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__3760 (
            .O(N__24350),
            .I(N__24347));
    InMux I__3759 (
            .O(N__24347),
            .I(N__24344));
    LocalMux I__3758 (
            .O(N__24344),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__3757 (
            .O(N__24341),
            .I(N__24338));
    LocalMux I__3756 (
            .O(N__24338),
            .I(N__24335));
    Span4Mux_v I__3755 (
            .O(N__24335),
            .I(N__24332));
    Sp12to4 I__3754 (
            .O(N__24332),
            .I(N__24329));
    Odrv12 I__3753 (
            .O(N__24329),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__3752 (
            .O(N__24326),
            .I(N__24322));
    InMux I__3751 (
            .O(N__24325),
            .I(N__24319));
    LocalMux I__3750 (
            .O(N__24322),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__3749 (
            .O(N__24319),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__3748 (
            .O(N__24314),
            .I(N__24311));
    InMux I__3747 (
            .O(N__24311),
            .I(N__24308));
    LocalMux I__3746 (
            .O(N__24308),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__3745 (
            .O(N__24305),
            .I(N__24301));
    InMux I__3744 (
            .O(N__24304),
            .I(N__24298));
    LocalMux I__3743 (
            .O(N__24301),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__3742 (
            .O(N__24298),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__3741 (
            .O(N__24293),
            .I(N__24290));
    InMux I__3740 (
            .O(N__24290),
            .I(N__24287));
    LocalMux I__3739 (
            .O(N__24287),
            .I(N__24284));
    Odrv12 I__3738 (
            .O(N__24284),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__3737 (
            .O(N__24281),
            .I(N__24278));
    LocalMux I__3736 (
            .O(N__24278),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__3735 (
            .O(N__24275),
            .I(N__24272));
    LocalMux I__3734 (
            .O(N__24272),
            .I(N__24269));
    Span4Mux_h I__3733 (
            .O(N__24269),
            .I(N__24266));
    Odrv4 I__3732 (
            .O(N__24266),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__3731 (
            .O(N__24263),
            .I(N__24259));
    InMux I__3730 (
            .O(N__24262),
            .I(N__24256));
    LocalMux I__3729 (
            .O(N__24259),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__3728 (
            .O(N__24256),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__3727 (
            .O(N__24251),
            .I(N__24248));
    InMux I__3726 (
            .O(N__24248),
            .I(N__24245));
    LocalMux I__3725 (
            .O(N__24245),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__3724 (
            .O(N__24242),
            .I(N__24239));
    LocalMux I__3723 (
            .O(N__24239),
            .I(N__24236));
    Span4Mux_h I__3722 (
            .O(N__24236),
            .I(N__24233));
    Odrv4 I__3721 (
            .O(N__24233),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__3720 (
            .O(N__24230),
            .I(N__24226));
    InMux I__3719 (
            .O(N__24229),
            .I(N__24223));
    LocalMux I__3718 (
            .O(N__24226),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__3717 (
            .O(N__24223),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__3716 (
            .O(N__24218),
            .I(N__24215));
    InMux I__3715 (
            .O(N__24215),
            .I(N__24212));
    LocalMux I__3714 (
            .O(N__24212),
            .I(N__24209));
    Odrv4 I__3713 (
            .O(N__24209),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    InMux I__3712 (
            .O(N__24206),
            .I(N__24203));
    LocalMux I__3711 (
            .O(N__24203),
            .I(N__24200));
    Span4Mux_h I__3710 (
            .O(N__24200),
            .I(N__24197));
    Span4Mux_h I__3709 (
            .O(N__24197),
            .I(N__24194));
    Odrv4 I__3708 (
            .O(N__24194),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__3707 (
            .O(N__24191),
            .I(N__24187));
    InMux I__3706 (
            .O(N__24190),
            .I(N__24184));
    LocalMux I__3705 (
            .O(N__24187),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__3704 (
            .O(N__24184),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__3703 (
            .O(N__24179),
            .I(N__24176));
    InMux I__3702 (
            .O(N__24176),
            .I(N__24173));
    LocalMux I__3701 (
            .O(N__24173),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    InMux I__3700 (
            .O(N__24170),
            .I(N__24167));
    LocalMux I__3699 (
            .O(N__24167),
            .I(N__24164));
    Span4Mux_h I__3698 (
            .O(N__24164),
            .I(N__24161));
    Span4Mux_h I__3697 (
            .O(N__24161),
            .I(N__24158));
    Odrv4 I__3696 (
            .O(N__24158),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    InMux I__3695 (
            .O(N__24155),
            .I(N__24151));
    InMux I__3694 (
            .O(N__24154),
            .I(N__24148));
    LocalMux I__3693 (
            .O(N__24151),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__3692 (
            .O(N__24148),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__3691 (
            .O(N__24143),
            .I(N__24140));
    InMux I__3690 (
            .O(N__24140),
            .I(N__24137));
    LocalMux I__3689 (
            .O(N__24137),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    InMux I__3688 (
            .O(N__24134),
            .I(N__24130));
    InMux I__3687 (
            .O(N__24133),
            .I(N__24127));
    LocalMux I__3686 (
            .O(N__24130),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__3685 (
            .O(N__24127),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__3684 (
            .O(N__24122),
            .I(N__24119));
    InMux I__3683 (
            .O(N__24119),
            .I(N__24116));
    LocalMux I__3682 (
            .O(N__24116),
            .I(N__24113));
    Odrv4 I__3681 (
            .O(N__24113),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__3680 (
            .O(N__24110),
            .I(N__24106));
    InMux I__3679 (
            .O(N__24109),
            .I(N__24103));
    LocalMux I__3678 (
            .O(N__24106),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__3677 (
            .O(N__24103),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__3676 (
            .O(N__24098),
            .I(N__24095));
    InMux I__3675 (
            .O(N__24095),
            .I(N__24092));
    LocalMux I__3674 (
            .O(N__24092),
            .I(N__24089));
    Odrv4 I__3673 (
            .O(N__24089),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__3672 (
            .O(N__24086),
            .I(N__24082));
    InMux I__3671 (
            .O(N__24085),
            .I(N__24079));
    LocalMux I__3670 (
            .O(N__24082),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__3669 (
            .O(N__24079),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__3668 (
            .O(N__24074),
            .I(N__24071));
    InMux I__3667 (
            .O(N__24071),
            .I(N__24068));
    LocalMux I__3666 (
            .O(N__24068),
            .I(N__24065));
    Odrv4 I__3665 (
            .O(N__24065),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__3664 (
            .O(N__24062),
            .I(N__24059));
    LocalMux I__3663 (
            .O(N__24059),
            .I(N__24056));
    Span4Mux_h I__3662 (
            .O(N__24056),
            .I(N__24053));
    Odrv4 I__3661 (
            .O(N__24053),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__3660 (
            .O(N__24050),
            .I(N__24046));
    InMux I__3659 (
            .O(N__24049),
            .I(N__24043));
    LocalMux I__3658 (
            .O(N__24046),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__3657 (
            .O(N__24043),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__3656 (
            .O(N__24038),
            .I(N__24035));
    InMux I__3655 (
            .O(N__24035),
            .I(N__24032));
    LocalMux I__3654 (
            .O(N__24032),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__3653 (
            .O(N__24029),
            .I(N__24025));
    InMux I__3652 (
            .O(N__24028),
            .I(N__24022));
    LocalMux I__3651 (
            .O(N__24025),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__3650 (
            .O(N__24022),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__3649 (
            .O(N__24017),
            .I(N__24014));
    InMux I__3648 (
            .O(N__24014),
            .I(N__24011));
    LocalMux I__3647 (
            .O(N__24011),
            .I(N__24008));
    Odrv4 I__3646 (
            .O(N__24008),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__3645 (
            .O(N__24005),
            .I(N__24002));
    LocalMux I__3644 (
            .O(N__24002),
            .I(N__23999));
    Span4Mux_v I__3643 (
            .O(N__23999),
            .I(N__23996));
    Odrv4 I__3642 (
            .O(N__23996),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__3641 (
            .O(N__23993),
            .I(N__23989));
    InMux I__3640 (
            .O(N__23992),
            .I(N__23986));
    LocalMux I__3639 (
            .O(N__23989),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__3638 (
            .O(N__23986),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__3637 (
            .O(N__23981),
            .I(N__23978));
    InMux I__3636 (
            .O(N__23978),
            .I(N__23975));
    LocalMux I__3635 (
            .O(N__23975),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__3634 (
            .O(N__23972),
            .I(N__23969));
    LocalMux I__3633 (
            .O(N__23969),
            .I(N__23966));
    Span4Mux_h I__3632 (
            .O(N__23966),
            .I(N__23963));
    Odrv4 I__3631 (
            .O(N__23963),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__3630 (
            .O(N__23960),
            .I(N__23956));
    InMux I__3629 (
            .O(N__23959),
            .I(N__23953));
    LocalMux I__3628 (
            .O(N__23956),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__3627 (
            .O(N__23953),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__3626 (
            .O(N__23948),
            .I(N__23945));
    InMux I__3625 (
            .O(N__23945),
            .I(N__23942));
    LocalMux I__3624 (
            .O(N__23942),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__3623 (
            .O(N__23939),
            .I(N__23935));
    InMux I__3622 (
            .O(N__23938),
            .I(N__23932));
    LocalMux I__3621 (
            .O(N__23935),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__3620 (
            .O(N__23932),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__3619 (
            .O(N__23927),
            .I(N__23924));
    LocalMux I__3618 (
            .O(N__23924),
            .I(N__23921));
    Span4Mux_v I__3617 (
            .O(N__23921),
            .I(N__23918));
    Odrv4 I__3616 (
            .O(N__23918),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__3615 (
            .O(N__23915),
            .I(N__23912));
    InMux I__3614 (
            .O(N__23912),
            .I(N__23909));
    LocalMux I__3613 (
            .O(N__23909),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    IoInMux I__3612 (
            .O(N__23906),
            .I(N__23903));
    LocalMux I__3611 (
            .O(N__23903),
            .I(N__23900));
    Odrv4 I__3610 (
            .O(N__23900),
            .I(s3_phy_c));
    InMux I__3609 (
            .O(N__23897),
            .I(N__23894));
    LocalMux I__3608 (
            .O(N__23894),
            .I(N__23891));
    Span4Mux_h I__3607 (
            .O(N__23891),
            .I(N__23888));
    Span4Mux_v I__3606 (
            .O(N__23888),
            .I(N__23885));
    Odrv4 I__3605 (
            .O(N__23885),
            .I(il_min_comp1_c));
    InMux I__3604 (
            .O(N__23882),
            .I(N__23879));
    LocalMux I__3603 (
            .O(N__23879),
            .I(N__23876));
    Odrv4 I__3602 (
            .O(N__23876),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__3601 (
            .O(N__23873),
            .I(N__23870));
    LocalMux I__3600 (
            .O(N__23870),
            .I(N__23867));
    Odrv4 I__3599 (
            .O(N__23867),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__3598 (
            .O(N__23864),
            .I(N__23861));
    LocalMux I__3597 (
            .O(N__23861),
            .I(N__23858));
    Odrv12 I__3596 (
            .O(N__23858),
            .I(il_min_comp1_D1));
    InMux I__3595 (
            .O(N__23855),
            .I(N__23852));
    LocalMux I__3594 (
            .O(N__23852),
            .I(N__23849));
    Span4Mux_h I__3593 (
            .O(N__23849),
            .I(N__23846));
    Span4Mux_v I__3592 (
            .O(N__23846),
            .I(N__23843));
    Span4Mux_v I__3591 (
            .O(N__23843),
            .I(N__23840));
    Odrv4 I__3590 (
            .O(N__23840),
            .I(il_max_comp1_c));
    CascadeMux I__3589 (
            .O(N__23837),
            .I(N__23834));
    InMux I__3588 (
            .O(N__23834),
            .I(N__23831));
    LocalMux I__3587 (
            .O(N__23831),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__3586 (
            .O(N__23828),
            .I(N__23824));
    InMux I__3585 (
            .O(N__23827),
            .I(N__23821));
    LocalMux I__3584 (
            .O(N__23824),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__3583 (
            .O(N__23821),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__3582 (
            .O(N__23816),
            .I(N__23813));
    InMux I__3581 (
            .O(N__23813),
            .I(N__23810));
    LocalMux I__3580 (
            .O(N__23810),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__3579 (
            .O(N__23807),
            .I(N__23803));
    InMux I__3578 (
            .O(N__23806),
            .I(N__23800));
    LocalMux I__3577 (
            .O(N__23803),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__3576 (
            .O(N__23800),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__3575 (
            .O(N__23795),
            .I(N__23792));
    InMux I__3574 (
            .O(N__23792),
            .I(N__23789));
    LocalMux I__3573 (
            .O(N__23789),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__3572 (
            .O(N__23786),
            .I(N__23782));
    InMux I__3571 (
            .O(N__23785),
            .I(N__23779));
    LocalMux I__3570 (
            .O(N__23782),
            .I(N__23776));
    LocalMux I__3569 (
            .O(N__23779),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4 ));
    Odrv4 I__3568 (
            .O(N__23776),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4 ));
    InMux I__3567 (
            .O(N__23771),
            .I(N__23768));
    LocalMux I__3566 (
            .O(N__23768),
            .I(N__23763));
    InMux I__3565 (
            .O(N__23767),
            .I(N__23758));
    InMux I__3564 (
            .O(N__23766),
            .I(N__23758));
    Odrv4 I__3563 (
            .O(N__23763),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ));
    LocalMux I__3562 (
            .O(N__23758),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ));
    InMux I__3561 (
            .O(N__23753),
            .I(N__23749));
    InMux I__3560 (
            .O(N__23752),
            .I(N__23746));
    LocalMux I__3559 (
            .O(N__23749),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ));
    LocalMux I__3558 (
            .O(N__23746),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ));
    InMux I__3557 (
            .O(N__23741),
            .I(N__23736));
    InMux I__3556 (
            .O(N__23740),
            .I(N__23731));
    InMux I__3555 (
            .O(N__23739),
            .I(N__23731));
    LocalMux I__3554 (
            .O(N__23736),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ));
    LocalMux I__3553 (
            .O(N__23731),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ));
    CascadeMux I__3552 (
            .O(N__23726),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_ ));
    CascadeMux I__3551 (
            .O(N__23723),
            .I(N__23719));
    InMux I__3550 (
            .O(N__23722),
            .I(N__23716));
    InMux I__3549 (
            .O(N__23719),
            .I(N__23713));
    LocalMux I__3548 (
            .O(N__23716),
            .I(N__23707));
    LocalMux I__3547 (
            .O(N__23713),
            .I(N__23707));
    InMux I__3546 (
            .O(N__23712),
            .I(N__23704));
    Odrv4 I__3545 (
            .O(N__23707),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    LocalMux I__3544 (
            .O(N__23704),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    CascadeMux I__3543 (
            .O(N__23699),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_ ));
    CascadeMux I__3542 (
            .O(N__23696),
            .I(N__23692));
    InMux I__3541 (
            .O(N__23695),
            .I(N__23688));
    InMux I__3540 (
            .O(N__23692),
            .I(N__23685));
    InMux I__3539 (
            .O(N__23691),
            .I(N__23682));
    LocalMux I__3538 (
            .O(N__23688),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__3537 (
            .O(N__23685),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__3536 (
            .O(N__23682),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    CascadeMux I__3535 (
            .O(N__23675),
            .I(N__23671));
    InMux I__3534 (
            .O(N__23674),
            .I(N__23667));
    InMux I__3533 (
            .O(N__23671),
            .I(N__23664));
    InMux I__3532 (
            .O(N__23670),
            .I(N__23661));
    LocalMux I__3531 (
            .O(N__23667),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__3530 (
            .O(N__23664),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__3529 (
            .O(N__23661),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    CEMux I__3528 (
            .O(N__23654),
            .I(N__23639));
    CEMux I__3527 (
            .O(N__23653),
            .I(N__23639));
    CEMux I__3526 (
            .O(N__23652),
            .I(N__23639));
    CEMux I__3525 (
            .O(N__23651),
            .I(N__23639));
    CEMux I__3524 (
            .O(N__23650),
            .I(N__23639));
    GlobalMux I__3523 (
            .O(N__23639),
            .I(N__23636));
    gio2CtrlBuf I__3522 (
            .O(N__23636),
            .I(\delay_measurement_inst.delay_hc_timer.N_432_i_g ));
    IoInMux I__3521 (
            .O(N__23633),
            .I(N__23630));
    LocalMux I__3520 (
            .O(N__23630),
            .I(N__23627));
    Span4Mux_s0_v I__3519 (
            .O(N__23627),
            .I(N__23624));
    Span4Mux_h I__3518 (
            .O(N__23624),
            .I(N__23621));
    Span4Mux_v I__3517 (
            .O(N__23621),
            .I(N__23618));
    Span4Mux_v I__3516 (
            .O(N__23618),
            .I(N__23615));
    Odrv4 I__3515 (
            .O(N__23615),
            .I(\delay_measurement_inst.delay_hc_timer.N_432_i ));
    InMux I__3514 (
            .O(N__23612),
            .I(N__23609));
    LocalMux I__3513 (
            .O(N__23609),
            .I(N__23606));
    Span4Mux_v I__3512 (
            .O(N__23606),
            .I(N__23603));
    Span4Mux_v I__3511 (
            .O(N__23603),
            .I(N__23600));
    Span4Mux_v I__3510 (
            .O(N__23600),
            .I(N__23597));
    Odrv4 I__3509 (
            .O(N__23597),
            .I(il_min_comp2_D1));
    InMux I__3508 (
            .O(N__23594),
            .I(N__23591));
    LocalMux I__3507 (
            .O(N__23591),
            .I(N__23587));
    InMux I__3506 (
            .O(N__23590),
            .I(N__23584));
    Span4Mux_h I__3505 (
            .O(N__23587),
            .I(N__23581));
    LocalMux I__3504 (
            .O(N__23584),
            .I(N__23578));
    Odrv4 I__3503 (
            .O(N__23581),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv12 I__3502 (
            .O(N__23578),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    CascadeMux I__3501 (
            .O(N__23573),
            .I(N__23570));
    InMux I__3500 (
            .O(N__23570),
            .I(N__23567));
    LocalMux I__3499 (
            .O(N__23567),
            .I(elapsed_time_ns_1_RNIT6ND11_0_25));
    CascadeMux I__3498 (
            .O(N__23564),
            .I(elapsed_time_ns_1_RNIT6ND11_0_25_cascade_));
    InMux I__3497 (
            .O(N__23561),
            .I(N__23558));
    LocalMux I__3496 (
            .O(N__23558),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_o5_6Z0Z_15 ));
    InMux I__3495 (
            .O(N__23555),
            .I(N__23551));
    InMux I__3494 (
            .O(N__23554),
            .I(N__23548));
    LocalMux I__3493 (
            .O(N__23551),
            .I(N__23543));
    LocalMux I__3492 (
            .O(N__23548),
            .I(N__23543));
    Span4Mux_h I__3491 (
            .O(N__23543),
            .I(N__23540));
    Odrv4 I__3490 (
            .O(N__23540),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__3489 (
            .O(N__23537),
            .I(N__23531));
    InMux I__3488 (
            .O(N__23536),
            .I(N__23531));
    LocalMux I__3487 (
            .O(N__23531),
            .I(elapsed_time_ns_1_RNIV8ND11_0_27));
    InMux I__3486 (
            .O(N__23528),
            .I(N__23524));
    InMux I__3485 (
            .O(N__23527),
            .I(N__23521));
    LocalMux I__3484 (
            .O(N__23524),
            .I(N__23516));
    LocalMux I__3483 (
            .O(N__23521),
            .I(N__23516));
    Span4Mux_h I__3482 (
            .O(N__23516),
            .I(N__23513));
    Odrv4 I__3481 (
            .O(N__23513),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__3480 (
            .O(N__23510),
            .I(N__23504));
    InMux I__3479 (
            .O(N__23509),
            .I(N__23504));
    LocalMux I__3478 (
            .O(N__23504),
            .I(elapsed_time_ns_1_RNIU7ND11_0_26));
    InMux I__3477 (
            .O(N__23501),
            .I(N__23498));
    LocalMux I__3476 (
            .O(N__23498),
            .I(N__23494));
    InMux I__3475 (
            .O(N__23497),
            .I(N__23491));
    Span4Mux_h I__3474 (
            .O(N__23494),
            .I(N__23488));
    LocalMux I__3473 (
            .O(N__23491),
            .I(N__23485));
    Odrv4 I__3472 (
            .O(N__23488),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    Odrv12 I__3471 (
            .O(N__23485),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    CascadeMux I__3470 (
            .O(N__23480),
            .I(N__23477));
    InMux I__3469 (
            .O(N__23477),
            .I(N__23473));
    InMux I__3468 (
            .O(N__23476),
            .I(N__23470));
    LocalMux I__3467 (
            .O(N__23473),
            .I(elapsed_time_ns_1_RNI0AND11_0_28));
    LocalMux I__3466 (
            .O(N__23470),
            .I(elapsed_time_ns_1_RNI0AND11_0_28));
    CascadeMux I__3465 (
            .O(N__23465),
            .I(N__23461));
    InMux I__3464 (
            .O(N__23464),
            .I(N__23458));
    InMux I__3463 (
            .O(N__23461),
            .I(N__23455));
    LocalMux I__3462 (
            .O(N__23458),
            .I(N__23452));
    LocalMux I__3461 (
            .O(N__23455),
            .I(N__23449));
    Span4Mux_h I__3460 (
            .O(N__23452),
            .I(N__23446));
    Span4Mux_h I__3459 (
            .O(N__23449),
            .I(N__23443));
    Odrv4 I__3458 (
            .O(N__23446),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__3457 (
            .O(N__23443),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__3456 (
            .O(N__23438),
            .I(N__23434));
    InMux I__3455 (
            .O(N__23437),
            .I(N__23431));
    LocalMux I__3454 (
            .O(N__23434),
            .I(N__23428));
    LocalMux I__3453 (
            .O(N__23431),
            .I(elapsed_time_ns_1_RNIP3OD11_0_30));
    Odrv4 I__3452 (
            .O(N__23428),
            .I(elapsed_time_ns_1_RNIP3OD11_0_30));
    InMux I__3451 (
            .O(N__23423),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__3450 (
            .O(N__23420),
            .I(N__23417));
    LocalMux I__3449 (
            .O(N__23417),
            .I(N__23413));
    InMux I__3448 (
            .O(N__23416),
            .I(N__23408));
    Span4Mux_v I__3447 (
            .O(N__23413),
            .I(N__23405));
    InMux I__3446 (
            .O(N__23412),
            .I(N__23402));
    InMux I__3445 (
            .O(N__23411),
            .I(N__23398));
    LocalMux I__3444 (
            .O(N__23408),
            .I(N__23391));
    Span4Mux_h I__3443 (
            .O(N__23405),
            .I(N__23391));
    LocalMux I__3442 (
            .O(N__23402),
            .I(N__23391));
    InMux I__3441 (
            .O(N__23401),
            .I(N__23388));
    LocalMux I__3440 (
            .O(N__23398),
            .I(elapsed_time_ns_1_RNI40CED1_0_17));
    Odrv4 I__3439 (
            .O(N__23391),
            .I(elapsed_time_ns_1_RNI40CED1_0_17));
    LocalMux I__3438 (
            .O(N__23388),
            .I(elapsed_time_ns_1_RNI40CED1_0_17));
    InMux I__3437 (
            .O(N__23381),
            .I(N__23378));
    LocalMux I__3436 (
            .O(N__23378),
            .I(N__23372));
    InMux I__3435 (
            .O(N__23377),
            .I(N__23369));
    InMux I__3434 (
            .O(N__23376),
            .I(N__23366));
    InMux I__3433 (
            .O(N__23375),
            .I(N__23363));
    Span4Mux_h I__3432 (
            .O(N__23372),
            .I(N__23360));
    LocalMux I__3431 (
            .O(N__23369),
            .I(N__23357));
    LocalMux I__3430 (
            .O(N__23366),
            .I(N__23354));
    LocalMux I__3429 (
            .O(N__23363),
            .I(elapsed_time_ns_1_RNI51CED1_0_18));
    Odrv4 I__3428 (
            .O(N__23360),
            .I(elapsed_time_ns_1_RNI51CED1_0_18));
    Odrv4 I__3427 (
            .O(N__23357),
            .I(elapsed_time_ns_1_RNI51CED1_0_18));
    Odrv4 I__3426 (
            .O(N__23354),
            .I(elapsed_time_ns_1_RNI51CED1_0_18));
    InMux I__3425 (
            .O(N__23345),
            .I(N__23342));
    LocalMux I__3424 (
            .O(N__23342),
            .I(N__23337));
    InMux I__3423 (
            .O(N__23341),
            .I(N__23333));
    InMux I__3422 (
            .O(N__23340),
            .I(N__23330));
    Span4Mux_v I__3421 (
            .O(N__23337),
            .I(N__23327));
    InMux I__3420 (
            .O(N__23336),
            .I(N__23324));
    LocalMux I__3419 (
            .O(N__23333),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16));
    LocalMux I__3418 (
            .O(N__23330),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16));
    Odrv4 I__3417 (
            .O(N__23327),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16));
    LocalMux I__3416 (
            .O(N__23324),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16));
    CascadeMux I__3415 (
            .O(N__23315),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3Z0Z_2_cascade_ ));
    InMux I__3414 (
            .O(N__23312),
            .I(N__23309));
    LocalMux I__3413 (
            .O(N__23309),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    InMux I__3412 (
            .O(N__23306),
            .I(N__23303));
    LocalMux I__3411 (
            .O(N__23303),
            .I(N__23300));
    Span4Mux_h I__3410 (
            .O(N__23300),
            .I(N__23296));
    InMux I__3409 (
            .O(N__23299),
            .I(N__23293));
    Span4Mux_h I__3408 (
            .O(N__23296),
            .I(N__23288));
    LocalMux I__3407 (
            .O(N__23293),
            .I(N__23288));
    Odrv4 I__3406 (
            .O(N__23288),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    CascadeMux I__3405 (
            .O(N__23285),
            .I(N__23282));
    InMux I__3404 (
            .O(N__23282),
            .I(N__23279));
    LocalMux I__3403 (
            .O(N__23279),
            .I(N__23276));
    Span4Mux_h I__3402 (
            .O(N__23276),
            .I(N__23272));
    InMux I__3401 (
            .O(N__23275),
            .I(N__23269));
    Span4Mux_v I__3400 (
            .O(N__23272),
            .I(N__23266));
    LocalMux I__3399 (
            .O(N__23269),
            .I(N__23263));
    Odrv4 I__3398 (
            .O(N__23266),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    Odrv12 I__3397 (
            .O(N__23263),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__3396 (
            .O(N__23258),
            .I(N__23255));
    LocalMux I__3395 (
            .O(N__23255),
            .I(elapsed_time_ns_1_RNI1BND11_0_29));
    InMux I__3394 (
            .O(N__23252),
            .I(N__23246));
    InMux I__3393 (
            .O(N__23251),
            .I(N__23246));
    LocalMux I__3392 (
            .O(N__23246),
            .I(elapsed_time_ns_1_RNIP2ND11_0_21));
    CascadeMux I__3391 (
            .O(N__23243),
            .I(elapsed_time_ns_1_RNI1BND11_0_29_cascade_));
    InMux I__3390 (
            .O(N__23240),
            .I(N__23237));
    LocalMux I__3389 (
            .O(N__23237),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_o5_0Z0Z_15 ));
    CascadeMux I__3388 (
            .O(N__23234),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_o5_7Z0Z_15_cascade_ ));
    InMux I__3387 (
            .O(N__23231),
            .I(N__23228));
    LocalMux I__3386 (
            .O(N__23228),
            .I(N__23225));
    Span4Mux_h I__3385 (
            .O(N__23225),
            .I(N__23221));
    InMux I__3384 (
            .O(N__23224),
            .I(N__23218));
    Span4Mux_h I__3383 (
            .O(N__23221),
            .I(N__23213));
    LocalMux I__3382 (
            .O(N__23218),
            .I(N__23213));
    Odrv4 I__3381 (
            .O(N__23213),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__3380 (
            .O(N__23210),
            .I(N__23204));
    InMux I__3379 (
            .O(N__23209),
            .I(N__23204));
    LocalMux I__3378 (
            .O(N__23204),
            .I(elapsed_time_ns_1_RNIO1ND11_0_20));
    InMux I__3377 (
            .O(N__23201),
            .I(N__23198));
    LocalMux I__3376 (
            .O(N__23198),
            .I(N__23194));
    InMux I__3375 (
            .O(N__23197),
            .I(N__23191));
    Span4Mux_h I__3374 (
            .O(N__23194),
            .I(N__23186));
    LocalMux I__3373 (
            .O(N__23191),
            .I(N__23186));
    Span4Mux_v I__3372 (
            .O(N__23186),
            .I(N__23183));
    Odrv4 I__3371 (
            .O(N__23183),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__3370 (
            .O(N__23180),
            .I(N__23174));
    InMux I__3369 (
            .O(N__23179),
            .I(N__23174));
    LocalMux I__3368 (
            .O(N__23174),
            .I(elapsed_time_ns_1_RNIQ3ND11_0_22));
    InMux I__3367 (
            .O(N__23171),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__3366 (
            .O(N__23168),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__3365 (
            .O(N__23165),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__3364 (
            .O(N__23162),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__3363 (
            .O(N__23159),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__3362 (
            .O(N__23156),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__3361 (
            .O(N__23153),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__3360 (
            .O(N__23150),
            .I(bfn_9_15_0_));
    InMux I__3359 (
            .O(N__23147),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__3358 (
            .O(N__23144),
            .I(N__23141));
    LocalMux I__3357 (
            .O(N__23141),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    InMux I__3356 (
            .O(N__23138),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__3355 (
            .O(N__23135),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__3354 (
            .O(N__23132),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__3353 (
            .O(N__23129),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__3352 (
            .O(N__23126),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__3351 (
            .O(N__23123),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__3350 (
            .O(N__23120),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__3349 (
            .O(N__23117),
            .I(bfn_9_14_0_));
    IoInMux I__3348 (
            .O(N__23114),
            .I(N__23111));
    LocalMux I__3347 (
            .O(N__23111),
            .I(s4_phy_c));
    CascadeMux I__3346 (
            .O(N__23108),
            .I(N__23105));
    InMux I__3345 (
            .O(N__23105),
            .I(N__23102));
    LocalMux I__3344 (
            .O(N__23102),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__3343 (
            .O(N__23099),
            .I(N__23096));
    InMux I__3342 (
            .O(N__23096),
            .I(N__23093));
    LocalMux I__3341 (
            .O(N__23093),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    InMux I__3340 (
            .O(N__23090),
            .I(N__23087));
    LocalMux I__3339 (
            .O(N__23087),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__3338 (
            .O(N__23084),
            .I(N__23081));
    InMux I__3337 (
            .O(N__23081),
            .I(N__23078));
    LocalMux I__3336 (
            .O(N__23078),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__3335 (
            .O(N__23075),
            .I(N__23072));
    LocalMux I__3334 (
            .O(N__23072),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__3333 (
            .O(N__23069),
            .I(N__23066));
    LocalMux I__3332 (
            .O(N__23066),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__3331 (
            .O(N__23063),
            .I(N__23060));
    LocalMux I__3330 (
            .O(N__23060),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__3329 (
            .O(N__23057),
            .I(N__23050));
    CascadeMux I__3328 (
            .O(N__23056),
            .I(N__23046));
    CascadeMux I__3327 (
            .O(N__23055),
            .I(N__23042));
    InMux I__3326 (
            .O(N__23054),
            .I(N__23018));
    InMux I__3325 (
            .O(N__23053),
            .I(N__23018));
    InMux I__3324 (
            .O(N__23050),
            .I(N__23018));
    InMux I__3323 (
            .O(N__23049),
            .I(N__23018));
    InMux I__3322 (
            .O(N__23046),
            .I(N__23018));
    InMux I__3321 (
            .O(N__23045),
            .I(N__23018));
    InMux I__3320 (
            .O(N__23042),
            .I(N__23018));
    InMux I__3319 (
            .O(N__23041),
            .I(N__23018));
    CascadeMux I__3318 (
            .O(N__23040),
            .I(N__23014));
    CascadeMux I__3317 (
            .O(N__23039),
            .I(N__23010));
    CascadeMux I__3316 (
            .O(N__23038),
            .I(N__23006));
    CascadeMux I__3315 (
            .O(N__23037),
            .I(N__23002));
    CascadeMux I__3314 (
            .O(N__23036),
            .I(N__22999));
    CascadeMux I__3313 (
            .O(N__23035),
            .I(N__22995));
    LocalMux I__3312 (
            .O(N__23018),
            .I(N__22991));
    InMux I__3311 (
            .O(N__23017),
            .I(N__22974));
    InMux I__3310 (
            .O(N__23014),
            .I(N__22974));
    InMux I__3309 (
            .O(N__23013),
            .I(N__22974));
    InMux I__3308 (
            .O(N__23010),
            .I(N__22974));
    InMux I__3307 (
            .O(N__23009),
            .I(N__22974));
    InMux I__3306 (
            .O(N__23006),
            .I(N__22974));
    InMux I__3305 (
            .O(N__23005),
            .I(N__22974));
    InMux I__3304 (
            .O(N__23002),
            .I(N__22974));
    InMux I__3303 (
            .O(N__22999),
            .I(N__22965));
    InMux I__3302 (
            .O(N__22998),
            .I(N__22965));
    InMux I__3301 (
            .O(N__22995),
            .I(N__22965));
    InMux I__3300 (
            .O(N__22994),
            .I(N__22965));
    Odrv4 I__3299 (
            .O(N__22991),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    LocalMux I__3298 (
            .O(N__22974),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    LocalMux I__3297 (
            .O(N__22965),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    CascadeMux I__3296 (
            .O(N__22958),
            .I(N__22955));
    InMux I__3295 (
            .O(N__22955),
            .I(N__22950));
    InMux I__3294 (
            .O(N__22954),
            .I(N__22947));
    InMux I__3293 (
            .O(N__22953),
            .I(N__22944));
    LocalMux I__3292 (
            .O(N__22950),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__3291 (
            .O(N__22947),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__3290 (
            .O(N__22944),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__3289 (
            .O(N__22937),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__3288 (
            .O(N__22934),
            .I(N__22929));
    InMux I__3287 (
            .O(N__22933),
            .I(N__22924));
    InMux I__3286 (
            .O(N__22932),
            .I(N__22924));
    LocalMux I__3285 (
            .O(N__22929),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__3284 (
            .O(N__22924),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__3283 (
            .O(N__22919),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__3282 (
            .O(N__22916),
            .I(N__22911));
    InMux I__3281 (
            .O(N__22915),
            .I(N__22906));
    InMux I__3280 (
            .O(N__22914),
            .I(N__22906));
    LocalMux I__3279 (
            .O(N__22911),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__3278 (
            .O(N__22906),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__3277 (
            .O(N__22901),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    CascadeMux I__3276 (
            .O(N__22898),
            .I(N__22894));
    CascadeMux I__3275 (
            .O(N__22897),
            .I(N__22891));
    InMux I__3274 (
            .O(N__22894),
            .I(N__22887));
    InMux I__3273 (
            .O(N__22891),
            .I(N__22884));
    InMux I__3272 (
            .O(N__22890),
            .I(N__22881));
    LocalMux I__3271 (
            .O(N__22887),
            .I(N__22878));
    LocalMux I__3270 (
            .O(N__22884),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__3269 (
            .O(N__22881),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__3268 (
            .O(N__22878),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__3267 (
            .O(N__22871),
            .I(bfn_8_22_0_));
    CascadeMux I__3266 (
            .O(N__22868),
            .I(N__22864));
    CascadeMux I__3265 (
            .O(N__22867),
            .I(N__22861));
    InMux I__3264 (
            .O(N__22864),
            .I(N__22857));
    InMux I__3263 (
            .O(N__22861),
            .I(N__22854));
    InMux I__3262 (
            .O(N__22860),
            .I(N__22851));
    LocalMux I__3261 (
            .O(N__22857),
            .I(N__22848));
    LocalMux I__3260 (
            .O(N__22854),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__3259 (
            .O(N__22851),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__3258 (
            .O(N__22848),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__3257 (
            .O(N__22841),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__3256 (
            .O(N__22838),
            .I(N__22835));
    InMux I__3255 (
            .O(N__22835),
            .I(N__22830));
    InMux I__3254 (
            .O(N__22834),
            .I(N__22827));
    InMux I__3253 (
            .O(N__22833),
            .I(N__22824));
    LocalMux I__3252 (
            .O(N__22830),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__3251 (
            .O(N__22827),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__3250 (
            .O(N__22824),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__3249 (
            .O(N__22817),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__3248 (
            .O(N__22814),
            .I(N__22811));
    InMux I__3247 (
            .O(N__22811),
            .I(N__22806));
    InMux I__3246 (
            .O(N__22810),
            .I(N__22803));
    InMux I__3245 (
            .O(N__22809),
            .I(N__22800));
    LocalMux I__3244 (
            .O(N__22806),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__3243 (
            .O(N__22803),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__3242 (
            .O(N__22800),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__3241 (
            .O(N__22793),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__3240 (
            .O(N__22790),
            .I(N__22786));
    InMux I__3239 (
            .O(N__22789),
            .I(N__22783));
    LocalMux I__3238 (
            .O(N__22786),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__3237 (
            .O(N__22783),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__3236 (
            .O(N__22778),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__3235 (
            .O(N__22775),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__3234 (
            .O(N__22772),
            .I(N__22768));
    InMux I__3233 (
            .O(N__22771),
            .I(N__22765));
    LocalMux I__3232 (
            .O(N__22768),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__3231 (
            .O(N__22765),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__3230 (
            .O(N__22760),
            .I(N__22757));
    InMux I__3229 (
            .O(N__22757),
            .I(N__22752));
    InMux I__3228 (
            .O(N__22756),
            .I(N__22749));
    InMux I__3227 (
            .O(N__22755),
            .I(N__22746));
    LocalMux I__3226 (
            .O(N__22752),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__3225 (
            .O(N__22749),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__3224 (
            .O(N__22746),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__3223 (
            .O(N__22739),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__3222 (
            .O(N__22736),
            .I(N__22731));
    InMux I__3221 (
            .O(N__22735),
            .I(N__22726));
    InMux I__3220 (
            .O(N__22734),
            .I(N__22726));
    LocalMux I__3219 (
            .O(N__22731),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__3218 (
            .O(N__22726),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__3217 (
            .O(N__22721),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__3216 (
            .O(N__22718),
            .I(N__22713));
    InMux I__3215 (
            .O(N__22717),
            .I(N__22708));
    InMux I__3214 (
            .O(N__22716),
            .I(N__22708));
    LocalMux I__3213 (
            .O(N__22713),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__3212 (
            .O(N__22708),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__3211 (
            .O(N__22703),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    CascadeMux I__3210 (
            .O(N__22700),
            .I(N__22696));
    CascadeMux I__3209 (
            .O(N__22699),
            .I(N__22693));
    InMux I__3208 (
            .O(N__22696),
            .I(N__22689));
    InMux I__3207 (
            .O(N__22693),
            .I(N__22686));
    InMux I__3206 (
            .O(N__22692),
            .I(N__22683));
    LocalMux I__3205 (
            .O(N__22689),
            .I(N__22680));
    LocalMux I__3204 (
            .O(N__22686),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__3203 (
            .O(N__22683),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__3202 (
            .O(N__22680),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__3201 (
            .O(N__22673),
            .I(bfn_8_21_0_));
    CascadeMux I__3200 (
            .O(N__22670),
            .I(N__22666));
    CascadeMux I__3199 (
            .O(N__22669),
            .I(N__22663));
    InMux I__3198 (
            .O(N__22666),
            .I(N__22659));
    InMux I__3197 (
            .O(N__22663),
            .I(N__22656));
    InMux I__3196 (
            .O(N__22662),
            .I(N__22653));
    LocalMux I__3195 (
            .O(N__22659),
            .I(N__22650));
    LocalMux I__3194 (
            .O(N__22656),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__3193 (
            .O(N__22653),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__3192 (
            .O(N__22650),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__3191 (
            .O(N__22643),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    CascadeMux I__3190 (
            .O(N__22640),
            .I(N__22637));
    InMux I__3189 (
            .O(N__22637),
            .I(N__22632));
    InMux I__3188 (
            .O(N__22636),
            .I(N__22629));
    InMux I__3187 (
            .O(N__22635),
            .I(N__22626));
    LocalMux I__3186 (
            .O(N__22632),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__3185 (
            .O(N__22629),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__3184 (
            .O(N__22626),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__3183 (
            .O(N__22619),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    CascadeMux I__3182 (
            .O(N__22616),
            .I(N__22613));
    InMux I__3181 (
            .O(N__22613),
            .I(N__22608));
    InMux I__3180 (
            .O(N__22612),
            .I(N__22605));
    InMux I__3179 (
            .O(N__22611),
            .I(N__22602));
    LocalMux I__3178 (
            .O(N__22608),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__3177 (
            .O(N__22605),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__3176 (
            .O(N__22602),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__3175 (
            .O(N__22595),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    CascadeMux I__3174 (
            .O(N__22592),
            .I(N__22589));
    InMux I__3173 (
            .O(N__22589),
            .I(N__22584));
    InMux I__3172 (
            .O(N__22588),
            .I(N__22581));
    InMux I__3171 (
            .O(N__22587),
            .I(N__22578));
    LocalMux I__3170 (
            .O(N__22584),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__3169 (
            .O(N__22581),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__3168 (
            .O(N__22578),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__3167 (
            .O(N__22571),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    CascadeMux I__3166 (
            .O(N__22568),
            .I(N__22565));
    InMux I__3165 (
            .O(N__22565),
            .I(N__22560));
    InMux I__3164 (
            .O(N__22564),
            .I(N__22557));
    InMux I__3163 (
            .O(N__22563),
            .I(N__22554));
    LocalMux I__3162 (
            .O(N__22560),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__3161 (
            .O(N__22557),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__3160 (
            .O(N__22554),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__3159 (
            .O(N__22547),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__3158 (
            .O(N__22544),
            .I(N__22539));
    InMux I__3157 (
            .O(N__22543),
            .I(N__22534));
    InMux I__3156 (
            .O(N__22542),
            .I(N__22534));
    LocalMux I__3155 (
            .O(N__22539),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__3154 (
            .O(N__22534),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__3153 (
            .O(N__22529),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__3152 (
            .O(N__22526),
            .I(N__22521));
    InMux I__3151 (
            .O(N__22525),
            .I(N__22516));
    InMux I__3150 (
            .O(N__22524),
            .I(N__22516));
    LocalMux I__3149 (
            .O(N__22521),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__3148 (
            .O(N__22516),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__3147 (
            .O(N__22511),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    CascadeMux I__3146 (
            .O(N__22508),
            .I(N__22505));
    InMux I__3145 (
            .O(N__22505),
            .I(N__22501));
    CascadeMux I__3144 (
            .O(N__22504),
            .I(N__22498));
    LocalMux I__3143 (
            .O(N__22501),
            .I(N__22494));
    InMux I__3142 (
            .O(N__22498),
            .I(N__22491));
    InMux I__3141 (
            .O(N__22497),
            .I(N__22488));
    Span4Mux_h I__3140 (
            .O(N__22494),
            .I(N__22485));
    LocalMux I__3139 (
            .O(N__22491),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__3138 (
            .O(N__22488),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__3137 (
            .O(N__22485),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__3136 (
            .O(N__22478),
            .I(bfn_8_20_0_));
    CascadeMux I__3135 (
            .O(N__22475),
            .I(N__22471));
    CascadeMux I__3134 (
            .O(N__22474),
            .I(N__22468));
    InMux I__3133 (
            .O(N__22471),
            .I(N__22464));
    InMux I__3132 (
            .O(N__22468),
            .I(N__22461));
    InMux I__3131 (
            .O(N__22467),
            .I(N__22458));
    LocalMux I__3130 (
            .O(N__22464),
            .I(N__22455));
    LocalMux I__3129 (
            .O(N__22461),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__3128 (
            .O(N__22458),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__3127 (
            .O(N__22455),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__3126 (
            .O(N__22448),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    CascadeMux I__3125 (
            .O(N__22445),
            .I(N__22442));
    InMux I__3124 (
            .O(N__22442),
            .I(N__22437));
    InMux I__3123 (
            .O(N__22441),
            .I(N__22434));
    InMux I__3122 (
            .O(N__22440),
            .I(N__22431));
    LocalMux I__3121 (
            .O(N__22437),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__3120 (
            .O(N__22434),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__3119 (
            .O(N__22431),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__3118 (
            .O(N__22424),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    CascadeMux I__3117 (
            .O(N__22421),
            .I(N__22418));
    InMux I__3116 (
            .O(N__22418),
            .I(N__22413));
    InMux I__3115 (
            .O(N__22417),
            .I(N__22410));
    InMux I__3114 (
            .O(N__22416),
            .I(N__22407));
    LocalMux I__3113 (
            .O(N__22413),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__3112 (
            .O(N__22410),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__3111 (
            .O(N__22407),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__3110 (
            .O(N__22400),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    CascadeMux I__3109 (
            .O(N__22397),
            .I(N__22394));
    InMux I__3108 (
            .O(N__22394),
            .I(N__22389));
    InMux I__3107 (
            .O(N__22393),
            .I(N__22386));
    InMux I__3106 (
            .O(N__22392),
            .I(N__22383));
    LocalMux I__3105 (
            .O(N__22389),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__3104 (
            .O(N__22386),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__3103 (
            .O(N__22383),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__3102 (
            .O(N__22376),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__3101 (
            .O(N__22373),
            .I(N__22369));
    InMux I__3100 (
            .O(N__22372),
            .I(N__22366));
    LocalMux I__3099 (
            .O(N__22369),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    LocalMux I__3098 (
            .O(N__22366),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__3097 (
            .O(N__22361),
            .I(N__22358));
    LocalMux I__3096 (
            .O(N__22358),
            .I(N__22354));
    InMux I__3095 (
            .O(N__22357),
            .I(N__22351));
    Odrv4 I__3094 (
            .O(N__22354),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    LocalMux I__3093 (
            .O(N__22351),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__3092 (
            .O(N__22346),
            .I(N__22343));
    LocalMux I__3091 (
            .O(N__22343),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16 ));
    InMux I__3090 (
            .O(N__22340),
            .I(N__22335));
    InMux I__3089 (
            .O(N__22339),
            .I(N__22330));
    InMux I__3088 (
            .O(N__22338),
            .I(N__22330));
    LocalMux I__3087 (
            .O(N__22335),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ));
    LocalMux I__3086 (
            .O(N__22330),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ));
    CascadeMux I__3085 (
            .O(N__22325),
            .I(N__22321));
    CascadeMux I__3084 (
            .O(N__22324),
            .I(N__22318));
    InMux I__3083 (
            .O(N__22321),
            .I(N__22314));
    InMux I__3082 (
            .O(N__22318),
            .I(N__22309));
    InMux I__3081 (
            .O(N__22317),
            .I(N__22309));
    LocalMux I__3080 (
            .O(N__22314),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ));
    LocalMux I__3079 (
            .O(N__22309),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ));
    InMux I__3078 (
            .O(N__22304),
            .I(N__22301));
    LocalMux I__3077 (
            .O(N__22301),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15 ));
    InMux I__3076 (
            .O(N__22298),
            .I(N__22295));
    LocalMux I__3075 (
            .O(N__22295),
            .I(N__22291));
    InMux I__3074 (
            .O(N__22294),
            .I(N__22288));
    Odrv4 I__3073 (
            .O(N__22291),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ));
    LocalMux I__3072 (
            .O(N__22288),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ));
    CascadeMux I__3071 (
            .O(N__22283),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_ ));
    CascadeMux I__3070 (
            .O(N__22280),
            .I(N__22277));
    InMux I__3069 (
            .O(N__22277),
            .I(N__22273));
    InMux I__3068 (
            .O(N__22276),
            .I(N__22270));
    LocalMux I__3067 (
            .O(N__22273),
            .I(N__22266));
    LocalMux I__3066 (
            .O(N__22270),
            .I(N__22263));
    InMux I__3065 (
            .O(N__22269),
            .I(N__22260));
    Odrv4 I__3064 (
            .O(N__22266),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ));
    Odrv4 I__3063 (
            .O(N__22263),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ));
    LocalMux I__3062 (
            .O(N__22260),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ));
    InMux I__3061 (
            .O(N__22253),
            .I(bfn_8_19_0_));
    InMux I__3060 (
            .O(N__22250),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    CascadeMux I__3059 (
            .O(N__22247),
            .I(N__22244));
    InMux I__3058 (
            .O(N__22244),
            .I(N__22239));
    InMux I__3057 (
            .O(N__22243),
            .I(N__22236));
    InMux I__3056 (
            .O(N__22242),
            .I(N__22233));
    LocalMux I__3055 (
            .O(N__22239),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__3054 (
            .O(N__22236),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__3053 (
            .O(N__22233),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__3052 (
            .O(N__22226),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    CascadeMux I__3051 (
            .O(N__22223),
            .I(N__22220));
    InMux I__3050 (
            .O(N__22220),
            .I(N__22215));
    InMux I__3049 (
            .O(N__22219),
            .I(N__22212));
    InMux I__3048 (
            .O(N__22218),
            .I(N__22209));
    LocalMux I__3047 (
            .O(N__22215),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__3046 (
            .O(N__22212),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__3045 (
            .O(N__22209),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__3044 (
            .O(N__22202),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    CascadeMux I__3043 (
            .O(N__22199),
            .I(N__22196));
    InMux I__3042 (
            .O(N__22196),
            .I(N__22191));
    InMux I__3041 (
            .O(N__22195),
            .I(N__22188));
    InMux I__3040 (
            .O(N__22194),
            .I(N__22185));
    LocalMux I__3039 (
            .O(N__22191),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__3038 (
            .O(N__22188),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__3037 (
            .O(N__22185),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__3036 (
            .O(N__22178),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__3035 (
            .O(N__22175),
            .I(N__22172));
    LocalMux I__3034 (
            .O(N__22172),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31 ));
    CascadeMux I__3033 (
            .O(N__22169),
            .I(N__22166));
    InMux I__3032 (
            .O(N__22166),
            .I(N__22163));
    LocalMux I__3031 (
            .O(N__22163),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5 ));
    InMux I__3030 (
            .O(N__22160),
            .I(N__22157));
    LocalMux I__3029 (
            .O(N__22157),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6 ));
    CascadeMux I__3028 (
            .O(N__22154),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_ ));
    InMux I__3027 (
            .O(N__22151),
            .I(N__22147));
    InMux I__3026 (
            .O(N__22150),
            .I(N__22144));
    LocalMux I__3025 (
            .O(N__22147),
            .I(N__22141));
    LocalMux I__3024 (
            .O(N__22144),
            .I(N__22138));
    Span4Mux_v I__3023 (
            .O(N__22141),
            .I(N__22134));
    Span4Mux_h I__3022 (
            .O(N__22138),
            .I(N__22131));
    InMux I__3021 (
            .O(N__22137),
            .I(N__22128));
    Odrv4 I__3020 (
            .O(N__22134),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv4 I__3019 (
            .O(N__22131),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    LocalMux I__3018 (
            .O(N__22128),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__3017 (
            .O(N__22121),
            .I(N__22115));
    InMux I__3016 (
            .O(N__22120),
            .I(N__22115));
    LocalMux I__3015 (
            .O(N__22115),
            .I(N__22111));
    InMux I__3014 (
            .O(N__22114),
            .I(N__22108));
    Span4Mux_v I__3013 (
            .O(N__22111),
            .I(N__22105));
    LocalMux I__3012 (
            .O(N__22108),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    Odrv4 I__3011 (
            .O(N__22105),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__3010 (
            .O(N__22100),
            .I(N__22095));
    CascadeMux I__3009 (
            .O(N__22099),
            .I(N__22092));
    CascadeMux I__3008 (
            .O(N__22098),
            .I(N__22089));
    LocalMux I__3007 (
            .O(N__22095),
            .I(N__22086));
    InMux I__3006 (
            .O(N__22092),
            .I(N__22083));
    InMux I__3005 (
            .O(N__22089),
            .I(N__22080));
    Span4Mux_v I__3004 (
            .O(N__22086),
            .I(N__22075));
    LocalMux I__3003 (
            .O(N__22083),
            .I(N__22075));
    LocalMux I__3002 (
            .O(N__22080),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__3001 (
            .O(N__22075),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__3000 (
            .O(N__22070),
            .I(N__22066));
    InMux I__2999 (
            .O(N__22069),
            .I(N__22062));
    LocalMux I__2998 (
            .O(N__22066),
            .I(N__22058));
    InMux I__2997 (
            .O(N__22065),
            .I(N__22055));
    LocalMux I__2996 (
            .O(N__22062),
            .I(N__22052));
    InMux I__2995 (
            .O(N__22061),
            .I(N__22049));
    Odrv12 I__2994 (
            .O(N__22058),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    LocalMux I__2993 (
            .O(N__22055),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    Odrv4 I__2992 (
            .O(N__22052),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    LocalMux I__2991 (
            .O(N__22049),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    InMux I__2990 (
            .O(N__22040),
            .I(N__22037));
    LocalMux I__2989 (
            .O(N__22037),
            .I(N__22031));
    InMux I__2988 (
            .O(N__22036),
            .I(N__22028));
    InMux I__2987 (
            .O(N__22035),
            .I(N__22025));
    InMux I__2986 (
            .O(N__22034),
            .I(N__22022));
    Span4Mux_v I__2985 (
            .O(N__22031),
            .I(N__22015));
    LocalMux I__2984 (
            .O(N__22028),
            .I(N__22015));
    LocalMux I__2983 (
            .O(N__22025),
            .I(N__22015));
    LocalMux I__2982 (
            .O(N__22022),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ));
    Odrv4 I__2981 (
            .O(N__22015),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ));
    CascadeMux I__2980 (
            .O(N__22010),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_ ));
    CascadeMux I__2979 (
            .O(N__22007),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_ ));
    CascadeMux I__2978 (
            .O(N__22004),
            .I(N__22000));
    InMux I__2977 (
            .O(N__22003),
            .I(N__21997));
    InMux I__2976 (
            .O(N__22000),
            .I(N__21994));
    LocalMux I__2975 (
            .O(N__21997),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ));
    LocalMux I__2974 (
            .O(N__21994),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ));
    CascadeMux I__2973 (
            .O(N__21989),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_ ));
    InMux I__2972 (
            .O(N__21986),
            .I(N__21983));
    LocalMux I__2971 (
            .O(N__21983),
            .I(N__21980));
    Odrv4 I__2970 (
            .O(N__21980),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24 ));
    CascadeMux I__2969 (
            .O(N__21977),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_ ));
    InMux I__2968 (
            .O(N__21974),
            .I(N__21971));
    LocalMux I__2967 (
            .O(N__21971),
            .I(N__21968));
    Odrv12 I__2966 (
            .O(N__21968),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17 ));
    CascadeMux I__2965 (
            .O(N__21965),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_ ));
    CascadeMux I__2964 (
            .O(N__21962),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31_cascade_ ));
    CascadeMux I__2963 (
            .O(N__21959),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31_cascade_ ));
    InMux I__2962 (
            .O(N__21956),
            .I(N__21953));
    LocalMux I__2961 (
            .O(N__21953),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2 ));
    InMux I__2960 (
            .O(N__21950),
            .I(N__21947));
    LocalMux I__2959 (
            .O(N__21947),
            .I(N__21944));
    Span4Mux_v I__2958 (
            .O(N__21944),
            .I(N__21941));
    Odrv4 I__2957 (
            .O(N__21941),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14 ));
    CascadeMux I__2956 (
            .O(N__21938),
            .I(N__21935));
    InMux I__2955 (
            .O(N__21935),
            .I(N__21931));
    InMux I__2954 (
            .O(N__21934),
            .I(N__21926));
    LocalMux I__2953 (
            .O(N__21931),
            .I(N__21923));
    InMux I__2952 (
            .O(N__21930),
            .I(N__21917));
    InMux I__2951 (
            .O(N__21929),
            .I(N__21917));
    LocalMux I__2950 (
            .O(N__21926),
            .I(N__21912));
    Span12Mux_s8_h I__2949 (
            .O(N__21923),
            .I(N__21912));
    InMux I__2948 (
            .O(N__21922),
            .I(N__21909));
    LocalMux I__2947 (
            .O(N__21917),
            .I(N__21906));
    Odrv12 I__2946 (
            .O(N__21912),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    LocalMux I__2945 (
            .O(N__21909),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    Odrv4 I__2944 (
            .O(N__21906),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    CascadeMux I__2943 (
            .O(N__21899),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14_cascade_));
    InMux I__2942 (
            .O(N__21896),
            .I(N__21892));
    InMux I__2941 (
            .O(N__21895),
            .I(N__21889));
    LocalMux I__2940 (
            .O(N__21892),
            .I(N__21882));
    LocalMux I__2939 (
            .O(N__21889),
            .I(N__21882));
    InMux I__2938 (
            .O(N__21888),
            .I(N__21879));
    InMux I__2937 (
            .O(N__21887),
            .I(N__21876));
    Odrv4 I__2936 (
            .O(N__21882),
            .I(elapsed_time_ns_1_RNIL13KD1_0_9));
    LocalMux I__2935 (
            .O(N__21879),
            .I(elapsed_time_ns_1_RNIL13KD1_0_9));
    LocalMux I__2934 (
            .O(N__21876),
            .I(elapsed_time_ns_1_RNIL13KD1_0_9));
    InMux I__2933 (
            .O(N__21869),
            .I(N__21865));
    InMux I__2932 (
            .O(N__21868),
            .I(N__21862));
    LocalMux I__2931 (
            .O(N__21865),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_1Z0Z_9 ));
    LocalMux I__2930 (
            .O(N__21862),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_1Z0Z_9 ));
    CascadeMux I__2929 (
            .O(N__21857),
            .I(N__21853));
    InMux I__2928 (
            .O(N__21856),
            .I(N__21850));
    InMux I__2927 (
            .O(N__21853),
            .I(N__21846));
    LocalMux I__2926 (
            .O(N__21850),
            .I(N__21843));
    InMux I__2925 (
            .O(N__21849),
            .I(N__21840));
    LocalMux I__2924 (
            .O(N__21846),
            .I(elapsed_time_ns_1_RNINVLD11_0_10));
    Odrv4 I__2923 (
            .O(N__21843),
            .I(elapsed_time_ns_1_RNINVLD11_0_10));
    LocalMux I__2922 (
            .O(N__21840),
            .I(elapsed_time_ns_1_RNINVLD11_0_10));
    CascadeMux I__2921 (
            .O(N__21833),
            .I(N__21827));
    CascadeMux I__2920 (
            .O(N__21832),
            .I(N__21820));
    CascadeMux I__2919 (
            .O(N__21831),
            .I(N__21817));
    InMux I__2918 (
            .O(N__21830),
            .I(N__21811));
    InMux I__2917 (
            .O(N__21827),
            .I(N__21811));
    InMux I__2916 (
            .O(N__21826),
            .I(N__21806));
    InMux I__2915 (
            .O(N__21825),
            .I(N__21806));
    InMux I__2914 (
            .O(N__21824),
            .I(N__21801));
    InMux I__2913 (
            .O(N__21823),
            .I(N__21801));
    InMux I__2912 (
            .O(N__21820),
            .I(N__21796));
    InMux I__2911 (
            .O(N__21817),
            .I(N__21796));
    InMux I__2910 (
            .O(N__21816),
            .I(N__21793));
    LocalMux I__2909 (
            .O(N__21811),
            .I(\phase_controller_inst1.stoper_hc.N_315 ));
    LocalMux I__2908 (
            .O(N__21806),
            .I(\phase_controller_inst1.stoper_hc.N_315 ));
    LocalMux I__2907 (
            .O(N__21801),
            .I(\phase_controller_inst1.stoper_hc.N_315 ));
    LocalMux I__2906 (
            .O(N__21796),
            .I(\phase_controller_inst1.stoper_hc.N_315 ));
    LocalMux I__2905 (
            .O(N__21793),
            .I(\phase_controller_inst1.stoper_hc.N_315 ));
    InMux I__2904 (
            .O(N__21782),
            .I(N__21778));
    InMux I__2903 (
            .O(N__21781),
            .I(N__21773));
    LocalMux I__2902 (
            .O(N__21778),
            .I(N__21770));
    InMux I__2901 (
            .O(N__21777),
            .I(N__21765));
    InMux I__2900 (
            .O(N__21776),
            .I(N__21765));
    LocalMux I__2899 (
            .O(N__21773),
            .I(elapsed_time_ns_1_RNIO0MD11_0_11));
    Odrv4 I__2898 (
            .O(N__21770),
            .I(elapsed_time_ns_1_RNIO0MD11_0_11));
    LocalMux I__2897 (
            .O(N__21765),
            .I(elapsed_time_ns_1_RNIO0MD11_0_11));
    InMux I__2896 (
            .O(N__21758),
            .I(N__21754));
    InMux I__2895 (
            .O(N__21757),
            .I(N__21751));
    LocalMux I__2894 (
            .O(N__21754),
            .I(elapsed_time_ns_1_RNIR4ND11_0_23));
    LocalMux I__2893 (
            .O(N__21751),
            .I(elapsed_time_ns_1_RNIR4ND11_0_23));
    InMux I__2892 (
            .O(N__21746),
            .I(N__21742));
    InMux I__2891 (
            .O(N__21745),
            .I(N__21739));
    LocalMux I__2890 (
            .O(N__21742),
            .I(N__21734));
    LocalMux I__2889 (
            .O(N__21739),
            .I(N__21734));
    Odrv4 I__2888 (
            .O(N__21734),
            .I(elapsed_time_ns_1_RNIS5ND11_0_24));
    CascadeMux I__2887 (
            .O(N__21731),
            .I(N__21728));
    InMux I__2886 (
            .O(N__21728),
            .I(N__21724));
    CascadeMux I__2885 (
            .O(N__21727),
            .I(N__21721));
    LocalMux I__2884 (
            .O(N__21724),
            .I(N__21718));
    InMux I__2883 (
            .O(N__21721),
            .I(N__21715));
    Span4Mux_h I__2882 (
            .O(N__21718),
            .I(N__21712));
    LocalMux I__2881 (
            .O(N__21715),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    Odrv4 I__2880 (
            .O(N__21712),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2879 (
            .O(N__21707),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__2878 (
            .O(N__21704),
            .I(N__21701));
    LocalMux I__2877 (
            .O(N__21701),
            .I(N__21697));
    InMux I__2876 (
            .O(N__21700),
            .I(N__21694));
    Span4Mux_v I__2875 (
            .O(N__21697),
            .I(N__21691));
    LocalMux I__2874 (
            .O(N__21694),
            .I(N__21688));
    Odrv4 I__2873 (
            .O(N__21691),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    Odrv4 I__2872 (
            .O(N__21688),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2871 (
            .O(N__21683),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2870 (
            .O(N__21680),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2869 (
            .O(N__21677),
            .I(N__21674));
    LocalMux I__2868 (
            .O(N__21674),
            .I(N__21667));
    InMux I__2867 (
            .O(N__21673),
            .I(N__21664));
    InMux I__2866 (
            .O(N__21672),
            .I(N__21656));
    InMux I__2865 (
            .O(N__21671),
            .I(N__21656));
    InMux I__2864 (
            .O(N__21670),
            .I(N__21653));
    Span4Mux_v I__2863 (
            .O(N__21667),
            .I(N__21646));
    LocalMux I__2862 (
            .O(N__21664),
            .I(N__21646));
    InMux I__2861 (
            .O(N__21663),
            .I(N__21643));
    InMux I__2860 (
            .O(N__21662),
            .I(N__21638));
    InMux I__2859 (
            .O(N__21661),
            .I(N__21638));
    LocalMux I__2858 (
            .O(N__21656),
            .I(N__21635));
    LocalMux I__2857 (
            .O(N__21653),
            .I(N__21632));
    InMux I__2856 (
            .O(N__21652),
            .I(N__21627));
    InMux I__2855 (
            .O(N__21651),
            .I(N__21627));
    Span4Mux_v I__2854 (
            .O(N__21646),
            .I(N__21624));
    LocalMux I__2853 (
            .O(N__21643),
            .I(N__21619));
    LocalMux I__2852 (
            .O(N__21638),
            .I(N__21619));
    Span4Mux_v I__2851 (
            .O(N__21635),
            .I(N__21616));
    Span12Mux_s8_h I__2850 (
            .O(N__21632),
            .I(N__21613));
    LocalMux I__2849 (
            .O(N__21627),
            .I(N__21610));
    Span4Mux_h I__2848 (
            .O(N__21624),
            .I(N__21605));
    Span4Mux_v I__2847 (
            .O(N__21619),
            .I(N__21605));
    Span4Mux_h I__2846 (
            .O(N__21616),
            .I(N__21602));
    Odrv12 I__2845 (
            .O(N__21613),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv12 I__2844 (
            .O(N__21610),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2843 (
            .O(N__21605),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2842 (
            .O(N__21602),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__2841 (
            .O(N__21593),
            .I(N__21590));
    LocalMux I__2840 (
            .O(N__21590),
            .I(N__21586));
    InMux I__2839 (
            .O(N__21589),
            .I(N__21583));
    Odrv12 I__2838 (
            .O(N__21586),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_14 ));
    LocalMux I__2837 (
            .O(N__21583),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_14 ));
    InMux I__2836 (
            .O(N__21578),
            .I(N__21572));
    InMux I__2835 (
            .O(N__21577),
            .I(N__21572));
    LocalMux I__2834 (
            .O(N__21572),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2833 (
            .O(N__21569),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    CascadeMux I__2832 (
            .O(N__21566),
            .I(N__21563));
    InMux I__2831 (
            .O(N__21563),
            .I(N__21560));
    LocalMux I__2830 (
            .O(N__21560),
            .I(N__21556));
    InMux I__2829 (
            .O(N__21559),
            .I(N__21553));
    Odrv12 I__2828 (
            .O(N__21556),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    LocalMux I__2827 (
            .O(N__21553),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2826 (
            .O(N__21548),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2825 (
            .O(N__21545),
            .I(N__21542));
    LocalMux I__2824 (
            .O(N__21542),
            .I(N__21538));
    InMux I__2823 (
            .O(N__21541),
            .I(N__21535));
    Odrv4 I__2822 (
            .O(N__21538),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    LocalMux I__2821 (
            .O(N__21535),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2820 (
            .O(N__21530),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2819 (
            .O(N__21527),
            .I(N__21521));
    InMux I__2818 (
            .O(N__21526),
            .I(N__21521));
    LocalMux I__2817 (
            .O(N__21521),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2816 (
            .O(N__21518),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    CascadeMux I__2815 (
            .O(N__21515),
            .I(N__21512));
    InMux I__2814 (
            .O(N__21512),
            .I(N__21508));
    InMux I__2813 (
            .O(N__21511),
            .I(N__21505));
    LocalMux I__2812 (
            .O(N__21508),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    LocalMux I__2811 (
            .O(N__21505),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2810 (
            .O(N__21500),
            .I(bfn_8_13_0_));
    CascadeMux I__2809 (
            .O(N__21497),
            .I(N__21494));
    InMux I__2808 (
            .O(N__21494),
            .I(N__21488));
    InMux I__2807 (
            .O(N__21493),
            .I(N__21488));
    LocalMux I__2806 (
            .O(N__21488),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2805 (
            .O(N__21485),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    InMux I__2804 (
            .O(N__21482),
            .I(N__21479));
    LocalMux I__2803 (
            .O(N__21479),
            .I(N__21475));
    InMux I__2802 (
            .O(N__21478),
            .I(N__21472));
    Span4Mux_h I__2801 (
            .O(N__21475),
            .I(N__21469));
    LocalMux I__2800 (
            .O(N__21472),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    Odrv4 I__2799 (
            .O(N__21469),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2798 (
            .O(N__21464),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2797 (
            .O(N__21461),
            .I(N__21457));
    InMux I__2796 (
            .O(N__21460),
            .I(N__21454));
    LocalMux I__2795 (
            .O(N__21457),
            .I(N__21451));
    LocalMux I__2794 (
            .O(N__21454),
            .I(N__21448));
    Span4Mux_h I__2793 (
            .O(N__21451),
            .I(N__21445));
    Odrv4 I__2792 (
            .O(N__21448),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    Odrv4 I__2791 (
            .O(N__21445),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2790 (
            .O(N__21440),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2789 (
            .O(N__21437),
            .I(N__21434));
    LocalMux I__2788 (
            .O(N__21434),
            .I(N__21431));
    Span4Mux_v I__2787 (
            .O(N__21431),
            .I(N__21427));
    InMux I__2786 (
            .O(N__21430),
            .I(N__21424));
    Odrv4 I__2785 (
            .O(N__21427),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    LocalMux I__2784 (
            .O(N__21424),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2783 (
            .O(N__21419),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    CascadeMux I__2782 (
            .O(N__21416),
            .I(N__21413));
    InMux I__2781 (
            .O(N__21413),
            .I(N__21410));
    LocalMux I__2780 (
            .O(N__21410),
            .I(N__21406));
    InMux I__2779 (
            .O(N__21409),
            .I(N__21403));
    Odrv12 I__2778 (
            .O(N__21406),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    LocalMux I__2777 (
            .O(N__21403),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2776 (
            .O(N__21398),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2775 (
            .O(N__21395),
            .I(N__21389));
    InMux I__2774 (
            .O(N__21394),
            .I(N__21389));
    LocalMux I__2773 (
            .O(N__21389),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2772 (
            .O(N__21386),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    CascadeMux I__2771 (
            .O(N__21383),
            .I(N__21379));
    InMux I__2770 (
            .O(N__21382),
            .I(N__21376));
    InMux I__2769 (
            .O(N__21379),
            .I(N__21373));
    LocalMux I__2768 (
            .O(N__21376),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    LocalMux I__2767 (
            .O(N__21373),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2766 (
            .O(N__21368),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2765 (
            .O(N__21365),
            .I(N__21362));
    LocalMux I__2764 (
            .O(N__21362),
            .I(N__21359));
    Span4Mux_h I__2763 (
            .O(N__21359),
            .I(N__21355));
    InMux I__2762 (
            .O(N__21358),
            .I(N__21352));
    Odrv4 I__2761 (
            .O(N__21355),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__2760 (
            .O(N__21352),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2759 (
            .O(N__21347),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    CascadeMux I__2758 (
            .O(N__21344),
            .I(N__21341));
    InMux I__2757 (
            .O(N__21341),
            .I(N__21338));
    LocalMux I__2756 (
            .O(N__21338),
            .I(N__21334));
    InMux I__2755 (
            .O(N__21337),
            .I(N__21331));
    Odrv12 I__2754 (
            .O(N__21334),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    LocalMux I__2753 (
            .O(N__21331),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2752 (
            .O(N__21326),
            .I(bfn_8_12_0_));
    InMux I__2751 (
            .O(N__21323),
            .I(N__21317));
    InMux I__2750 (
            .O(N__21322),
            .I(N__21317));
    LocalMux I__2749 (
            .O(N__21317),
            .I(N__21314));
    Odrv12 I__2748 (
            .O(N__21314),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2747 (
            .O(N__21311),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    CascadeMux I__2746 (
            .O(N__21308),
            .I(N__21305));
    InMux I__2745 (
            .O(N__21305),
            .I(N__21299));
    InMux I__2744 (
            .O(N__21304),
            .I(N__21299));
    LocalMux I__2743 (
            .O(N__21299),
            .I(N__21296));
    Span4Mux_v I__2742 (
            .O(N__21296),
            .I(N__21293));
    Odrv4 I__2741 (
            .O(N__21293),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2740 (
            .O(N__21290),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2739 (
            .O(N__21287),
            .I(N__21281));
    InMux I__2738 (
            .O(N__21286),
            .I(N__21281));
    LocalMux I__2737 (
            .O(N__21281),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2736 (
            .O(N__21278),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    CascadeMux I__2735 (
            .O(N__21275),
            .I(N__21271));
    InMux I__2734 (
            .O(N__21274),
            .I(N__21268));
    InMux I__2733 (
            .O(N__21271),
            .I(N__21265));
    LocalMux I__2732 (
            .O(N__21268),
            .I(N__21262));
    LocalMux I__2731 (
            .O(N__21265),
            .I(N__21259));
    Span4Mux_v I__2730 (
            .O(N__21262),
            .I(N__21256));
    Span12Mux_v I__2729 (
            .O(N__21259),
            .I(N__21250));
    Sp12to4 I__2728 (
            .O(N__21256),
            .I(N__21250));
    InMux I__2727 (
            .O(N__21255),
            .I(N__21247));
    Odrv12 I__2726 (
            .O(N__21250),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    LocalMux I__2725 (
            .O(N__21247),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2724 (
            .O(N__21242),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__2723 (
            .O(N__21239),
            .I(N__21235));
    InMux I__2722 (
            .O(N__21238),
            .I(N__21231));
    LocalMux I__2721 (
            .O(N__21235),
            .I(N__21228));
    InMux I__2720 (
            .O(N__21234),
            .I(N__21225));
    LocalMux I__2719 (
            .O(N__21231),
            .I(N__21220));
    Span4Mux_h I__2718 (
            .O(N__21228),
            .I(N__21220));
    LocalMux I__2717 (
            .O(N__21225),
            .I(N__21216));
    Span4Mux_h I__2716 (
            .O(N__21220),
            .I(N__21213));
    InMux I__2715 (
            .O(N__21219),
            .I(N__21210));
    Odrv12 I__2714 (
            .O(N__21216),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2713 (
            .O(N__21213),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    LocalMux I__2712 (
            .O(N__21210),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2711 (
            .O(N__21203),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    CascadeMux I__2710 (
            .O(N__21200),
            .I(N__21197));
    InMux I__2709 (
            .O(N__21197),
            .I(N__21194));
    LocalMux I__2708 (
            .O(N__21194),
            .I(N__21189));
    InMux I__2707 (
            .O(N__21193),
            .I(N__21186));
    InMux I__2706 (
            .O(N__21192),
            .I(N__21183));
    Span4Mux_v I__2705 (
            .O(N__21189),
            .I(N__21180));
    LocalMux I__2704 (
            .O(N__21186),
            .I(N__21175));
    LocalMux I__2703 (
            .O(N__21183),
            .I(N__21175));
    Span4Mux_h I__2702 (
            .O(N__21180),
            .I(N__21170));
    Span4Mux_v I__2701 (
            .O(N__21175),
            .I(N__21170));
    Odrv4 I__2700 (
            .O(N__21170),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2699 (
            .O(N__21167),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    CascadeMux I__2698 (
            .O(N__21164),
            .I(N__21161));
    InMux I__2697 (
            .O(N__21161),
            .I(N__21158));
    LocalMux I__2696 (
            .O(N__21158),
            .I(N__21154));
    InMux I__2695 (
            .O(N__21157),
            .I(N__21151));
    Span4Mux_h I__2694 (
            .O(N__21154),
            .I(N__21145));
    LocalMux I__2693 (
            .O(N__21151),
            .I(N__21145));
    InMux I__2692 (
            .O(N__21150),
            .I(N__21142));
    Span4Mux_v I__2691 (
            .O(N__21145),
            .I(N__21137));
    LocalMux I__2690 (
            .O(N__21142),
            .I(N__21137));
    Span4Mux_h I__2689 (
            .O(N__21137),
            .I(N__21134));
    Odrv4 I__2688 (
            .O(N__21134),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2687 (
            .O(N__21131),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    CascadeMux I__2686 (
            .O(N__21128),
            .I(N__21123));
    InMux I__2685 (
            .O(N__21127),
            .I(N__21120));
    InMux I__2684 (
            .O(N__21126),
            .I(N__21117));
    InMux I__2683 (
            .O(N__21123),
            .I(N__21114));
    LocalMux I__2682 (
            .O(N__21120),
            .I(N__21109));
    LocalMux I__2681 (
            .O(N__21117),
            .I(N__21109));
    LocalMux I__2680 (
            .O(N__21114),
            .I(N__21106));
    Span4Mux_v I__2679 (
            .O(N__21109),
            .I(N__21103));
    Odrv12 I__2678 (
            .O(N__21106),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__2677 (
            .O(N__21103),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2676 (
            .O(N__21098),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    CascadeMux I__2675 (
            .O(N__21095),
            .I(N__21092));
    InMux I__2674 (
            .O(N__21092),
            .I(N__21088));
    InMux I__2673 (
            .O(N__21091),
            .I(N__21085));
    LocalMux I__2672 (
            .O(N__21088),
            .I(N__21081));
    LocalMux I__2671 (
            .O(N__21085),
            .I(N__21078));
    InMux I__2670 (
            .O(N__21084),
            .I(N__21075));
    Span4Mux_h I__2669 (
            .O(N__21081),
            .I(N__21072));
    Span4Mux_v I__2668 (
            .O(N__21078),
            .I(N__21067));
    LocalMux I__2667 (
            .O(N__21075),
            .I(N__21067));
    Span4Mux_h I__2666 (
            .O(N__21072),
            .I(N__21064));
    Span4Mux_h I__2665 (
            .O(N__21067),
            .I(N__21061));
    Odrv4 I__2664 (
            .O(N__21064),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2663 (
            .O(N__21061),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2662 (
            .O(N__21056),
            .I(bfn_8_11_0_));
    InMux I__2661 (
            .O(N__21053),
            .I(N__21050));
    LocalMux I__2660 (
            .O(N__21050),
            .I(N__21045));
    InMux I__2659 (
            .O(N__21049),
            .I(N__21042));
    InMux I__2658 (
            .O(N__21048),
            .I(N__21039));
    Span4Mux_h I__2657 (
            .O(N__21045),
            .I(N__21034));
    LocalMux I__2656 (
            .O(N__21042),
            .I(N__21034));
    LocalMux I__2655 (
            .O(N__21039),
            .I(N__21031));
    Span4Mux_h I__2654 (
            .O(N__21034),
            .I(N__21028));
    Odrv12 I__2653 (
            .O(N__21031),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv4 I__2652 (
            .O(N__21028),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2651 (
            .O(N__21023),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    InMux I__2650 (
            .O(N__21020),
            .I(N__21014));
    InMux I__2649 (
            .O(N__21019),
            .I(N__21014));
    LocalMux I__2648 (
            .O(N__21014),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2647 (
            .O(N__21011),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2646 (
            .O(N__21008),
            .I(N__21005));
    LocalMux I__2645 (
            .O(N__21005),
            .I(N__21001));
    InMux I__2644 (
            .O(N__21004),
            .I(N__20998));
    Odrv4 I__2643 (
            .O(N__21001),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    LocalMux I__2642 (
            .O(N__20998),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2641 (
            .O(N__20993),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2640 (
            .O(N__20990),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__2639 (
            .O(N__20987),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__2638 (
            .O(N__20984),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__2637 (
            .O(N__20981),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__2636 (
            .O(N__20978),
            .I(N__20975));
    LocalMux I__2635 (
            .O(N__20975),
            .I(N__20972));
    Span4Mux_h I__2634 (
            .O(N__20972),
            .I(N__20969));
    Span4Mux_v I__2633 (
            .O(N__20969),
            .I(N__20966));
    Odrv4 I__2632 (
            .O(N__20966),
            .I(il_min_comp2_c));
    InMux I__2631 (
            .O(N__20963),
            .I(N__20960));
    LocalMux I__2630 (
            .O(N__20960),
            .I(N__20957));
    Span4Mux_h I__2629 (
            .O(N__20957),
            .I(N__20954));
    Span4Mux_h I__2628 (
            .O(N__20954),
            .I(N__20951));
    Odrv4 I__2627 (
            .O(N__20951),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__2626 (
            .O(N__20948),
            .I(N__20945));
    LocalMux I__2625 (
            .O(N__20945),
            .I(N__20942));
    Span4Mux_h I__2624 (
            .O(N__20942),
            .I(N__20939));
    Span4Mux_h I__2623 (
            .O(N__20939),
            .I(N__20936));
    Odrv4 I__2622 (
            .O(N__20936),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2621 (
            .O(N__20933),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    CascadeMux I__2620 (
            .O(N__20930),
            .I(N__20927));
    InMux I__2619 (
            .O(N__20927),
            .I(N__20924));
    LocalMux I__2618 (
            .O(N__20924),
            .I(N__20921));
    Span12Mux_s8_h I__2617 (
            .O(N__20921),
            .I(N__20918));
    Odrv12 I__2616 (
            .O(N__20918),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2615 (
            .O(N__20915),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2614 (
            .O(N__20912),
            .I(bfn_7_20_0_));
    InMux I__2613 (
            .O(N__20909),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__2612 (
            .O(N__20906),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__2611 (
            .O(N__20903),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__2610 (
            .O(N__20900),
            .I(N__20897));
    InMux I__2609 (
            .O(N__20897),
            .I(N__20894));
    LocalMux I__2608 (
            .O(N__20894),
            .I(N__20890));
    InMux I__2607 (
            .O(N__20893),
            .I(N__20887));
    Span4Mux_v I__2606 (
            .O(N__20890),
            .I(N__20882));
    LocalMux I__2605 (
            .O(N__20887),
            .I(N__20882));
    Odrv4 I__2604 (
            .O(N__20882),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__2603 (
            .O(N__20879),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__2602 (
            .O(N__20876),
            .I(N__20873));
    LocalMux I__2601 (
            .O(N__20873),
            .I(N__20869));
    InMux I__2600 (
            .O(N__20872),
            .I(N__20866));
    Span4Mux_h I__2599 (
            .O(N__20869),
            .I(N__20861));
    LocalMux I__2598 (
            .O(N__20866),
            .I(N__20861));
    Odrv4 I__2597 (
            .O(N__20861),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__2596 (
            .O(N__20858),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__2595 (
            .O(N__20855),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__2594 (
            .O(N__20852),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__2593 (
            .O(N__20849),
            .I(bfn_7_21_0_));
    CascadeMux I__2592 (
            .O(N__20846),
            .I(N__20843));
    InMux I__2591 (
            .O(N__20843),
            .I(N__20840));
    LocalMux I__2590 (
            .O(N__20840),
            .I(N__20836));
    InMux I__2589 (
            .O(N__20839),
            .I(N__20833));
    Odrv12 I__2588 (
            .O(N__20836),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__2587 (
            .O(N__20833),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__2586 (
            .O(N__20828),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__2585 (
            .O(N__20825),
            .I(N__20822));
    InMux I__2584 (
            .O(N__20822),
            .I(N__20819));
    LocalMux I__2583 (
            .O(N__20819),
            .I(N__20815));
    InMux I__2582 (
            .O(N__20818),
            .I(N__20812));
    Span4Mux_h I__2581 (
            .O(N__20815),
            .I(N__20809));
    LocalMux I__2580 (
            .O(N__20812),
            .I(N__20806));
    Odrv4 I__2579 (
            .O(N__20809),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    Odrv4 I__2578 (
            .O(N__20806),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__2577 (
            .O(N__20801),
            .I(bfn_7_19_0_));
    CascadeMux I__2576 (
            .O(N__20798),
            .I(N__20795));
    InMux I__2575 (
            .O(N__20795),
            .I(N__20791));
    InMux I__2574 (
            .O(N__20794),
            .I(N__20788));
    LocalMux I__2573 (
            .O(N__20791),
            .I(N__20785));
    LocalMux I__2572 (
            .O(N__20788),
            .I(N__20782));
    Odrv12 I__2571 (
            .O(N__20785),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__2570 (
            .O(N__20782),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__2569 (
            .O(N__20777),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__2568 (
            .O(N__20774),
            .I(N__20770));
    CascadeMux I__2567 (
            .O(N__20773),
            .I(N__20767));
    InMux I__2566 (
            .O(N__20770),
            .I(N__20764));
    InMux I__2565 (
            .O(N__20767),
            .I(N__20761));
    LocalMux I__2564 (
            .O(N__20764),
            .I(N__20758));
    LocalMux I__2563 (
            .O(N__20761),
            .I(N__20755));
    Odrv12 I__2562 (
            .O(N__20758),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv4 I__2561 (
            .O(N__20755),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__2560 (
            .O(N__20750),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__2559 (
            .O(N__20747),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__2558 (
            .O(N__20744),
            .I(N__20741));
    InMux I__2557 (
            .O(N__20741),
            .I(N__20736));
    InMux I__2556 (
            .O(N__20740),
            .I(N__20731));
    InMux I__2555 (
            .O(N__20739),
            .I(N__20731));
    LocalMux I__2554 (
            .O(N__20736),
            .I(N__20726));
    LocalMux I__2553 (
            .O(N__20731),
            .I(N__20726));
    Odrv4 I__2552 (
            .O(N__20726),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ));
    InMux I__2551 (
            .O(N__20723),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__2550 (
            .O(N__20720),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__2549 (
            .O(N__20717),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__2548 (
            .O(N__20714),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__2547 (
            .O(N__20711),
            .I(N__20708));
    LocalMux I__2546 (
            .O(N__20708),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10 ));
    CascadeMux I__2545 (
            .O(N__20705),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_ ));
    InMux I__2544 (
            .O(N__20702),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__2543 (
            .O(N__20699),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__2542 (
            .O(N__20696),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__2541 (
            .O(N__20693),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__2540 (
            .O(N__20690),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__2539 (
            .O(N__20687),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__2538 (
            .O(N__20684),
            .I(N__20681));
    LocalMux I__2537 (
            .O(N__20681),
            .I(N__20678));
    Odrv12 I__2536 (
            .O(N__20678),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ));
    CascadeMux I__2535 (
            .O(N__20675),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_ ));
    CascadeMux I__2534 (
            .O(N__20672),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4_cascade_ ));
    InMux I__2533 (
            .O(N__20669),
            .I(N__20666));
    LocalMux I__2532 (
            .O(N__20666),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5 ));
    CascadeMux I__2531 (
            .O(N__20663),
            .I(elapsed_time_ns_1_RNIP1MD11_0_12_cascade_));
    CascadeMux I__2530 (
            .O(N__20660),
            .I(N__20657));
    InMux I__2529 (
            .O(N__20657),
            .I(N__20654));
    LocalMux I__2528 (
            .O(N__20654),
            .I(N__20649));
    InMux I__2527 (
            .O(N__20653),
            .I(N__20644));
    InMux I__2526 (
            .O(N__20652),
            .I(N__20644));
    Odrv4 I__2525 (
            .O(N__20649),
            .I(elapsed_time_ns_1_RNIP1MD11_0_12));
    LocalMux I__2524 (
            .O(N__20644),
            .I(elapsed_time_ns_1_RNIP1MD11_0_12));
    CascadeMux I__2523 (
            .O(N__20639),
            .I(elapsed_time_ns_1_RNINVLD11_0_10_cascade_));
    CascadeMux I__2522 (
            .O(N__20636),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2_cascade_ ));
    InMux I__2521 (
            .O(N__20633),
            .I(N__20629));
    CascadeMux I__2520 (
            .O(N__20632),
            .I(N__20625));
    LocalMux I__2519 (
            .O(N__20629),
            .I(N__20621));
    InMux I__2518 (
            .O(N__20628),
            .I(N__20614));
    InMux I__2517 (
            .O(N__20625),
            .I(N__20614));
    InMux I__2516 (
            .O(N__20624),
            .I(N__20614));
    Odrv4 I__2515 (
            .O(N__20621),
            .I(elapsed_time_ns_1_RNIQ2MD11_0_13));
    LocalMux I__2514 (
            .O(N__20614),
            .I(elapsed_time_ns_1_RNIQ2MD11_0_13));
    CascadeMux I__2513 (
            .O(N__20609),
            .I(elapsed_time_ns_1_RNI51CED1_0_18_cascade_));
    InMux I__2512 (
            .O(N__20606),
            .I(N__20603));
    LocalMux I__2511 (
            .O(N__20603),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18 ));
    CascadeMux I__2510 (
            .O(N__20600),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ));
    CascadeMux I__2509 (
            .O(N__20597),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16_cascade_));
    CascadeMux I__2508 (
            .O(N__20594),
            .I(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9_cascade_ ));
    InMux I__2507 (
            .O(N__20591),
            .I(N__20588));
    LocalMux I__2506 (
            .O(N__20588),
            .I(N__20585));
    Span4Mux_h I__2505 (
            .O(N__20585),
            .I(N__20582));
    Odrv4 I__2504 (
            .O(N__20582),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    CascadeMux I__2503 (
            .O(N__20579),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ));
    InMux I__2502 (
            .O(N__20576),
            .I(N__20573));
    LocalMux I__2501 (
            .O(N__20573),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ));
    InMux I__2500 (
            .O(N__20570),
            .I(N__20567));
    LocalMux I__2499 (
            .O(N__20567),
            .I(N__20564));
    Odrv4 I__2498 (
            .O(N__20564),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__2497 (
            .O(N__20561),
            .I(N__20558));
    LocalMux I__2496 (
            .O(N__20558),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__2495 (
            .O(N__20555),
            .I(N__20549));
    InMux I__2494 (
            .O(N__20554),
            .I(N__20541));
    InMux I__2493 (
            .O(N__20553),
            .I(N__20541));
    CascadeMux I__2492 (
            .O(N__20552),
            .I(N__20538));
    LocalMux I__2491 (
            .O(N__20549),
            .I(N__20535));
    InMux I__2490 (
            .O(N__20548),
            .I(N__20531));
    InMux I__2489 (
            .O(N__20547),
            .I(N__20526));
    InMux I__2488 (
            .O(N__20546),
            .I(N__20526));
    LocalMux I__2487 (
            .O(N__20541),
            .I(N__20522));
    InMux I__2486 (
            .O(N__20538),
            .I(N__20519));
    Span4Mux_s3_h I__2485 (
            .O(N__20535),
            .I(N__20516));
    InMux I__2484 (
            .O(N__20534),
            .I(N__20513));
    LocalMux I__2483 (
            .O(N__20531),
            .I(N__20510));
    LocalMux I__2482 (
            .O(N__20526),
            .I(N__20507));
    InMux I__2481 (
            .O(N__20525),
            .I(N__20504));
    Span4Mux_v I__2480 (
            .O(N__20522),
            .I(N__20499));
    LocalMux I__2479 (
            .O(N__20519),
            .I(N__20499));
    Span4Mux_v I__2478 (
            .O(N__20516),
            .I(N__20494));
    LocalMux I__2477 (
            .O(N__20513),
            .I(N__20494));
    Odrv4 I__2476 (
            .O(N__20510),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv12 I__2475 (
            .O(N__20507),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    LocalMux I__2474 (
            .O(N__20504),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2473 (
            .O(N__20499),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2472 (
            .O(N__20494),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    InMux I__2471 (
            .O(N__20483),
            .I(N__20480));
    LocalMux I__2470 (
            .O(N__20480),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ));
    InMux I__2469 (
            .O(N__20477),
            .I(N__20474));
    LocalMux I__2468 (
            .O(N__20474),
            .I(N__20471));
    Span12Mux_v I__2467 (
            .O(N__20471),
            .I(N__20468));
    Odrv12 I__2466 (
            .O(N__20468),
            .I(il_max_comp2_D1));
    InMux I__2465 (
            .O(N__20465),
            .I(N__20462));
    LocalMux I__2464 (
            .O(N__20462),
            .I(N__20459));
    Glb2LocalMux I__2463 (
            .O(N__20459),
            .I(N__20456));
    GlobalMux I__2462 (
            .O(N__20456),
            .I(clk_12mhz));
    IoInMux I__2461 (
            .O(N__20453),
            .I(N__20450));
    LocalMux I__2460 (
            .O(N__20450),
            .I(N__20447));
    IoSpan4Mux I__2459 (
            .O(N__20447),
            .I(N__20444));
    Span4Mux_s0_v I__2458 (
            .O(N__20444),
            .I(N__20441));
    Odrv4 I__2457 (
            .O(N__20441),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__2456 (
            .O(N__20438),
            .I(N__20435));
    LocalMux I__2455 (
            .O(N__20435),
            .I(N__20432));
    Odrv4 I__2454 (
            .O(N__20432),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    CascadeMux I__2453 (
            .O(N__20429),
            .I(N__20426));
    InMux I__2452 (
            .O(N__20426),
            .I(N__20423));
    LocalMux I__2451 (
            .O(N__20423),
            .I(N__20420));
    Span4Mux_h I__2450 (
            .O(N__20420),
            .I(N__20417));
    Odrv4 I__2449 (
            .O(N__20417),
            .I(\current_shift_inst.PI_CTRL.N_155 ));
    InMux I__2448 (
            .O(N__20414),
            .I(N__20411));
    LocalMux I__2447 (
            .O(N__20411),
            .I(N__20408));
    Odrv4 I__2446 (
            .O(N__20408),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__2445 (
            .O(N__20405),
            .I(N__20402));
    LocalMux I__2444 (
            .O(N__20402),
            .I(N__20399));
    Odrv12 I__2443 (
            .O(N__20399),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__2442 (
            .O(N__20396),
            .I(N__20393));
    LocalMux I__2441 (
            .O(N__20393),
            .I(N__20390));
    Odrv4 I__2440 (
            .O(N__20390),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9 ));
    InMux I__2439 (
            .O(N__20387),
            .I(N__20384));
    LocalMux I__2438 (
            .O(N__20384),
            .I(N__20381));
    Odrv4 I__2437 (
            .O(N__20381),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    InMux I__2436 (
            .O(N__20378),
            .I(N__20373));
    InMux I__2435 (
            .O(N__20377),
            .I(N__20370));
    InMux I__2434 (
            .O(N__20376),
            .I(N__20367));
    LocalMux I__2433 (
            .O(N__20373),
            .I(N__20364));
    LocalMux I__2432 (
            .O(N__20370),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2431 (
            .O(N__20367),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__2430 (
            .O(N__20364),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    CascadeMux I__2429 (
            .O(N__20357),
            .I(N__20354));
    InMux I__2428 (
            .O(N__20354),
            .I(N__20351));
    LocalMux I__2427 (
            .O(N__20351),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2426 (
            .O(N__20348),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2425 (
            .O(N__20345),
            .I(N__20342));
    LocalMux I__2424 (
            .O(N__20342),
            .I(N__20339));
    IoSpan4Mux I__2423 (
            .O(N__20339),
            .I(N__20336));
    Sp12to4 I__2422 (
            .O(N__20336),
            .I(N__20333));
    Span12Mux_s9_v I__2421 (
            .O(N__20333),
            .I(N__20330));
    Span12Mux_h I__2420 (
            .O(N__20330),
            .I(N__20327));
    Odrv12 I__2419 (
            .O(N__20327),
            .I(pwm_output_c));
    CascadeMux I__2418 (
            .O(N__20324),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ));
    CascadeMux I__2417 (
            .O(N__20321),
            .I(N__20316));
    InMux I__2416 (
            .O(N__20320),
            .I(N__20312));
    InMux I__2415 (
            .O(N__20319),
            .I(N__20305));
    InMux I__2414 (
            .O(N__20316),
            .I(N__20305));
    InMux I__2413 (
            .O(N__20315),
            .I(N__20302));
    LocalMux I__2412 (
            .O(N__20312),
            .I(N__20299));
    InMux I__2411 (
            .O(N__20311),
            .I(N__20294));
    InMux I__2410 (
            .O(N__20310),
            .I(N__20294));
    LocalMux I__2409 (
            .O(N__20305),
            .I(N__20291));
    LocalMux I__2408 (
            .O(N__20302),
            .I(N__20287));
    Span4Mux_h I__2407 (
            .O(N__20299),
            .I(N__20284));
    LocalMux I__2406 (
            .O(N__20294),
            .I(N__20279));
    Span4Mux_h I__2405 (
            .O(N__20291),
            .I(N__20279));
    InMux I__2404 (
            .O(N__20290),
            .I(N__20276));
    Odrv12 I__2403 (
            .O(N__20287),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__2402 (
            .O(N__20284),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__2401 (
            .O(N__20279),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    LocalMux I__2400 (
            .O(N__20276),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__2399 (
            .O(N__20267),
            .I(N__20264));
    LocalMux I__2398 (
            .O(N__20264),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    InMux I__2397 (
            .O(N__20261),
            .I(N__20258));
    LocalMux I__2396 (
            .O(N__20258),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    CascadeMux I__2395 (
            .O(N__20255),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ));
    InMux I__2394 (
            .O(N__20252),
            .I(N__20249));
    LocalMux I__2393 (
            .O(N__20249),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    InMux I__2392 (
            .O(N__20246),
            .I(N__20242));
    InMux I__2391 (
            .O(N__20245),
            .I(N__20238));
    LocalMux I__2390 (
            .O(N__20242),
            .I(N__20235));
    InMux I__2389 (
            .O(N__20241),
            .I(N__20232));
    LocalMux I__2388 (
            .O(N__20238),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__2387 (
            .O(N__20235),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2386 (
            .O(N__20232),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    CascadeMux I__2385 (
            .O(N__20225),
            .I(N__20222));
    InMux I__2384 (
            .O(N__20222),
            .I(N__20219));
    LocalMux I__2383 (
            .O(N__20219),
            .I(\pwm_generator_inst.counter_i_1 ));
    InMux I__2382 (
            .O(N__20216),
            .I(N__20213));
    LocalMux I__2381 (
            .O(N__20213),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    InMux I__2380 (
            .O(N__20210),
            .I(N__20205));
    InMux I__2379 (
            .O(N__20209),
            .I(N__20202));
    InMux I__2378 (
            .O(N__20208),
            .I(N__20199));
    LocalMux I__2377 (
            .O(N__20205),
            .I(N__20196));
    LocalMux I__2376 (
            .O(N__20202),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2375 (
            .O(N__20199),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__2374 (
            .O(N__20196),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    CascadeMux I__2373 (
            .O(N__20189),
            .I(N__20186));
    InMux I__2372 (
            .O(N__20186),
            .I(N__20183));
    LocalMux I__2371 (
            .O(N__20183),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__2370 (
            .O(N__20180),
            .I(N__20176));
    InMux I__2369 (
            .O(N__20179),
            .I(N__20172));
    LocalMux I__2368 (
            .O(N__20176),
            .I(N__20169));
    InMux I__2367 (
            .O(N__20175),
            .I(N__20166));
    LocalMux I__2366 (
            .O(N__20172),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__2365 (
            .O(N__20169),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2364 (
            .O(N__20166),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__2363 (
            .O(N__20159),
            .I(N__20156));
    LocalMux I__2362 (
            .O(N__20156),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    CascadeMux I__2361 (
            .O(N__20153),
            .I(N__20150));
    InMux I__2360 (
            .O(N__20150),
            .I(N__20147));
    LocalMux I__2359 (
            .O(N__20147),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__2358 (
            .O(N__20144),
            .I(N__20141));
    LocalMux I__2357 (
            .O(N__20141),
            .I(N__20138));
    Odrv4 I__2356 (
            .O(N__20138),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    InMux I__2355 (
            .O(N__20135),
            .I(N__20131));
    InMux I__2354 (
            .O(N__20134),
            .I(N__20127));
    LocalMux I__2353 (
            .O(N__20131),
            .I(N__20124));
    InMux I__2352 (
            .O(N__20130),
            .I(N__20121));
    LocalMux I__2351 (
            .O(N__20127),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__2350 (
            .O(N__20124),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2349 (
            .O(N__20121),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    CascadeMux I__2348 (
            .O(N__20114),
            .I(N__20111));
    InMux I__2347 (
            .O(N__20111),
            .I(N__20108));
    LocalMux I__2346 (
            .O(N__20108),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__2345 (
            .O(N__20105),
            .I(N__20102));
    LocalMux I__2344 (
            .O(N__20102),
            .I(N__20097));
    InMux I__2343 (
            .O(N__20101),
            .I(N__20094));
    InMux I__2342 (
            .O(N__20100),
            .I(N__20091));
    Odrv4 I__2341 (
            .O(N__20097),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2340 (
            .O(N__20094),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2339 (
            .O(N__20091),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__2338 (
            .O(N__20084),
            .I(N__20081));
    LocalMux I__2337 (
            .O(N__20081),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    CascadeMux I__2336 (
            .O(N__20078),
            .I(N__20075));
    InMux I__2335 (
            .O(N__20075),
            .I(N__20072));
    LocalMux I__2334 (
            .O(N__20072),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__2333 (
            .O(N__20069),
            .I(N__20066));
    LocalMux I__2332 (
            .O(N__20066),
            .I(N__20063));
    Span4Mux_h I__2331 (
            .O(N__20063),
            .I(N__20060));
    Odrv4 I__2330 (
            .O(N__20060),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    InMux I__2329 (
            .O(N__20057),
            .I(N__20054));
    LocalMux I__2328 (
            .O(N__20054),
            .I(N__20049));
    InMux I__2327 (
            .O(N__20053),
            .I(N__20046));
    InMux I__2326 (
            .O(N__20052),
            .I(N__20043));
    Odrv4 I__2325 (
            .O(N__20049),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2324 (
            .O(N__20046),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2323 (
            .O(N__20043),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    CascadeMux I__2322 (
            .O(N__20036),
            .I(N__20033));
    InMux I__2321 (
            .O(N__20033),
            .I(N__20030));
    LocalMux I__2320 (
            .O(N__20030),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__2319 (
            .O(N__20027),
            .I(N__20024));
    LocalMux I__2318 (
            .O(N__20024),
            .I(N__20021));
    Odrv12 I__2317 (
            .O(N__20021),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    InMux I__2316 (
            .O(N__20018),
            .I(N__20014));
    InMux I__2315 (
            .O(N__20017),
            .I(N__20010));
    LocalMux I__2314 (
            .O(N__20014),
            .I(N__20007));
    InMux I__2313 (
            .O(N__20013),
            .I(N__20004));
    LocalMux I__2312 (
            .O(N__20010),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__2311 (
            .O(N__20007),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2310 (
            .O(N__20004),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    CascadeMux I__2309 (
            .O(N__19997),
            .I(N__19994));
    InMux I__2308 (
            .O(N__19994),
            .I(N__19991));
    LocalMux I__2307 (
            .O(N__19991),
            .I(\pwm_generator_inst.counter_i_7 ));
    InMux I__2306 (
            .O(N__19988),
            .I(N__19985));
    LocalMux I__2305 (
            .O(N__19985),
            .I(N__19982));
    Odrv12 I__2304 (
            .O(N__19982),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    InMux I__2303 (
            .O(N__19979),
            .I(N__19974));
    InMux I__2302 (
            .O(N__19978),
            .I(N__19971));
    InMux I__2301 (
            .O(N__19977),
            .I(N__19968));
    LocalMux I__2300 (
            .O(N__19974),
            .I(N__19965));
    LocalMux I__2299 (
            .O(N__19971),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__2298 (
            .O(N__19968),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__2297 (
            .O(N__19965),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    CascadeMux I__2296 (
            .O(N__19958),
            .I(N__19955));
    InMux I__2295 (
            .O(N__19955),
            .I(N__19952));
    LocalMux I__2294 (
            .O(N__19952),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__2293 (
            .O(N__19949),
            .I(N__19946));
    InMux I__2292 (
            .O(N__19946),
            .I(N__19941));
    InMux I__2291 (
            .O(N__19945),
            .I(N__19936));
    InMux I__2290 (
            .O(N__19944),
            .I(N__19936));
    LocalMux I__2289 (
            .O(N__19941),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__2288 (
            .O(N__19936),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__2287 (
            .O(N__19931),
            .I(N__19928));
    LocalMux I__2286 (
            .O(N__19928),
            .I(N__19925));
    Odrv12 I__2285 (
            .O(N__19925),
            .I(il_max_comp2_c));
    InMux I__2284 (
            .O(N__19922),
            .I(N__19919));
    LocalMux I__2283 (
            .O(N__19919),
            .I(N__19916));
    Odrv4 I__2282 (
            .O(N__19916),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__2281 (
            .O(N__19913),
            .I(N__19910));
    LocalMux I__2280 (
            .O(N__19910),
            .I(N__19907));
    Odrv4 I__2279 (
            .O(N__19907),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    InMux I__2278 (
            .O(N__19904),
            .I(N__19901));
    LocalMux I__2277 (
            .O(N__19901),
            .I(N__19898));
    Odrv12 I__2276 (
            .O(N__19898),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    InMux I__2275 (
            .O(N__19895),
            .I(N__19892));
    LocalMux I__2274 (
            .O(N__19892),
            .I(N__19889));
    Odrv4 I__2273 (
            .O(N__19889),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    InMux I__2272 (
            .O(N__19886),
            .I(N__19883));
    LocalMux I__2271 (
            .O(N__19883),
            .I(N__19880));
    Odrv4 I__2270 (
            .O(N__19880),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    CascadeMux I__2269 (
            .O(N__19877),
            .I(N__19874));
    InMux I__2268 (
            .O(N__19874),
            .I(N__19871));
    LocalMux I__2267 (
            .O(N__19871),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    InMux I__2266 (
            .O(N__19868),
            .I(N__19863));
    InMux I__2265 (
            .O(N__19867),
            .I(N__19860));
    InMux I__2264 (
            .O(N__19866),
            .I(N__19857));
    LocalMux I__2263 (
            .O(N__19863),
            .I(N__19854));
    LocalMux I__2262 (
            .O(N__19860),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2261 (
            .O(N__19857),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__2260 (
            .O(N__19854),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2259 (
            .O(N__19847),
            .I(N__19844));
    LocalMux I__2258 (
            .O(N__19844),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__2257 (
            .O(N__19841),
            .I(N__19837));
    InMux I__2256 (
            .O(N__19840),
            .I(N__19834));
    InMux I__2255 (
            .O(N__19837),
            .I(N__19831));
    LocalMux I__2254 (
            .O(N__19834),
            .I(N__19828));
    LocalMux I__2253 (
            .O(N__19831),
            .I(N__19823));
    Span4Mux_v I__2252 (
            .O(N__19828),
            .I(N__19823));
    Odrv4 I__2251 (
            .O(N__19823),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    InMux I__2250 (
            .O(N__19820),
            .I(N__19817));
    LocalMux I__2249 (
            .O(N__19817),
            .I(N__19813));
    InMux I__2248 (
            .O(N__19816),
            .I(N__19809));
    Span4Mux_h I__2247 (
            .O(N__19813),
            .I(N__19806));
    InMux I__2246 (
            .O(N__19812),
            .I(N__19803));
    LocalMux I__2245 (
            .O(N__19809),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    Odrv4 I__2244 (
            .O(N__19806),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    LocalMux I__2243 (
            .O(N__19803),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    CascadeMux I__2242 (
            .O(N__19796),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ));
    InMux I__2241 (
            .O(N__19793),
            .I(N__19790));
    LocalMux I__2240 (
            .O(N__19790),
            .I(N__19786));
    InMux I__2239 (
            .O(N__19789),
            .I(N__19783));
    Span4Mux_v I__2238 (
            .O(N__19786),
            .I(N__19777));
    LocalMux I__2237 (
            .O(N__19783),
            .I(N__19777));
    InMux I__2236 (
            .O(N__19782),
            .I(N__19774));
    Odrv4 I__2235 (
            .O(N__19777),
            .I(pwm_duty_input_9));
    LocalMux I__2234 (
            .O(N__19774),
            .I(pwm_duty_input_9));
    CascadeMux I__2233 (
            .O(N__19769),
            .I(N__19764));
    InMux I__2232 (
            .O(N__19768),
            .I(N__19761));
    InMux I__2231 (
            .O(N__19767),
            .I(N__19758));
    InMux I__2230 (
            .O(N__19764),
            .I(N__19755));
    LocalMux I__2229 (
            .O(N__19761),
            .I(N__19752));
    LocalMux I__2228 (
            .O(N__19758),
            .I(N__19749));
    LocalMux I__2227 (
            .O(N__19755),
            .I(N__19742));
    Span4Mux_v I__2226 (
            .O(N__19752),
            .I(N__19742));
    Span4Mux_v I__2225 (
            .O(N__19749),
            .I(N__19742));
    Odrv4 I__2224 (
            .O(N__19742),
            .I(pwm_duty_input_6));
    InMux I__2223 (
            .O(N__19739),
            .I(N__19734));
    CascadeMux I__2222 (
            .O(N__19738),
            .I(N__19731));
    InMux I__2221 (
            .O(N__19737),
            .I(N__19728));
    LocalMux I__2220 (
            .O(N__19734),
            .I(N__19725));
    InMux I__2219 (
            .O(N__19731),
            .I(N__19722));
    LocalMux I__2218 (
            .O(N__19728),
            .I(N__19719));
    Span4Mux_h I__2217 (
            .O(N__19725),
            .I(N__19716));
    LocalMux I__2216 (
            .O(N__19722),
            .I(N__19711));
    Span4Mux_h I__2215 (
            .O(N__19719),
            .I(N__19711));
    Odrv4 I__2214 (
            .O(N__19716),
            .I(pwm_duty_input_7));
    Odrv4 I__2213 (
            .O(N__19711),
            .I(pwm_duty_input_7));
    InMux I__2212 (
            .O(N__19706),
            .I(N__19702));
    InMux I__2211 (
            .O(N__19705),
            .I(N__19699));
    LocalMux I__2210 (
            .O(N__19702),
            .I(N__19696));
    LocalMux I__2209 (
            .O(N__19699),
            .I(N__19693));
    Span4Mux_h I__2208 (
            .O(N__19696),
            .I(N__19689));
    Span4Mux_v I__2207 (
            .O(N__19693),
            .I(N__19686));
    InMux I__2206 (
            .O(N__19692),
            .I(N__19683));
    Odrv4 I__2205 (
            .O(N__19689),
            .I(pwm_duty_input_8));
    Odrv4 I__2204 (
            .O(N__19686),
            .I(pwm_duty_input_8));
    LocalMux I__2203 (
            .O(N__19683),
            .I(pwm_duty_input_8));
    InMux I__2202 (
            .O(N__19676),
            .I(N__19673));
    LocalMux I__2201 (
            .O(N__19673),
            .I(N__19670));
    Odrv4 I__2200 (
            .O(N__19670),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ));
    InMux I__2199 (
            .O(N__19667),
            .I(N__19664));
    LocalMux I__2198 (
            .O(N__19664),
            .I(N__19661));
    Odrv4 I__2197 (
            .O(N__19661),
            .I(\current_shift_inst.PI_CTRL.N_149 ));
    CascadeMux I__2196 (
            .O(N__19658),
            .I(N__19655));
    InMux I__2195 (
            .O(N__19655),
            .I(N__19651));
    InMux I__2194 (
            .O(N__19654),
            .I(N__19648));
    LocalMux I__2193 (
            .O(N__19651),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__2192 (
            .O(N__19648),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__2191 (
            .O(N__19643),
            .I(N__19637));
    CascadeMux I__2190 (
            .O(N__19642),
            .I(N__19634));
    InMux I__2189 (
            .O(N__19641),
            .I(N__19624));
    InMux I__2188 (
            .O(N__19640),
            .I(N__19624));
    InMux I__2187 (
            .O(N__19637),
            .I(N__19624));
    InMux I__2186 (
            .O(N__19634),
            .I(N__19624));
    InMux I__2185 (
            .O(N__19633),
            .I(N__19621));
    LocalMux I__2184 (
            .O(N__19624),
            .I(N__19618));
    LocalMux I__2183 (
            .O(N__19621),
            .I(N__19615));
    Odrv12 I__2182 (
            .O(N__19618),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    Odrv4 I__2181 (
            .O(N__19615),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    CascadeMux I__2180 (
            .O(N__19610),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__2179 (
            .O(N__19607),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__2178 (
            .O(N__19604),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__2177 (
            .O(N__19601),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__2176 (
            .O(N__19598),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__2175 (
            .O(N__19595),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__2174 (
            .O(N__19592),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__2173 (
            .O(N__19589),
            .I(bfn_4_10_0_));
    InMux I__2172 (
            .O(N__19586),
            .I(N__19568));
    InMux I__2171 (
            .O(N__19585),
            .I(N__19568));
    InMux I__2170 (
            .O(N__19584),
            .I(N__19568));
    InMux I__2169 (
            .O(N__19583),
            .I(N__19568));
    InMux I__2168 (
            .O(N__19582),
            .I(N__19563));
    InMux I__2167 (
            .O(N__19581),
            .I(N__19563));
    InMux I__2166 (
            .O(N__19580),
            .I(N__19554));
    InMux I__2165 (
            .O(N__19579),
            .I(N__19554));
    InMux I__2164 (
            .O(N__19578),
            .I(N__19554));
    InMux I__2163 (
            .O(N__19577),
            .I(N__19554));
    LocalMux I__2162 (
            .O(N__19568),
            .I(N__19547));
    LocalMux I__2161 (
            .O(N__19563),
            .I(N__19547));
    LocalMux I__2160 (
            .O(N__19554),
            .I(N__19547));
    Odrv4 I__2159 (
            .O(N__19547),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__2158 (
            .O(N__19544),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__2157 (
            .O(N__19541),
            .I(N__19537));
    InMux I__2156 (
            .O(N__19540),
            .I(N__19534));
    LocalMux I__2155 (
            .O(N__19537),
            .I(N__19531));
    LocalMux I__2154 (
            .O(N__19534),
            .I(N__19527));
    Span4Mux_v I__2153 (
            .O(N__19531),
            .I(N__19524));
    InMux I__2152 (
            .O(N__19530),
            .I(N__19521));
    Span4Mux_h I__2151 (
            .O(N__19527),
            .I(N__19518));
    Odrv4 I__2150 (
            .O(N__19524),
            .I(pwm_duty_input_4));
    LocalMux I__2149 (
            .O(N__19521),
            .I(pwm_duty_input_4));
    Odrv4 I__2148 (
            .O(N__19518),
            .I(pwm_duty_input_4));
    InMux I__2147 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__2146 (
            .O(N__19508),
            .I(N__19505));
    Odrv4 I__2145 (
            .O(N__19505),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    InMux I__2144 (
            .O(N__19502),
            .I(N__19488));
    InMux I__2143 (
            .O(N__19501),
            .I(N__19488));
    InMux I__2142 (
            .O(N__19500),
            .I(N__19483));
    InMux I__2141 (
            .O(N__19499),
            .I(N__19483));
    InMux I__2140 (
            .O(N__19498),
            .I(N__19480));
    InMux I__2139 (
            .O(N__19497),
            .I(N__19469));
    InMux I__2138 (
            .O(N__19496),
            .I(N__19469));
    InMux I__2137 (
            .O(N__19495),
            .I(N__19469));
    InMux I__2136 (
            .O(N__19494),
            .I(N__19469));
    InMux I__2135 (
            .O(N__19493),
            .I(N__19469));
    LocalMux I__2134 (
            .O(N__19488),
            .I(N__19466));
    LocalMux I__2133 (
            .O(N__19483),
            .I(N__19463));
    LocalMux I__2132 (
            .O(N__19480),
            .I(N__19460));
    LocalMux I__2131 (
            .O(N__19469),
            .I(N__19457));
    Span4Mux_s3_h I__2130 (
            .O(N__19466),
            .I(N__19450));
    Span4Mux_v I__2129 (
            .O(N__19463),
            .I(N__19450));
    Span4Mux_h I__2128 (
            .O(N__19460),
            .I(N__19450));
    Odrv12 I__2127 (
            .O(N__19457),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__2126 (
            .O(N__19450),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__2125 (
            .O(N__19445),
            .I(N__19437));
    CascadeMux I__2124 (
            .O(N__19444),
            .I(N__19434));
    CascadeMux I__2123 (
            .O(N__19443),
            .I(N__19428));
    CascadeMux I__2122 (
            .O(N__19442),
            .I(N__19425));
    CascadeMux I__2121 (
            .O(N__19441),
            .I(N__19422));
    CascadeMux I__2120 (
            .O(N__19440),
            .I(N__19419));
    InMux I__2119 (
            .O(N__19437),
            .I(N__19406));
    InMux I__2118 (
            .O(N__19434),
            .I(N__19406));
    InMux I__2117 (
            .O(N__19433),
            .I(N__19403));
    InMux I__2116 (
            .O(N__19432),
            .I(N__19392));
    InMux I__2115 (
            .O(N__19431),
            .I(N__19392));
    InMux I__2114 (
            .O(N__19428),
            .I(N__19392));
    InMux I__2113 (
            .O(N__19425),
            .I(N__19392));
    InMux I__2112 (
            .O(N__19422),
            .I(N__19392));
    InMux I__2111 (
            .O(N__19419),
            .I(N__19387));
    InMux I__2110 (
            .O(N__19418),
            .I(N__19387));
    InMux I__2109 (
            .O(N__19417),
            .I(N__19382));
    InMux I__2108 (
            .O(N__19416),
            .I(N__19382));
    CascadeMux I__2107 (
            .O(N__19415),
            .I(N__19379));
    CascadeMux I__2106 (
            .O(N__19414),
            .I(N__19376));
    InMux I__2105 (
            .O(N__19413),
            .I(N__19369));
    InMux I__2104 (
            .O(N__19412),
            .I(N__19369));
    InMux I__2103 (
            .O(N__19411),
            .I(N__19369));
    LocalMux I__2102 (
            .O(N__19406),
            .I(N__19366));
    LocalMux I__2101 (
            .O(N__19403),
            .I(N__19346));
    LocalMux I__2100 (
            .O(N__19392),
            .I(N__19346));
    LocalMux I__2099 (
            .O(N__19387),
            .I(N__19341));
    LocalMux I__2098 (
            .O(N__19382),
            .I(N__19341));
    InMux I__2097 (
            .O(N__19379),
            .I(N__19336));
    InMux I__2096 (
            .O(N__19376),
            .I(N__19336));
    LocalMux I__2095 (
            .O(N__19369),
            .I(N__19333));
    Span4Mux_h I__2094 (
            .O(N__19366),
            .I(N__19330));
    InMux I__2093 (
            .O(N__19365),
            .I(N__19313));
    InMux I__2092 (
            .O(N__19364),
            .I(N__19313));
    InMux I__2091 (
            .O(N__19363),
            .I(N__19313));
    InMux I__2090 (
            .O(N__19362),
            .I(N__19313));
    InMux I__2089 (
            .O(N__19361),
            .I(N__19313));
    InMux I__2088 (
            .O(N__19360),
            .I(N__19313));
    InMux I__2087 (
            .O(N__19359),
            .I(N__19313));
    InMux I__2086 (
            .O(N__19358),
            .I(N__19313));
    InMux I__2085 (
            .O(N__19357),
            .I(N__19298));
    InMux I__2084 (
            .O(N__19356),
            .I(N__19298));
    InMux I__2083 (
            .O(N__19355),
            .I(N__19298));
    InMux I__2082 (
            .O(N__19354),
            .I(N__19298));
    InMux I__2081 (
            .O(N__19353),
            .I(N__19298));
    InMux I__2080 (
            .O(N__19352),
            .I(N__19298));
    InMux I__2079 (
            .O(N__19351),
            .I(N__19298));
    Span4Mux_h I__2078 (
            .O(N__19346),
            .I(N__19293));
    Span4Mux_v I__2077 (
            .O(N__19341),
            .I(N__19293));
    LocalMux I__2076 (
            .O(N__19336),
            .I(N__19288));
    Span4Mux_v I__2075 (
            .O(N__19333),
            .I(N__19288));
    Odrv4 I__2074 (
            .O(N__19330),
            .I(N_19_1));
    LocalMux I__2073 (
            .O(N__19313),
            .I(N_19_1));
    LocalMux I__2072 (
            .O(N__19298),
            .I(N_19_1));
    Odrv4 I__2071 (
            .O(N__19293),
            .I(N_19_1));
    Odrv4 I__2070 (
            .O(N__19288),
            .I(N_19_1));
    CascadeMux I__2069 (
            .O(N__19277),
            .I(N__19274));
    InMux I__2068 (
            .O(N__19274),
            .I(N__19271));
    LocalMux I__2067 (
            .O(N__19271),
            .I(N__19268));
    Odrv4 I__2066 (
            .O(N__19268),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__2065 (
            .O(N__19265),
            .I(N__19259));
    InMux I__2064 (
            .O(N__19264),
            .I(N__19259));
    LocalMux I__2063 (
            .O(N__19259),
            .I(N__19250));
    InMux I__2062 (
            .O(N__19258),
            .I(N__19247));
    InMux I__2061 (
            .O(N__19257),
            .I(N__19236));
    InMux I__2060 (
            .O(N__19256),
            .I(N__19236));
    InMux I__2059 (
            .O(N__19255),
            .I(N__19236));
    InMux I__2058 (
            .O(N__19254),
            .I(N__19236));
    InMux I__2057 (
            .O(N__19253),
            .I(N__19236));
    Span4Mux_v I__2056 (
            .O(N__19250),
            .I(N__19227));
    LocalMux I__2055 (
            .O(N__19247),
            .I(N__19227));
    LocalMux I__2054 (
            .O(N__19236),
            .I(N__19227));
    InMux I__2053 (
            .O(N__19235),
            .I(N__19222));
    InMux I__2052 (
            .O(N__19234),
            .I(N__19222));
    Span4Mux_v I__2051 (
            .O(N__19227),
            .I(N__19219));
    LocalMux I__2050 (
            .O(N__19222),
            .I(N__19216));
    Odrv4 I__2049 (
            .O(N__19219),
            .I(\pwm_generator_inst.N_17 ));
    Odrv12 I__2048 (
            .O(N__19216),
            .I(\pwm_generator_inst.N_17 ));
    InMux I__2047 (
            .O(N__19211),
            .I(N__19208));
    LocalMux I__2046 (
            .O(N__19208),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__2045 (
            .O(N__19205),
            .I(N__19202));
    LocalMux I__2044 (
            .O(N__19202),
            .I(N__19199));
    Odrv4 I__2043 (
            .O(N__19199),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    InMux I__2042 (
            .O(N__19196),
            .I(N__19193));
    LocalMux I__2041 (
            .O(N__19193),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    InMux I__2040 (
            .O(N__19190),
            .I(N__19187));
    LocalMux I__2039 (
            .O(N__19187),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    InMux I__2038 (
            .O(N__19184),
            .I(bfn_4_9_0_));
    InMux I__2037 (
            .O(N__19181),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__2036 (
            .O(N__19178),
            .I(N__19175));
    LocalMux I__2035 (
            .O(N__19175),
            .I(N__19171));
    InMux I__2034 (
            .O(N__19174),
            .I(N__19168));
    Span4Mux_h I__2033 (
            .O(N__19171),
            .I(N__19165));
    LocalMux I__2032 (
            .O(N__19168),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    Odrv4 I__2031 (
            .O(N__19165),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    InMux I__2030 (
            .O(N__19160),
            .I(N__19157));
    LocalMux I__2029 (
            .O(N__19157),
            .I(N__19152));
    InMux I__2028 (
            .O(N__19156),
            .I(N__19149));
    InMux I__2027 (
            .O(N__19155),
            .I(N__19146));
    Span4Mux_s3_h I__2026 (
            .O(N__19152),
            .I(N__19141));
    LocalMux I__2025 (
            .O(N__19149),
            .I(N__19141));
    LocalMux I__2024 (
            .O(N__19146),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    Odrv4 I__2023 (
            .O(N__19141),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    InMux I__2022 (
            .O(N__19136),
            .I(N__19133));
    LocalMux I__2021 (
            .O(N__19133),
            .I(N__19129));
    InMux I__2020 (
            .O(N__19132),
            .I(N__19126));
    Odrv4 I__2019 (
            .O(N__19129),
            .I(pwm_duty_input_0));
    LocalMux I__2018 (
            .O(N__19126),
            .I(pwm_duty_input_0));
    InMux I__2017 (
            .O(N__19121),
            .I(N__19118));
    LocalMux I__2016 (
            .O(N__19118),
            .I(N__19114));
    InMux I__2015 (
            .O(N__19117),
            .I(N__19111));
    Odrv4 I__2014 (
            .O(N__19114),
            .I(pwm_duty_input_1));
    LocalMux I__2013 (
            .O(N__19111),
            .I(pwm_duty_input_1));
    InMux I__2012 (
            .O(N__19106),
            .I(N__19103));
    LocalMux I__2011 (
            .O(N__19103),
            .I(N__19099));
    InMux I__2010 (
            .O(N__19102),
            .I(N__19096));
    Odrv4 I__2009 (
            .O(N__19099),
            .I(pwm_duty_input_2));
    LocalMux I__2008 (
            .O(N__19096),
            .I(pwm_duty_input_2));
    InMux I__2007 (
            .O(N__19091),
            .I(N__19088));
    LocalMux I__2006 (
            .O(N__19088),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__2005 (
            .O(N__19085),
            .I(N__19081));
    InMux I__2004 (
            .O(N__19084),
            .I(N__19078));
    LocalMux I__2003 (
            .O(N__19081),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__2002 (
            .O(N__19078),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    InMux I__2001 (
            .O(N__19073),
            .I(N__19067));
    InMux I__2000 (
            .O(N__19072),
            .I(N__19067));
    LocalMux I__1999 (
            .O(N__19067),
            .I(N__19064));
    Span4Mux_h I__1998 (
            .O(N__19064),
            .I(N__19061));
    Odrv4 I__1997 (
            .O(N__19061),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    InMux I__1996 (
            .O(N__19058),
            .I(N__19055));
    LocalMux I__1995 (
            .O(N__19055),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    CascadeMux I__1994 (
            .O(N__19052),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ));
    CascadeMux I__1993 (
            .O(N__19049),
            .I(N__19042));
    CascadeMux I__1992 (
            .O(N__19048),
            .I(N__19039));
    CascadeMux I__1991 (
            .O(N__19047),
            .I(N__19036));
    InMux I__1990 (
            .O(N__19046),
            .I(N__19033));
    CascadeMux I__1989 (
            .O(N__19045),
            .I(N__19030));
    InMux I__1988 (
            .O(N__19042),
            .I(N__19023));
    InMux I__1987 (
            .O(N__19039),
            .I(N__19023));
    InMux I__1986 (
            .O(N__19036),
            .I(N__19019));
    LocalMux I__1985 (
            .O(N__19033),
            .I(N__19015));
    InMux I__1984 (
            .O(N__19030),
            .I(N__19008));
    InMux I__1983 (
            .O(N__19029),
            .I(N__19008));
    InMux I__1982 (
            .O(N__19028),
            .I(N__19008));
    LocalMux I__1981 (
            .O(N__19023),
            .I(N__19003));
    InMux I__1980 (
            .O(N__19022),
            .I(N__19000));
    LocalMux I__1979 (
            .O(N__19019),
            .I(N__18997));
    InMux I__1978 (
            .O(N__19018),
            .I(N__18994));
    Span4Mux_h I__1977 (
            .O(N__19015),
            .I(N__18989));
    LocalMux I__1976 (
            .O(N__19008),
            .I(N__18989));
    InMux I__1975 (
            .O(N__19007),
            .I(N__18984));
    InMux I__1974 (
            .O(N__19006),
            .I(N__18984));
    Span4Mux_s3_h I__1973 (
            .O(N__19003),
            .I(N__18979));
    LocalMux I__1972 (
            .O(N__19000),
            .I(N__18979));
    Odrv12 I__1971 (
            .O(N__18997),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__1970 (
            .O(N__18994),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__1969 (
            .O(N__18989),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__1968 (
            .O(N__18984),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__1967 (
            .O(N__18979),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    InMux I__1966 (
            .O(N__18968),
            .I(N__18965));
    LocalMux I__1965 (
            .O(N__18965),
            .I(N__18962));
    Span4Mux_v I__1964 (
            .O(N__18962),
            .I(N__18959));
    Odrv4 I__1963 (
            .O(N__18959),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    InMux I__1962 (
            .O(N__18956),
            .I(N__18953));
    LocalMux I__1961 (
            .O(N__18953),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ));
    CascadeMux I__1960 (
            .O(N__18950),
            .I(N__18947));
    InMux I__1959 (
            .O(N__18947),
            .I(N__18944));
    LocalMux I__1958 (
            .O(N__18944),
            .I(N__18941));
    Odrv4 I__1957 (
            .O(N__18941),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    CascadeMux I__1956 (
            .O(N__18938),
            .I(N__18935));
    InMux I__1955 (
            .O(N__18935),
            .I(N__18931));
    InMux I__1954 (
            .O(N__18934),
            .I(N__18928));
    LocalMux I__1953 (
            .O(N__18931),
            .I(N__18925));
    LocalMux I__1952 (
            .O(N__18928),
            .I(N__18922));
    Span4Mux_h I__1951 (
            .O(N__18925),
            .I(N__18919));
    Span4Mux_h I__1950 (
            .O(N__18922),
            .I(N__18916));
    Odrv4 I__1949 (
            .O(N__18919),
            .I(\pwm_generator_inst.O_10 ));
    Odrv4 I__1948 (
            .O(N__18916),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__1947 (
            .O(N__18911),
            .I(N__18906));
    InMux I__1946 (
            .O(N__18910),
            .I(N__18903));
    InMux I__1945 (
            .O(N__18909),
            .I(N__18900));
    LocalMux I__1944 (
            .O(N__18906),
            .I(N__18897));
    LocalMux I__1943 (
            .O(N__18903),
            .I(N__18894));
    LocalMux I__1942 (
            .O(N__18900),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    Odrv4 I__1941 (
            .O(N__18897),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    Odrv12 I__1940 (
            .O(N__18894),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    InMux I__1939 (
            .O(N__18887),
            .I(N__18884));
    LocalMux I__1938 (
            .O(N__18884),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    InMux I__1937 (
            .O(N__18881),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    InMux I__1936 (
            .O(N__18878),
            .I(N__18875));
    LocalMux I__1935 (
            .O(N__18875),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    InMux I__1934 (
            .O(N__18872),
            .I(bfn_3_11_0_));
    InMux I__1933 (
            .O(N__18869),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__1932 (
            .O(N__18866),
            .I(N__18861));
    InMux I__1931 (
            .O(N__18865),
            .I(N__18858));
    InMux I__1930 (
            .O(N__18864),
            .I(N__18855));
    LocalMux I__1929 (
            .O(N__18861),
            .I(N__18852));
    LocalMux I__1928 (
            .O(N__18858),
            .I(N__18849));
    LocalMux I__1927 (
            .O(N__18855),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    Odrv4 I__1926 (
            .O(N__18852),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    Odrv4 I__1925 (
            .O(N__18849),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__1924 (
            .O(N__18842),
            .I(N__18839));
    LocalMux I__1923 (
            .O(N__18839),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    InMux I__1922 (
            .O(N__18836),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__1921 (
            .O(N__18833),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__1920 (
            .O(N__18830),
            .I(N__18827));
    LocalMux I__1919 (
            .O(N__18827),
            .I(N__18824));
    Odrv4 I__1918 (
            .O(N__18824),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    InMux I__1917 (
            .O(N__18821),
            .I(N__18818));
    LocalMux I__1916 (
            .O(N__18818),
            .I(N__18814));
    InMux I__1915 (
            .O(N__18817),
            .I(N__18810));
    Span4Mux_h I__1914 (
            .O(N__18814),
            .I(N__18807));
    InMux I__1913 (
            .O(N__18813),
            .I(N__18804));
    LocalMux I__1912 (
            .O(N__18810),
            .I(pwm_duty_input_3));
    Odrv4 I__1911 (
            .O(N__18807),
            .I(pwm_duty_input_3));
    LocalMux I__1910 (
            .O(N__18804),
            .I(pwm_duty_input_3));
    InMux I__1909 (
            .O(N__18797),
            .I(N__18793));
    InMux I__1908 (
            .O(N__18796),
            .I(N__18790));
    LocalMux I__1907 (
            .O(N__18793),
            .I(N__18787));
    LocalMux I__1906 (
            .O(N__18790),
            .I(N__18784));
    Span4Mux_h I__1905 (
            .O(N__18787),
            .I(N__18781));
    Odrv4 I__1904 (
            .O(N__18784),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    Odrv4 I__1903 (
            .O(N__18781),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    CascadeMux I__1902 (
            .O(N__18776),
            .I(N__18773));
    InMux I__1901 (
            .O(N__18773),
            .I(N__18768));
    InMux I__1900 (
            .O(N__18772),
            .I(N__18763));
    InMux I__1899 (
            .O(N__18771),
            .I(N__18763));
    LocalMux I__1898 (
            .O(N__18768),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__1897 (
            .O(N__18763),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    InMux I__1896 (
            .O(N__18758),
            .I(N__18755));
    LocalMux I__1895 (
            .O(N__18755),
            .I(N__18751));
    InMux I__1894 (
            .O(N__18754),
            .I(N__18748));
    Odrv4 I__1893 (
            .O(N__18751),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    LocalMux I__1892 (
            .O(N__18748),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    InMux I__1891 (
            .O(N__18743),
            .I(N__18734));
    InMux I__1890 (
            .O(N__18742),
            .I(N__18734));
    InMux I__1889 (
            .O(N__18741),
            .I(N__18734));
    LocalMux I__1888 (
            .O(N__18734),
            .I(N__18731));
    Odrv4 I__1887 (
            .O(N__18731),
            .I(\current_shift_inst.PI_CTRL.N_154 ));
    InMux I__1886 (
            .O(N__18728),
            .I(N__18725));
    LocalMux I__1885 (
            .O(N__18725),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    InMux I__1884 (
            .O(N__18722),
            .I(N__18719));
    LocalMux I__1883 (
            .O(N__18719),
            .I(N__18716));
    Span4Mux_v I__1882 (
            .O(N__18716),
            .I(N__18713));
    Odrv4 I__1881 (
            .O(N__18713),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1880 (
            .O(N__18710),
            .I(N__18707));
    LocalMux I__1879 (
            .O(N__18707),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    InMux I__1878 (
            .O(N__18704),
            .I(N__18701));
    LocalMux I__1877 (
            .O(N__18701),
            .I(N__18698));
    Span4Mux_v I__1876 (
            .O(N__18698),
            .I(N__18695));
    Odrv4 I__1875 (
            .O(N__18695),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1874 (
            .O(N__18692),
            .I(N__18689));
    LocalMux I__1873 (
            .O(N__18689),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__1872 (
            .O(N__18686),
            .I(N__18683));
    LocalMux I__1871 (
            .O(N__18683),
            .I(N__18680));
    Odrv4 I__1870 (
            .O(N__18680),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    InMux I__1869 (
            .O(N__18677),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    InMux I__1868 (
            .O(N__18674),
            .I(N__18671));
    LocalMux I__1867 (
            .O(N__18671),
            .I(N__18667));
    InMux I__1866 (
            .O(N__18670),
            .I(N__18664));
    Span4Mux_h I__1865 (
            .O(N__18667),
            .I(N__18661));
    LocalMux I__1864 (
            .O(N__18664),
            .I(N__18658));
    Odrv4 I__1863 (
            .O(N__18661),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    Odrv4 I__1862 (
            .O(N__18658),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__1861 (
            .O(N__18653),
            .I(N__18650));
    LocalMux I__1860 (
            .O(N__18650),
            .I(N__18647));
    Odrv4 I__1859 (
            .O(N__18647),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    InMux I__1858 (
            .O(N__18644),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    InMux I__1857 (
            .O(N__18641),
            .I(N__18636));
    InMux I__1856 (
            .O(N__18640),
            .I(N__18633));
    InMux I__1855 (
            .O(N__18639),
            .I(N__18630));
    LocalMux I__1854 (
            .O(N__18636),
            .I(N__18627));
    LocalMux I__1853 (
            .O(N__18633),
            .I(N__18624));
    LocalMux I__1852 (
            .O(N__18630),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    Odrv4 I__1851 (
            .O(N__18627),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    Odrv4 I__1850 (
            .O(N__18624),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    InMux I__1849 (
            .O(N__18617),
            .I(N__18614));
    LocalMux I__1848 (
            .O(N__18614),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    InMux I__1847 (
            .O(N__18611),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    InMux I__1846 (
            .O(N__18608),
            .I(N__18605));
    LocalMux I__1845 (
            .O(N__18605),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    InMux I__1844 (
            .O(N__18602),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__1843 (
            .O(N__18599),
            .I(N__18596));
    LocalMux I__1842 (
            .O(N__18596),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    InMux I__1841 (
            .O(N__18593),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    InMux I__1840 (
            .O(N__18590),
            .I(N__18583));
    InMux I__1839 (
            .O(N__18589),
            .I(N__18583));
    InMux I__1838 (
            .O(N__18588),
            .I(N__18580));
    LocalMux I__1837 (
            .O(N__18583),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__1836 (
            .O(N__18580),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    InMux I__1835 (
            .O(N__18575),
            .I(N__18572));
    LocalMux I__1834 (
            .O(N__18572),
            .I(N__18569));
    Span4Mux_v I__1833 (
            .O(N__18569),
            .I(N__18566));
    Odrv4 I__1832 (
            .O(N__18566),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1831 (
            .O(N__18563),
            .I(N__18560));
    LocalMux I__1830 (
            .O(N__18560),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__1829 (
            .O(N__18557),
            .I(N__18554));
    LocalMux I__1828 (
            .O(N__18554),
            .I(N__18551));
    Span4Mux_v I__1827 (
            .O(N__18551),
            .I(N__18548));
    Odrv4 I__1826 (
            .O(N__18548),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1825 (
            .O(N__18545),
            .I(N__18542));
    LocalMux I__1824 (
            .O(N__18542),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__1823 (
            .O(N__18539),
            .I(N__18536));
    LocalMux I__1822 (
            .O(N__18536),
            .I(N__18533));
    Span4Mux_h I__1821 (
            .O(N__18533),
            .I(N__18530));
    Odrv4 I__1820 (
            .O(N__18530),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1819 (
            .O(N__18527),
            .I(N__18524));
    LocalMux I__1818 (
            .O(N__18524),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    InMux I__1817 (
            .O(N__18521),
            .I(N__18518));
    LocalMux I__1816 (
            .O(N__18518),
            .I(N__18515));
    Span4Mux_h I__1815 (
            .O(N__18515),
            .I(N__18512));
    Odrv4 I__1814 (
            .O(N__18512),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1813 (
            .O(N__18509),
            .I(N__18506));
    LocalMux I__1812 (
            .O(N__18506),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__1811 (
            .O(N__18503),
            .I(N__18500));
    LocalMux I__1810 (
            .O(N__18500),
            .I(N__18497));
    Span4Mux_h I__1809 (
            .O(N__18497),
            .I(N__18494));
    Odrv4 I__1808 (
            .O(N__18494),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1807 (
            .O(N__18491),
            .I(N__18488));
    LocalMux I__1806 (
            .O(N__18488),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__1805 (
            .O(N__18485),
            .I(N__18482));
    LocalMux I__1804 (
            .O(N__18482),
            .I(N__18479));
    Span4Mux_h I__1803 (
            .O(N__18479),
            .I(N__18476));
    Odrv4 I__1802 (
            .O(N__18476),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1801 (
            .O(N__18473),
            .I(N__18470));
    LocalMux I__1800 (
            .O(N__18470),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__1799 (
            .O(N__18467),
            .I(N__18464));
    LocalMux I__1798 (
            .O(N__18464),
            .I(N__18461));
    Span4Mux_h I__1797 (
            .O(N__18461),
            .I(N__18458));
    Odrv4 I__1796 (
            .O(N__18458),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1795 (
            .O(N__18455),
            .I(N__18452));
    LocalMux I__1794 (
            .O(N__18452),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    InMux I__1793 (
            .O(N__18449),
            .I(N__18446));
    LocalMux I__1792 (
            .O(N__18446),
            .I(N__18443));
    Span4Mux_h I__1791 (
            .O(N__18443),
            .I(N__18440));
    Odrv4 I__1790 (
            .O(N__18440),
            .I(\pwm_generator_inst.O_7 ));
    CascadeMux I__1789 (
            .O(N__18437),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    CascadeMux I__1788 (
            .O(N__18434),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__1787 (
            .O(N__18431),
            .I(N__18428));
    LocalMux I__1786 (
            .O(N__18428),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    InMux I__1785 (
            .O(N__18425),
            .I(N__18422));
    LocalMux I__1784 (
            .O(N__18422),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    InMux I__1783 (
            .O(N__18419),
            .I(N__18416));
    LocalMux I__1782 (
            .O(N__18416),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    InMux I__1781 (
            .O(N__18413),
            .I(N__18410));
    LocalMux I__1780 (
            .O(N__18410),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    CascadeMux I__1779 (
            .O(N__18407),
            .I(N__18404));
    InMux I__1778 (
            .O(N__18404),
            .I(N__18401));
    LocalMux I__1777 (
            .O(N__18401),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    InMux I__1776 (
            .O(N__18398),
            .I(N__18395));
    LocalMux I__1775 (
            .O(N__18395),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    CascadeMux I__1774 (
            .O(N__18392),
            .I(N__18389));
    InMux I__1773 (
            .O(N__18389),
            .I(N__18386));
    LocalMux I__1772 (
            .O(N__18386),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__1771 (
            .O(N__18383),
            .I(N__18380));
    LocalMux I__1770 (
            .O(N__18380),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    CascadeMux I__1769 (
            .O(N__18377),
            .I(N__18368));
    CascadeMux I__1768 (
            .O(N__18376),
            .I(N__18365));
    CascadeMux I__1767 (
            .O(N__18375),
            .I(N__18362));
    CascadeMux I__1766 (
            .O(N__18374),
            .I(N__18358));
    CascadeMux I__1765 (
            .O(N__18373),
            .I(N__18355));
    InMux I__1764 (
            .O(N__18372),
            .I(N__18350));
    InMux I__1763 (
            .O(N__18371),
            .I(N__18350));
    InMux I__1762 (
            .O(N__18368),
            .I(N__18345));
    InMux I__1761 (
            .O(N__18365),
            .I(N__18345));
    InMux I__1760 (
            .O(N__18362),
            .I(N__18336));
    InMux I__1759 (
            .O(N__18361),
            .I(N__18336));
    InMux I__1758 (
            .O(N__18358),
            .I(N__18336));
    InMux I__1757 (
            .O(N__18355),
            .I(N__18336));
    LocalMux I__1756 (
            .O(N__18350),
            .I(N__18329));
    LocalMux I__1755 (
            .O(N__18345),
            .I(N__18329));
    LocalMux I__1754 (
            .O(N__18336),
            .I(N__18329));
    Span4Mux_h I__1753 (
            .O(N__18329),
            .I(N__18326));
    Odrv4 I__1752 (
            .O(N__18326),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    InMux I__1751 (
            .O(N__18323),
            .I(N__18320));
    LocalMux I__1750 (
            .O(N__18320),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__1749 (
            .O(N__18317),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__1748 (
            .O(N__18314),
            .I(N__18311));
    LocalMux I__1747 (
            .O(N__18311),
            .I(N__18308));
    Odrv4 I__1746 (
            .O(N__18308),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    InMux I__1745 (
            .O(N__18305),
            .I(N__18302));
    LocalMux I__1744 (
            .O(N__18302),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    InMux I__1743 (
            .O(N__18299),
            .I(bfn_2_12_0_));
    InMux I__1742 (
            .O(N__18296),
            .I(N__18293));
    LocalMux I__1741 (
            .O(N__18293),
            .I(N__18289));
    InMux I__1740 (
            .O(N__18292),
            .I(N__18286));
    Odrv4 I__1739 (
            .O(N__18289),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    LocalMux I__1738 (
            .O(N__18286),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    CascadeMux I__1737 (
            .O(N__18281),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ));
    CascadeMux I__1736 (
            .O(N__18278),
            .I(N__18275));
    InMux I__1735 (
            .O(N__18275),
            .I(N__18272));
    LocalMux I__1734 (
            .O(N__18272),
            .I(N__18269));
    Odrv4 I__1733 (
            .O(N__18269),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    InMux I__1732 (
            .O(N__18266),
            .I(N__18257));
    InMux I__1731 (
            .O(N__18265),
            .I(N__18257));
    InMux I__1730 (
            .O(N__18264),
            .I(N__18257));
    LocalMux I__1729 (
            .O(N__18257),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1728 (
            .O(N__18254),
            .I(N__18251));
    LocalMux I__1727 (
            .O(N__18251),
            .I(N__18248));
    Odrv12 I__1726 (
            .O(N__18248),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    InMux I__1725 (
            .O(N__18245),
            .I(N__18242));
    LocalMux I__1724 (
            .O(N__18242),
            .I(N__18239));
    Span4Mux_v I__1723 (
            .O(N__18239),
            .I(N__18236));
    Odrv4 I__1722 (
            .O(N__18236),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    CascadeMux I__1721 (
            .O(N__18233),
            .I(N__18228));
    InMux I__1720 (
            .O(N__18232),
            .I(N__18225));
    InMux I__1719 (
            .O(N__18231),
            .I(N__18222));
    InMux I__1718 (
            .O(N__18228),
            .I(N__18219));
    LocalMux I__1717 (
            .O(N__18225),
            .I(N__18216));
    LocalMux I__1716 (
            .O(N__18222),
            .I(N__18213));
    LocalMux I__1715 (
            .O(N__18219),
            .I(N__18210));
    Span4Mux_v I__1714 (
            .O(N__18216),
            .I(N__18207));
    Span4Mux_v I__1713 (
            .O(N__18213),
            .I(N__18204));
    Odrv12 I__1712 (
            .O(N__18210),
            .I(pwm_duty_input_5));
    Odrv4 I__1711 (
            .O(N__18207),
            .I(pwm_duty_input_5));
    Odrv4 I__1710 (
            .O(N__18204),
            .I(pwm_duty_input_5));
    InMux I__1709 (
            .O(N__18197),
            .I(N__18194));
    LocalMux I__1708 (
            .O(N__18194),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__1707 (
            .O(N__18191),
            .I(N__18188));
    LocalMux I__1706 (
            .O(N__18188),
            .I(N__18185));
    Span4Mux_h I__1705 (
            .O(N__18185),
            .I(N__18182));
    Span4Mux_v I__1704 (
            .O(N__18182),
            .I(N__18179));
    Odrv4 I__1703 (
            .O(N__18179),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    CascadeMux I__1702 (
            .O(N__18176),
            .I(N__18173));
    InMux I__1701 (
            .O(N__18173),
            .I(N__18170));
    LocalMux I__1700 (
            .O(N__18170),
            .I(N__18167));
    Span4Mux_h I__1699 (
            .O(N__18167),
            .I(N__18164));
    Odrv4 I__1698 (
            .O(N__18164),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    InMux I__1697 (
            .O(N__18161),
            .I(N__18158));
    LocalMux I__1696 (
            .O(N__18158),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    InMux I__1695 (
            .O(N__18155),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__1694 (
            .O(N__18152),
            .I(N__18149));
    LocalMux I__1693 (
            .O(N__18149),
            .I(N__18146));
    Span4Mux_h I__1692 (
            .O(N__18146),
            .I(N__18143));
    Span4Mux_v I__1691 (
            .O(N__18143),
            .I(N__18140));
    Odrv4 I__1690 (
            .O(N__18140),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    CascadeMux I__1689 (
            .O(N__18137),
            .I(N__18134));
    InMux I__1688 (
            .O(N__18134),
            .I(N__18131));
    LocalMux I__1687 (
            .O(N__18131),
            .I(N__18128));
    Span4Mux_h I__1686 (
            .O(N__18128),
            .I(N__18125));
    Odrv4 I__1685 (
            .O(N__18125),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    InMux I__1684 (
            .O(N__18122),
            .I(N__18119));
    LocalMux I__1683 (
            .O(N__18119),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__1682 (
            .O(N__18116),
            .I(bfn_2_11_0_));
    InMux I__1681 (
            .O(N__18113),
            .I(N__18110));
    LocalMux I__1680 (
            .O(N__18110),
            .I(N__18107));
    Span4Mux_h I__1679 (
            .O(N__18107),
            .I(N__18104));
    Span4Mux_v I__1678 (
            .O(N__18104),
            .I(N__18101));
    Odrv4 I__1677 (
            .O(N__18101),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    CascadeMux I__1676 (
            .O(N__18098),
            .I(N__18095));
    InMux I__1675 (
            .O(N__18095),
            .I(N__18092));
    LocalMux I__1674 (
            .O(N__18092),
            .I(N__18089));
    Span4Mux_h I__1673 (
            .O(N__18089),
            .I(N__18086));
    Span4Mux_s0_h I__1672 (
            .O(N__18086),
            .I(N__18083));
    Odrv4 I__1671 (
            .O(N__18083),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    InMux I__1670 (
            .O(N__18080),
            .I(N__18077));
    LocalMux I__1669 (
            .O(N__18077),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__1668 (
            .O(N__18074),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    InMux I__1667 (
            .O(N__18071),
            .I(N__18068));
    LocalMux I__1666 (
            .O(N__18068),
            .I(N__18065));
    Span4Mux_h I__1665 (
            .O(N__18065),
            .I(N__18062));
    Span4Mux_v I__1664 (
            .O(N__18062),
            .I(N__18059));
    Odrv4 I__1663 (
            .O(N__18059),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1662 (
            .O(N__18056),
            .I(N__18053));
    LocalMux I__1661 (
            .O(N__18053),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__1660 (
            .O(N__18050),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    InMux I__1659 (
            .O(N__18047),
            .I(N__18044));
    LocalMux I__1658 (
            .O(N__18044),
            .I(N__18041));
    Span4Mux_h I__1657 (
            .O(N__18041),
            .I(N__18038));
    Span4Mux_v I__1656 (
            .O(N__18038),
            .I(N__18035));
    Odrv4 I__1655 (
            .O(N__18035),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    InMux I__1654 (
            .O(N__18032),
            .I(N__18029));
    LocalMux I__1653 (
            .O(N__18029),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__1652 (
            .O(N__18026),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    InMux I__1651 (
            .O(N__18023),
            .I(N__18020));
    LocalMux I__1650 (
            .O(N__18020),
            .I(N__18017));
    Span4Mux_v I__1649 (
            .O(N__18017),
            .I(N__18014));
    Span4Mux_v I__1648 (
            .O(N__18014),
            .I(N__18011));
    Odrv4 I__1647 (
            .O(N__18011),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1646 (
            .O(N__18008),
            .I(N__18005));
    LocalMux I__1645 (
            .O(N__18005),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__1644 (
            .O(N__18002),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    CascadeMux I__1643 (
            .O(N__17999),
            .I(N__17996));
    InMux I__1642 (
            .O(N__17996),
            .I(N__17993));
    LocalMux I__1641 (
            .O(N__17993),
            .I(N__17990));
    Span12Mux_h I__1640 (
            .O(N__17990),
            .I(N__17987));
    Odrv12 I__1639 (
            .O(N__17987),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    InMux I__1638 (
            .O(N__17984),
            .I(N__17981));
    LocalMux I__1637 (
            .O(N__17981),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__1636 (
            .O(N__17978),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    InMux I__1635 (
            .O(N__17975),
            .I(N__17972));
    LocalMux I__1634 (
            .O(N__17972),
            .I(N__17969));
    Span12Mux_v I__1633 (
            .O(N__17969),
            .I(N__17966));
    Odrv12 I__1632 (
            .O(N__17966),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__1631 (
            .O(N__17963),
            .I(N__17960));
    LocalMux I__1630 (
            .O(N__17960),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__1629 (
            .O(N__17957),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    InMux I__1628 (
            .O(N__17954),
            .I(N__17951));
    LocalMux I__1627 (
            .O(N__17951),
            .I(N__17948));
    Span4Mux_h I__1626 (
            .O(N__17948),
            .I(N__17945));
    Span4Mux_v I__1625 (
            .O(N__17945),
            .I(N__17942));
    Odrv4 I__1624 (
            .O(N__17942),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1623 (
            .O(N__17939),
            .I(N__17936));
    InMux I__1622 (
            .O(N__17936),
            .I(N__17933));
    LocalMux I__1621 (
            .O(N__17933),
            .I(N__17930));
    Span4Mux_h I__1620 (
            .O(N__17930),
            .I(N__17927));
    Odrv4 I__1619 (
            .O(N__17927),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    InMux I__1618 (
            .O(N__17924),
            .I(N__17921));
    LocalMux I__1617 (
            .O(N__17921),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    InMux I__1616 (
            .O(N__17918),
            .I(N__17915));
    LocalMux I__1615 (
            .O(N__17915),
            .I(N__17912));
    Span4Mux_h I__1614 (
            .O(N__17912),
            .I(N__17909));
    Span4Mux_v I__1613 (
            .O(N__17909),
            .I(N__17906));
    Odrv4 I__1612 (
            .O(N__17906),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    CascadeMux I__1611 (
            .O(N__17903),
            .I(N__17900));
    InMux I__1610 (
            .O(N__17900),
            .I(N__17897));
    LocalMux I__1609 (
            .O(N__17897),
            .I(N__17894));
    Span4Mux_h I__1608 (
            .O(N__17894),
            .I(N__17891));
    Odrv4 I__1607 (
            .O(N__17891),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    CascadeMux I__1606 (
            .O(N__17888),
            .I(N__17885));
    InMux I__1605 (
            .O(N__17885),
            .I(N__17882));
    LocalMux I__1604 (
            .O(N__17882),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__1603 (
            .O(N__17879),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1602 (
            .O(N__17876),
            .I(N__17873));
    LocalMux I__1601 (
            .O(N__17873),
            .I(N__17870));
    Span4Mux_h I__1600 (
            .O(N__17870),
            .I(N__17867));
    Span4Mux_v I__1599 (
            .O(N__17867),
            .I(N__17864));
    Odrv4 I__1598 (
            .O(N__17864),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    CascadeMux I__1597 (
            .O(N__17861),
            .I(N__17858));
    InMux I__1596 (
            .O(N__17858),
            .I(N__17855));
    LocalMux I__1595 (
            .O(N__17855),
            .I(N__17852));
    Span4Mux_h I__1594 (
            .O(N__17852),
            .I(N__17849));
    Odrv4 I__1593 (
            .O(N__17849),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    InMux I__1592 (
            .O(N__17846),
            .I(N__17843));
    LocalMux I__1591 (
            .O(N__17843),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__1590 (
            .O(N__17840),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1589 (
            .O(N__17837),
            .I(N__17834));
    LocalMux I__1588 (
            .O(N__17834),
            .I(N__17831));
    Span4Mux_h I__1587 (
            .O(N__17831),
            .I(N__17828));
    Span4Mux_v I__1586 (
            .O(N__17828),
            .I(N__17825));
    Odrv4 I__1585 (
            .O(N__17825),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    CascadeMux I__1584 (
            .O(N__17822),
            .I(N__17819));
    InMux I__1583 (
            .O(N__17819),
            .I(N__17816));
    LocalMux I__1582 (
            .O(N__17816),
            .I(N__17813));
    Span4Mux_v I__1581 (
            .O(N__17813),
            .I(N__17810));
    Odrv4 I__1580 (
            .O(N__17810),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    CascadeMux I__1579 (
            .O(N__17807),
            .I(N__17804));
    InMux I__1578 (
            .O(N__17804),
            .I(N__17801));
    LocalMux I__1577 (
            .O(N__17801),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    InMux I__1576 (
            .O(N__17798),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1575 (
            .O(N__17795),
            .I(N__17792));
    LocalMux I__1574 (
            .O(N__17792),
            .I(N__17789));
    Span4Mux_v I__1573 (
            .O(N__17789),
            .I(N__17786));
    Span4Mux_v I__1572 (
            .O(N__17786),
            .I(N__17783));
    Odrv4 I__1571 (
            .O(N__17783),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    CascadeMux I__1570 (
            .O(N__17780),
            .I(N__17777));
    InMux I__1569 (
            .O(N__17777),
            .I(N__17774));
    LocalMux I__1568 (
            .O(N__17774),
            .I(N__17771));
    Span4Mux_v I__1567 (
            .O(N__17771),
            .I(N__17768));
    Odrv4 I__1566 (
            .O(N__17768),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    InMux I__1565 (
            .O(N__17765),
            .I(N__17762));
    LocalMux I__1564 (
            .O(N__17762),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    InMux I__1563 (
            .O(N__17759),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1562 (
            .O(N__17756),
            .I(N__17753));
    LocalMux I__1561 (
            .O(N__17753),
            .I(N__17750));
    Span12Mux_h I__1560 (
            .O(N__17750),
            .I(N__17747));
    Odrv12 I__1559 (
            .O(N__17747),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    CascadeMux I__1558 (
            .O(N__17744),
            .I(N__17741));
    InMux I__1557 (
            .O(N__17741),
            .I(N__17738));
    LocalMux I__1556 (
            .O(N__17738),
            .I(N__17735));
    Span4Mux_h I__1555 (
            .O(N__17735),
            .I(N__17732));
    Span4Mux_s0_h I__1554 (
            .O(N__17732),
            .I(N__17729));
    Odrv4 I__1553 (
            .O(N__17729),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    InMux I__1552 (
            .O(N__17726),
            .I(N__17723));
    LocalMux I__1551 (
            .O(N__17723),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__1550 (
            .O(N__17720),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__1549 (
            .O(N__17717),
            .I(N__17714));
    LocalMux I__1548 (
            .O(N__17714),
            .I(N__17711));
    Span12Mux_v I__1547 (
            .O(N__17711),
            .I(N__17708));
    Odrv12 I__1546 (
            .O(N__17708),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    CascadeMux I__1545 (
            .O(N__17705),
            .I(N__17702));
    InMux I__1544 (
            .O(N__17702),
            .I(N__17699));
    LocalMux I__1543 (
            .O(N__17699),
            .I(N__17696));
    Span4Mux_h I__1542 (
            .O(N__17696),
            .I(N__17693));
    Odrv4 I__1541 (
            .O(N__17693),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    InMux I__1540 (
            .O(N__17690),
            .I(N__17687));
    LocalMux I__1539 (
            .O(N__17687),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__1538 (
            .O(N__17684),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__1537 (
            .O(N__17681),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    InMux I__1536 (
            .O(N__17678),
            .I(N__17675));
    LocalMux I__1535 (
            .O(N__17675),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    InMux I__1534 (
            .O(N__17672),
            .I(bfn_2_9_0_));
    InMux I__1533 (
            .O(N__17669),
            .I(N__17666));
    LocalMux I__1532 (
            .O(N__17666),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    InMux I__1531 (
            .O(N__17663),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    InMux I__1530 (
            .O(N__17660),
            .I(N__17657));
    LocalMux I__1529 (
            .O(N__17657),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__1528 (
            .O(N__17654),
            .I(N__17648));
    InMux I__1527 (
            .O(N__17653),
            .I(N__17648));
    LocalMux I__1526 (
            .O(N__17648),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    CascadeMux I__1525 (
            .O(N__17645),
            .I(N__17642));
    InMux I__1524 (
            .O(N__17642),
            .I(N__17639));
    LocalMux I__1523 (
            .O(N__17639),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    CascadeMux I__1522 (
            .O(N__17636),
            .I(N__17632));
    InMux I__1521 (
            .O(N__17635),
            .I(N__17629));
    InMux I__1520 (
            .O(N__17632),
            .I(N__17626));
    LocalMux I__1519 (
            .O(N__17629),
            .I(N__17623));
    LocalMux I__1518 (
            .O(N__17626),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    Odrv4 I__1517 (
            .O(N__17623),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    InMux I__1516 (
            .O(N__17618),
            .I(N__17615));
    LocalMux I__1515 (
            .O(N__17615),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    InMux I__1514 (
            .O(N__17612),
            .I(N__17609));
    LocalMux I__1513 (
            .O(N__17609),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    InMux I__1512 (
            .O(N__17606),
            .I(N__17603));
    LocalMux I__1511 (
            .O(N__17603),
            .I(rgb_drv_RNOZ0));
    InMux I__1510 (
            .O(N__17600),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__1509 (
            .O(N__17597),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    InMux I__1508 (
            .O(N__17594),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__1507 (
            .O(N__17591),
            .I(N__17588));
    LocalMux I__1506 (
            .O(N__17588),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    InMux I__1505 (
            .O(N__17585),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    InMux I__1504 (
            .O(N__17582),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__1503 (
            .O(N__17579),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__1502 (
            .O(N__17576),
            .I(N__17573));
    LocalMux I__1501 (
            .O(N__17573),
            .I(N__17570));
    Span4Mux_v I__1500 (
            .O(N__17570),
            .I(N__17567));
    Odrv4 I__1499 (
            .O(N__17567),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    InMux I__1498 (
            .O(N__17564),
            .I(N__17560));
    InMux I__1497 (
            .O(N__17563),
            .I(N__17557));
    LocalMux I__1496 (
            .O(N__17560),
            .I(N__17552));
    LocalMux I__1495 (
            .O(N__17557),
            .I(N__17552));
    Span4Mux_v I__1494 (
            .O(N__17552),
            .I(N__17549));
    Odrv4 I__1493 (
            .O(N__17549),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    InMux I__1492 (
            .O(N__17546),
            .I(N__17543));
    LocalMux I__1491 (
            .O(N__17543),
            .I(N_38_i_i));
    InMux I__1490 (
            .O(N__17540),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    InMux I__1489 (
            .O(N__17537),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    InMux I__1488 (
            .O(N__17534),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    InMux I__1487 (
            .O(N__17531),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    InMux I__1486 (
            .O(N__17528),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    InMux I__1485 (
            .O(N__17525),
            .I(bfn_1_10_0_));
    InMux I__1484 (
            .O(N__17522),
            .I(N__17519));
    LocalMux I__1483 (
            .O(N__17519),
            .I(N__17516));
    Odrv4 I__1482 (
            .O(N__17516),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1481 (
            .O(N__17513),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    CascadeMux I__1480 (
            .O(N__17510),
            .I(N__17507));
    InMux I__1479 (
            .O(N__17507),
            .I(N__17504));
    LocalMux I__1478 (
            .O(N__17504),
            .I(N__17501));
    Odrv4 I__1477 (
            .O(N__17501),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1476 (
            .O(N__17498),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__1475 (
            .O(N__17495),
            .I(N__17492));
    LocalMux I__1474 (
            .O(N__17492),
            .I(N__17489));
    Odrv4 I__1473 (
            .O(N__17489),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1472 (
            .O(N__17486),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    IoInMux I__1471 (
            .O(N__17483),
            .I(N__17480));
    LocalMux I__1470 (
            .O(N__17480),
            .I(N__17477));
    Span4Mux_s3_v I__1469 (
            .O(N__17477),
            .I(N__17474));
    Span4Mux_h I__1468 (
            .O(N__17474),
            .I(N__17471));
    Sp12to4 I__1467 (
            .O(N__17471),
            .I(N__17468));
    Span12Mux_v I__1466 (
            .O(N__17468),
            .I(N__17465));
    Span12Mux_v I__1465 (
            .O(N__17465),
            .I(N__17462));
    Odrv12 I__1464 (
            .O(N__17462),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1463 (
            .O(N__17459),
            .I(N__17456));
    LocalMux I__1462 (
            .O(N__17456),
            .I(N__17453));
    IoSpan4Mux I__1461 (
            .O(N__17453),
            .I(N__17450));
    IoSpan4Mux I__1460 (
            .O(N__17450),
            .I(N__17447));
    Odrv4 I__1459 (
            .O(N__17447),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_6 ),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_14 ),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_22 ),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_18_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_21_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_18_21_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_3_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_10_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_3_10_0_));
    defparam IN_MUX_bfv_3_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_11_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_3_11_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_18_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_7_0_));
    defparam IN_MUX_bfv_18_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_18_8_0_));
    defparam IN_MUX_bfv_18_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_18_9_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_7_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_18_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_13_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_27_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_13_27_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_7 ),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_13_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .carryinitout(bfn_13_14_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_12_12_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__17483),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__17459),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__27833),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_166_i_g ));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__36653),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_434_i_g ));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__23633),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_432_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__40376),
            .CLKHFEN(N__40378),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__40377),
            .RGB2PWM(N__17546),
            .RGB1(rgb_g),
            .CURREN(N__40485),
            .RGB2(rgb_b),
            .RGB1PWM(N__17606),
            .RGB0PWM(N__44337),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21677),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44951),
            .ce(),
            .sr(N__44170));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_8_0 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_8_0  (
            .in0(N__21670),
            .in1(N__20555),
            .in2(N__21200),
            .in3(N__20320),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44950),
            .ce(),
            .sr(N__44183));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_1_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_1_8_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_1_8_5 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_1_8_5  (
            .in0(N__19501),
            .in1(N__17591),
            .in2(N__19414),
            .in3(N__19234),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44950),
            .ce(),
            .sr(N__44183));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_1_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_1_8_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_1_8_7 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_1_8_7  (
            .in0(N__19502),
            .in1(N__17678),
            .in2(N__19415),
            .in3(N__19235),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44950),
            .ce(),
            .sr(N__44183));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__18670),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__17522),
            .in2(_gnd_net_),
            .in3(N__17513),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17510),
            .in3(N__17498),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__17495),
            .in2(_gnd_net_),
            .in3(N__17486),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__17924),
            .in2(_gnd_net_),
            .in3(N__17537),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(N__40547),
            .in2(N__17888),
            .in3(N__17534),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(N__17846),
            .in2(N__40607),
            .in3(N__17531),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(N__40551),
            .in2(N__17807),
            .in3(N__17528),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__17765),
            .in2(_gnd_net_),
            .in3(N__17525),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__17726),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__17690),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__18161),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__18122),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__18080),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__18056),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(N__18032),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__18008),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__17984),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__17963),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__18323),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17540),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_5  (
            .in0(N__18372),
            .in1(N__17563),
            .in2(_gnd_net_),
            .in3(N__19418),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6  (
            .in0(N__17576),
            .in1(N__17564),
            .in2(N__19440),
            .in3(N__18371),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_1_11_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_1_11_7 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_1_11_7  (
            .in0(N__19676),
            .in1(N__18817),
            .in2(N__18233),
            .in3(N__19541),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_12_0 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_12_0  (
            .in0(N__18741),
            .in1(N__18265),
            .in2(N__19642),
            .in3(N__20963),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44942),
            .ce(),
            .sr(N__44217));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_12_2 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_12_2  (
            .in0(N__18742),
            .in1(N__18266),
            .in2(N__19643),
            .in3(N__20948),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44942),
            .ce(),
            .sr(N__44217));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_12_3 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_12_3  (
            .in0(N__18264),
            .in1(N__18743),
            .in2(N__20930),
            .in3(N__19640),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44942),
            .ce(),
            .sr(N__44217));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_12_4 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_12_4  (
            .in0(N__21673),
            .in1(N__20547),
            .in2(N__21095),
            .in3(N__20315),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44942),
            .ce(),
            .sr(N__44217));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_12_5 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_12_5  (
            .in0(N__20546),
            .in1(N__18758),
            .in2(N__21275),
            .in3(N__19641),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44942),
            .ce(),
            .sr(N__44217));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_13_0 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_13_0  (
            .in0(N__21651),
            .in1(N__20554),
            .in2(N__21164),
            .in3(N__20319),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44939),
            .ce(),
            .sr(N__44224));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_13_1 .LUT_INIT=16'b1111001100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_13_1  (
            .in0(N__20553),
            .in1(N__21652),
            .in2(N__20321),
            .in3(N__21053),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44939),
            .ce(),
            .sr(N__44224));
    defparam rgb_drv_RNO_0_LC_1_29_4.C_ON=1'b0;
    defparam rgb_drv_RNO_0_LC_1_29_4.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_0_LC_1_29_4.LUT_INIT=16'b1010101001010101;
    LogicCell40 rgb_drv_RNO_0_LC_1_29_4 (
            .in0(N__44335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26719),
            .lcout(N_38_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_LC_1_30_6.C_ON=1'b0;
    defparam rgb_drv_RNO_LC_1_30_6.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_LC_1_30_6.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_drv_RNO_LC_1_30_6 (
            .in0(N__44336),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26723),
            .lcout(rgb_drv_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_7_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_7_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(N__17635),
            .in2(_gnd_net_),
            .in3(N__18639),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(N__18245),
            .in2(N__19047),
            .in3(N__19046),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__18653),
            .in2(_gnd_net_),
            .in3(N__17600),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__17618),
            .in2(_gnd_net_),
            .in3(N__17597),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_8_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17645),
            .in3(N__17594),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__17612),
            .in2(_gnd_net_),
            .in3(N__17585),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__17660),
            .in2(_gnd_net_),
            .in3(N__17582),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__18254),
            .in2(_gnd_net_),
            .in3(N__17579),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(N__18968),
            .in2(_gnd_net_),
            .in3(N__17681),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_9_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18278),
            .in3(N__17672),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_9_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_9_1  (
            .in0(N__18830),
            .in1(N__17669),
            .in2(N__19049),
            .in3(N__17663),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2  (
            .in0(N__17654),
            .in1(N__18887),
            .in2(N__19045),
            .in3(N__18589),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_3  (
            .in0(N__18590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17653),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_4 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_4  (
            .in0(N__19028),
            .in1(N__18608),
            .in2(N__19841),
            .in3(N__19820),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_5 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_5  (
            .in0(N__18617),
            .in1(N__18641),
            .in2(N__17636),
            .in3(N__19029),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_6  (
            .in0(N__18864),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18292),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_7  (
            .in0(N__19160),
            .in1(N__18599),
            .in2(N__19048),
            .in3(N__19174),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__17954),
            .in2(N__17939),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__17918),
            .in2(N__17903),
            .in3(N__17879),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__17876),
            .in2(N__17861),
            .in3(N__17840),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__17837),
            .in2(N__17822),
            .in3(N__17798),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__17795),
            .in2(N__17780),
            .in3(N__17759),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(N__17756),
            .in2(N__17744),
            .in3(N__17720),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(N__17717),
            .in2(N__17705),
            .in3(N__17684),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(N__18191),
            .in2(N__18176),
            .in3(N__18155),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__18152),
            .in2(N__18137),
            .in3(N__18116),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__18113),
            .in2(N__18098),
            .in3(N__18074),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__18071),
            .in2(N__18373),
            .in3(N__18050),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__18047),
            .in2(N__18376),
            .in3(N__18026),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__18023),
            .in2(N__18374),
            .in3(N__18002),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__18361),
            .in2(N__17999),
            .in3(N__17978),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__17975),
            .in2(N__18375),
            .in3(N__17957),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__18383),
            .in2(N__18377),
            .in3(N__18317),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_12_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_12_0  (
            .in0(N__18314),
            .in1(N__18305),
            .in2(_gnd_net_),
            .in3(N__18299),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_12_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_12_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_12_1  (
            .in0(N__18296),
            .in1(N__18865),
            .in2(N__18281),
            .in3(N__18842),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_12_3 .LUT_INIT=16'b0011001100000010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_12_3  (
            .in0(N__18754),
            .in1(N__21274),
            .in2(N__20552),
            .in3(N__19633),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_4 .LUT_INIT=16'b1011011110000100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_4  (
            .in0(N__18878),
            .in1(N__19007),
            .in2(N__18776),
            .in3(N__18796),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_12_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_12_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_12_6  (
            .in0(N__18686),
            .in1(N__18911),
            .in2(N__18938),
            .in3(N__19006),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_13_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_13_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__19739),
            .in2(_gnd_net_),
            .in3(N__18232),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_7_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_7_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_7_0 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_3_7_0  (
            .in0(N__19499),
            .in1(N__18197),
            .in2(N__19444),
            .in3(N__19264),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44949),
            .ce(),
            .sr(N__44162));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_3_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_3_7_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_3_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_3_7_2  (
            .in0(_gnd_net_),
            .in1(N__20210),
            .in2(_gnd_net_),
            .in3(N__19868),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_3_7_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_3_7_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_3_7_3 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_3_7_3  (
            .in0(N__20135),
            .in1(N__20180),
            .in2(N__18437),
            .in3(N__20246),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_3_7_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_3_7_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_3_7_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_3_7_4  (
            .in0(N__20057),
            .in1(N__20105),
            .in2(N__18434),
            .in3(N__19511),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_7_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_7_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_7_6 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_3_7_6  (
            .in0(N__19500),
            .in1(N__18431),
            .in2(N__19445),
            .in3(N__19265),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44949),
            .ce(),
            .sr(N__44162));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_8_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_8_0 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_3_8_0  (
            .in0(N__19257),
            .in1(N__19497),
            .in2(N__19443),
            .in3(N__18425),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44947),
            .ce(),
            .sr(N__44171));
    defparam \pwm_generator_inst.threshold_6_LC_3_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_3_8_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_3_8_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_3_8_1  (
            .in0(_gnd_net_),
            .in1(N__18419),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44947),
            .ce(),
            .sr(N__44171));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_8_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_8_2 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_3_8_2  (
            .in0(N__19255),
            .in1(N__19496),
            .in2(N__19442),
            .in3(N__18413),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44947),
            .ce(),
            .sr(N__44171));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_8_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_8_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_8_3 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_3_8_3  (
            .in0(N__19494),
            .in1(N__19432),
            .in2(N__18407),
            .in3(N__19256),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44947),
            .ce(),
            .sr(N__44171));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_8_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_8_4 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_3_8_4  (
            .in0(N__19254),
            .in1(N__19495),
            .in2(N__19441),
            .in3(N__18398),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44947),
            .ce(),
            .sr(N__44171));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_8_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_8_5 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_3_8_5  (
            .in0(N__19493),
            .in1(N__19431),
            .in2(N__18392),
            .in3(N__19253),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44947),
            .ce(),
            .sr(N__44171));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(N__18563),
            .in2(_gnd_net_),
            .in3(N__18575),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1  (
            .in0(_gnd_net_),
            .in1(N__18545),
            .in2(_gnd_net_),
            .in3(N__18557),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(N__18527),
            .in2(_gnd_net_),
            .in3(N__18539),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3  (
            .in0(_gnd_net_),
            .in1(N__18509),
            .in2(_gnd_net_),
            .in3(N__18521),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4  (
            .in0(_gnd_net_),
            .in1(N__18491),
            .in2(_gnd_net_),
            .in3(N__18503),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5  (
            .in0(_gnd_net_),
            .in1(N__18473),
            .in2(_gnd_net_),
            .in3(N__18485),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(N__18455),
            .in2(_gnd_net_),
            .in3(N__18467),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7  (
            .in0(_gnd_net_),
            .in1(N__18728),
            .in2(_gnd_net_),
            .in3(N__18449),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(N__18710),
            .in2(_gnd_net_),
            .in3(N__18722),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_3_10_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1  (
            .in0(_gnd_net_),
            .in1(N__18692),
            .in2(_gnd_net_),
            .in3(N__18704),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(N__18910),
            .in2(_gnd_net_),
            .in3(N__18677),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3  (
            .in0(N__19022),
            .in1(N__18674),
            .in2(_gnd_net_),
            .in3(N__18644),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4  (
            .in0(_gnd_net_),
            .in1(N__18640),
            .in2(_gnd_net_),
            .in3(N__18611),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5  (
            .in0(_gnd_net_),
            .in1(N__19812),
            .in2(_gnd_net_),
            .in3(N__18602),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6  (
            .in0(_gnd_net_),
            .in1(N__19156),
            .in2(_gnd_net_),
            .in3(N__18593),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7  (
            .in0(_gnd_net_),
            .in1(N__18588),
            .in2(_gnd_net_),
            .in3(N__18881),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0  (
            .in0(_gnd_net_),
            .in1(N__18771),
            .in2(_gnd_net_),
            .in3(N__18872),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_3_11_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1  (
            .in0(_gnd_net_),
            .in1(N__19084),
            .in2(_gnd_net_),
            .in3(N__18869),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__18866),
            .in2(_gnd_net_),
            .in3(N__18836),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18833),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_11_6 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_3_11_6  (
            .in0(N__19091),
            .in1(N__18821),
            .in2(N__18950),
            .in3(N__19530),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_3_11_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_3_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_3_11_7  (
            .in0(N__18772),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18797),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_3_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_3_12_1 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_3_12_1  (
            .in0(N__19944),
            .in1(N__21671),
            .in2(_gnd_net_),
            .in3(N__21239),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_12_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_12_2  (
            .in0(N__21672),
            .in1(N__19945),
            .in2(_gnd_net_),
            .in3(N__20534),
            .lcout(\current_shift_inst.PI_CTRL.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_12_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_12_3  (
            .in0(N__19155),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19178),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_3_12_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_3_12_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_3_12_4  (
            .in0(N__19136),
            .in1(N__19121),
            .in2(_gnd_net_),
            .in3(N__19106),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_3_12_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_3_12_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_3_12_5  (
            .in0(_gnd_net_),
            .in1(N__19072),
            .in2(_gnd_net_),
            .in3(N__19085),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_3_12_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_3_12_6 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_3_12_6  (
            .in0(N__19073),
            .in1(N__19058),
            .in2(N__19052),
            .in3(N__19018),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_13_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_13_3 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_13_3  (
            .in0(N__19705),
            .in1(N__19789),
            .in2(N__19769),
            .in3(N__18956),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_3_14_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_3_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_3_14_1  (
            .in0(N__18909),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18934),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_14_LC_3_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_14_LC_3_14_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_14_LC_3_14_4 .LUT_INIT=16'b0000000011111011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_14_LC_3_14_4  (
            .in0(N__24749),
            .in1(N__21593),
            .in2(N__21938),
            .in3(N__26032),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44927),
            .ce(N__25641),
            .sr(N__44218));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_19_LC_3_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_19_LC_3_14_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_19_LC_3_14_5 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_19_LC_3_14_5  (
            .in0(N__26030),
            .in1(N__24480),
            .in2(_gnd_net_),
            .in3(N__24751),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44927),
            .ce(N__25641),
            .sr(N__44218));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_18_LC_3_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_18_LC_3_14_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_18_LC_3_14_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_18_LC_3_14_6  (
            .in0(N__24748),
            .in1(N__26031),
            .in2(_gnd_net_),
            .in3(N__23381),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44927),
            .ce(N__25641),
            .sr(N__44218));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_17_LC_3_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_17_LC_3_14_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_17_LC_3_14_7 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_17_LC_3_14_7  (
            .in0(N__26029),
            .in1(N__23420),
            .in2(_gnd_net_),
            .in3(N__24750),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44927),
            .ce(N__25641),
            .sr(N__44218));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_4_7_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_4_7_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_4_7_6  (
            .in0(N__20378),
            .in1(N__19979),
            .in2(_gnd_net_),
            .in3(N__20018),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_0_LC_4_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_4_8_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_4_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19211),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44945),
            .ce(),
            .sr(N__44163));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_8_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_8_1 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_4_8_1  (
            .in0(N__19498),
            .in1(N__19433),
            .in2(N__19277),
            .in3(N__19258),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44945),
            .ce(),
            .sr(N__44163));
    defparam \pwm_generator_inst.threshold_4_LC_4_8_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_4_8_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_4_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19205),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44945),
            .ce(),
            .sr(N__44163));
    defparam \pwm_generator_inst.threshold_5_LC_4_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_4_8_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_4_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19196),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44945),
            .ce(),
            .sr(N__44163));
    defparam \pwm_generator_inst.threshold_2_LC_4_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_4_8_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_4_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_4_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19190),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44945),
            .ce(),
            .sr(N__44163));
    defparam \pwm_generator_inst.counter_0_LC_4_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_4_9_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_4_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_4_9_0  (
            .in0(N__19577),
            .in1(N__19867),
            .in2(_gnd_net_),
            .in3(N__19184),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__44943),
            .ce(),
            .sr(N__44172));
    defparam \pwm_generator_inst.counter_1_LC_4_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_4_9_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_4_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_4_9_1  (
            .in0(N__19583),
            .in1(N__20245),
            .in2(_gnd_net_),
            .in3(N__19181),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__44943),
            .ce(),
            .sr(N__44172));
    defparam \pwm_generator_inst.counter_2_LC_4_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_4_9_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_4_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_4_9_2  (
            .in0(N__19578),
            .in1(N__20209),
            .in2(_gnd_net_),
            .in3(N__19607),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__44943),
            .ce(),
            .sr(N__44172));
    defparam \pwm_generator_inst.counter_3_LC_4_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_4_9_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_4_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_4_9_3  (
            .in0(N__19584),
            .in1(N__20179),
            .in2(_gnd_net_),
            .in3(N__19604),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__44943),
            .ce(),
            .sr(N__44172));
    defparam \pwm_generator_inst.counter_4_LC_4_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_4_9_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_4_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_4_9_4  (
            .in0(N__19579),
            .in1(N__20134),
            .in2(_gnd_net_),
            .in3(N__19601),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__44943),
            .ce(),
            .sr(N__44172));
    defparam \pwm_generator_inst.counter_5_LC_4_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_4_9_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_4_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_4_9_5  (
            .in0(N__19585),
            .in1(N__20101),
            .in2(_gnd_net_),
            .in3(N__19598),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__44943),
            .ce(),
            .sr(N__44172));
    defparam \pwm_generator_inst.counter_6_LC_4_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_4_9_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_4_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_4_9_6  (
            .in0(N__19580),
            .in1(N__20053),
            .in2(_gnd_net_),
            .in3(N__19595),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__44943),
            .ce(),
            .sr(N__44172));
    defparam \pwm_generator_inst.counter_7_LC_4_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_4_9_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_4_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_4_9_7  (
            .in0(N__19586),
            .in1(N__20017),
            .in2(_gnd_net_),
            .in3(N__19592),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__44943),
            .ce(),
            .sr(N__44172));
    defparam \pwm_generator_inst.counter_8_LC_4_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_4_10_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_4_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_4_10_0  (
            .in0(N__19582),
            .in1(N__19978),
            .in2(_gnd_net_),
            .in3(N__19589),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__44940),
            .ce(),
            .sr(N__44178));
    defparam \pwm_generator_inst.counter_9_LC_4_10_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_4_10_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_4_10_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_4_10_1  (
            .in0(N__20377),
            .in1(N__19581),
            .in2(_gnd_net_),
            .in3(N__19544),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44940),
            .ce(),
            .sr(N__44178));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_4_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_4_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_4_10_4 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_4_10_4  (
            .in0(N__19667),
            .in1(N__21234),
            .in2(N__19658),
            .in3(N__20310),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44940),
            .ce(),
            .sr(N__44178));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_4_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_4_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_4_10_6 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_4_10_6  (
            .in0(N__20548),
            .in1(N__21663),
            .in2(N__21128),
            .in3(N__20311),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44940),
            .ce(),
            .sr(N__44178));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_4_11_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_4_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_4_11_0  (
            .in0(N__19816),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19840),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_4_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_4_11_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_4_11_4  (
            .in0(N__21192),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21091),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_11_5  (
            .in0(N__21126),
            .in1(N__21157),
            .in2(N__19796),
            .in3(N__21048),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_11_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_11_6  (
            .in0(N__19793),
            .in1(N__19768),
            .in2(N__19738),
            .in3(N__19706),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_4_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_4_12_0 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_4_12_0  (
            .in0(N__21238),
            .in1(N__21662),
            .in2(N__19949),
            .in3(N__20525),
            .lcout(\current_shift_inst.PI_CTRL.N_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_4_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_4_12_7 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_4_12_7  (
            .in0(N__21661),
            .in1(N__19654),
            .in2(N__20429),
            .in3(N__20290),
            .lcout(\current_shift_inst.PI_CTRL.N_153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_4_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_4_13_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_4_13_0  (
            .in0(N__21193),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21049),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_4_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_4_13_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_4_13_1  (
            .in0(N__21127),
            .in1(N__21084),
            .in2(N__19610),
            .in3(N__21150),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_4_24_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_24_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_24_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_6_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_6_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_5_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19931),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44948),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_7_LC_5_7_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_5_7_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_5_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19922),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44946),
            .ce(),
            .sr(N__44151));
    defparam \pwm_generator_inst.threshold_3_LC_5_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_5_8_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_5_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19913),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44944),
            .ce(),
            .sr(N__44158));
    defparam \pwm_generator_inst.threshold_8_LC_5_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_5_8_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_5_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19904),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44944),
            .ce(),
            .sr(N__44158));
    defparam \pwm_generator_inst.threshold_9_LC_5_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_5_8_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_5_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19895),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44944),
            .ce(),
            .sr(N__44158));
    defparam \pwm_generator_inst.threshold_1_LC_5_8_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_5_8_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_5_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_5_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19886),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44944),
            .ce(),
            .sr(N__44158));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(N__19847),
            .in2(N__19877),
            .in3(N__19866),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__20252),
            .in2(N__20225),
            .in3(N__20241),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__20216),
            .in2(N__20189),
            .in3(N__20208),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_9_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_9_3  (
            .in0(N__20175),
            .in1(N__20159),
            .in2(N__20153),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__20144),
            .in2(N__20114),
            .in3(N__20130),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_9_5  (
            .in0(N__20100),
            .in1(N__20084),
            .in2(N__20078),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(N__20069),
            .in2(N__20036),
            .in3(N__20052),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__20027),
            .in2(N__19997),
            .in3(N__20013),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__19988),
            .in2(N__19958),
            .in3(N__19977),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__20387),
            .in2(N__20357),
            .in3(N__20376),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_5_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_5_10_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_5_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20348),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44936),
            .ce(),
            .sr(N__44173));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_5_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_5_11_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_5_11_7  (
            .in0(N__20261),
            .in1(N__20438),
            .in2(N__21416),
            .in3(N__21008),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_15_LC_5_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_15_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_15_LC_5_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_15_LC_5_12_0  (
            .in0(N__21482),
            .in1(N__21365),
            .in2(N__21344),
            .in3(N__20396),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_12_1  (
            .in0(N__20267),
            .in1(N__20591),
            .in2(N__20324),
            .in3(N__20570),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_5_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_5_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_5_12_4  (
            .in0(N__21704),
            .in1(N__21461),
            .in2(N__21308),
            .in3(N__21322),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_5_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_5_12_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_5_12_5  (
            .in0(N__21323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21304),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_5_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_5_12_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_5_12_6  (
            .in0(N__20483),
            .in1(N__21545),
            .in2(N__21566),
            .in3(N__21437),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_5_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_5_12_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_5_12_7  (
            .in0(N__20414),
            .in1(N__20405),
            .in2(N__20255),
            .in3(N__20561),
            .lcout(\current_shift_inst.PI_CTRL.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_5_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_5_13_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__21700),
            .in2(_gnd_net_),
            .in3(N__21460),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_19_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_19_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_5_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20477),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44891),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_7.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_7.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20465),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_7_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_7_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__21409),
            .in2(_gnd_net_),
            .in3(N__21019),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_7_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_7_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_7_11_3  (
            .in0(N__21020),
            .in1(N__21358),
            .in2(N__21731),
            .in3(N__21337),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_7_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_7_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__21219),
            .in2(_gnd_net_),
            .in3(N__21255),
            .lcout(\current_shift_inst.PI_CTRL.N_155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_7_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_7_12_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_7_12_0  (
            .in0(N__21287),
            .in1(N__21478),
            .in2(N__21497),
            .in3(N__21578),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_7_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_7_12_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_7_12_2  (
            .in0(N__21527),
            .in1(N__21395),
            .in2(N__21515),
            .in3(N__21382),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPN72_22_LC_7_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPN72_22_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPN72_22_LC_7_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPN72_22_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__21493),
            .in2(_gnd_net_),
            .in3(N__21541),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_7_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_7_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_7_12_4  (
            .in0(N__21286),
            .in1(N__21577),
            .in2(N__21383),
            .in3(N__21394),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_7_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_7_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_7_12_5  (
            .in0(N__21511),
            .in1(N__21526),
            .in2(N__21727),
            .in3(N__21559),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_7_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_7_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_7_12_6  (
            .in0(N__21430),
            .in1(N__21004),
            .in2(N__20579),
            .in3(N__20576),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_9_LC_7_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_9_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_9_LC_7_13_0 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_9_LC_7_13_0  (
            .in0(N__24438),
            .in1(N__25996),
            .in2(N__24752),
            .in3(N__21869),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44911),
            .ce(N__25649),
            .sr(N__44179));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_16_LC_7_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_16_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_16_LC_7_13_1 .LUT_INIT=16'b0000111000001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_16_LC_7_13_1  (
            .in0(N__24737),
            .in1(N__23340),
            .in2(N__26034),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44911),
            .ce(N__25649),
            .sr(N__44179));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_10_LC_7_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_10_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_10_LC_7_13_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_10_LC_7_13_2  (
            .in0(N__24741),
            .in1(N__21856),
            .in2(N__21833),
            .in3(N__25997),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44911),
            .ce(N__25649),
            .sr(N__44179));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_11_LC_7_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_11_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_11_LC_7_13_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_11_LC_7_13_3  (
            .in0(N__26003),
            .in1(N__24743),
            .in2(N__21831),
            .in3(N__21782),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44911),
            .ce(N__25649),
            .sr(N__44179));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_12_LC_7_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_12_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_12_LC_7_13_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_12_LC_7_13_4  (
            .in0(N__21830),
            .in1(N__24738),
            .in2(N__20660),
            .in3(N__25998),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44911),
            .ce(N__25649),
            .sr(N__44179));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_13_LC_7_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_13_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_13_LC_7_13_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_13_LC_7_13_5  (
            .in0(N__26004),
            .in1(N__24744),
            .in2(N__21832),
            .in3(N__20633),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44911),
            .ce(N__25649),
            .sr(N__44179));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_15_LC_7_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_15_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_15_LC_7_13_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_15_LC_7_13_6  (
            .in0(N__24742),
            .in1(N__25999),
            .in2(N__24893),
            .in3(N__24408),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44911),
            .ce(N__25649),
            .sr(N__44179));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_7_LC_7_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_7_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_7_LC_7_13_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_7_LC_7_13_7  (
            .in0(N__25523),
            .in1(_gnd_net_),
            .in2(N__26033),
            .in3(N__25805),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44911),
            .ce(N__25649),
            .sr(N__44179));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_7_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_7_14_0 .LUT_INIT=16'b1111111011001110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_7_14_0  (
            .in0(N__21896),
            .in1(N__31638),
            .in2(N__31864),
            .in3(N__22070),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_7_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_7_14_1 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_7_14_1  (
            .in0(N__21929),
            .in1(N__22040),
            .in2(N__31649),
            .in3(N__31847),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_7_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_7_14_2 .LUT_INIT=16'b1110111111101100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_7_14_2  (
            .in0(N__22100),
            .in1(N__31637),
            .in2(N__31863),
            .in3(N__23336),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_7_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_7_14_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20600),
            .in3(N__25463),
            .lcout(elapsed_time_ns_1_RNI3VBED1_0_16),
            .ltout(elapsed_time_ns_1_RNI3VBED1_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_9_LC_7_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_9_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_9_LC_7_14_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_9_LC_7_14_4  (
            .in0(N__24464),
            .in1(N__23412),
            .in2(N__20597),
            .in3(N__23376),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_10_LC_7_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_10_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_10_LC_7_14_5 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_i_a2_10_LC_7_14_5  (
            .in0(N__21930),
            .in1(_gnd_net_),
            .in2(N__20594),
            .in3(N__24887),
            .lcout(\phase_controller_inst1.stoper_hc.N_315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_7_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_7_15_0 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_7_15_0  (
            .in0(N__26339),
            .in1(N__31817),
            .in2(N__20774),
            .in3(N__20628),
            .lcout(elapsed_time_ns_1_RNIQ2MD11_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_7_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_7_15_1 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_7_15_1  (
            .in0(N__31818),
            .in1(N__26340),
            .in2(N__20798),
            .in3(N__20653),
            .lcout(elapsed_time_ns_1_RNIP1MD11_0_12),
            .ltout(elapsed_time_ns_1_RNIP1MD11_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_12_LC_7_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_12_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_12_LC_7_15_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_12_LC_7_15_2  (
            .in0(N__24739),
            .in1(N__26038),
            .in2(N__20663),
            .in3(N__21824),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44903),
            .ce(N__31528),
            .sr(N__44188));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_7_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_7_15_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_7_15_3  (
            .in0(N__31819),
            .in1(N__26341),
            .in2(N__20825),
            .in3(N__21777),
            .lcout(elapsed_time_ns_1_RNIO0MD11_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_7_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_7_15_4 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_7_15_4  (
            .in0(N__26338),
            .in1(N__31816),
            .in2(N__20846),
            .in3(N__21849),
            .lcout(elapsed_time_ns_1_RNINVLD11_0_10),
            .ltout(elapsed_time_ns_1_RNINVLD11_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2_2_LC_7_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2_2_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2_2_LC_7_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_i_a2_2_2_LC_7_15_5  (
            .in0(N__20624),
            .in1(N__20652),
            .in2(N__20639),
            .in3(N__21776),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a0_6_LC_7_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a0_6_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a0_6_LC_7_15_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a0_6_LC_7_15_6  (
            .in0(N__21888),
            .in1(_gnd_net_),
            .in2(N__20636),
            .in3(N__24883),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_a5_1_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_13_LC_7_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_13_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_13_LC_7_15_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_13_LC_7_15_7  (
            .in0(N__21823),
            .in1(N__24740),
            .in2(N__20632),
            .in3(N__26039),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44903),
            .ce(N__31528),
            .sr(N__44188));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_7_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_7_16_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__20606),
            .in2(_gnd_net_),
            .in3(N__25449),
            .lcout(elapsed_time_ns_1_RNI51CED1_0_18),
            .ltout(elapsed_time_ns_1_RNI51CED1_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_7_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_7_16_1 .LUT_INIT=16'b1111111011011100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_7_16_1  (
            .in0(N__31777),
            .in1(N__31621),
            .in2(N__20609),
            .in3(N__22121),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_7_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_7_16_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_7_16_2  (
            .in0(N__23786),
            .in1(N__22069),
            .in2(N__22004),
            .in3(N__21956),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_7_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_7_16_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_7_16_3  (
            .in0(N__31775),
            .in1(N__21758),
            .in2(N__20900),
            .in3(N__26331),
            .lcout(elapsed_time_ns_1_RNIR4ND11_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_7_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_7_16_4 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_7_16_4  (
            .in0(N__26332),
            .in1(N__31778),
            .in2(N__20744),
            .in3(N__24882),
            .lcout(elapsed_time_ns_1_RNIS4MD11_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_7_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_7_16_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_7_16_5  (
            .in0(N__25450),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20684),
            .lcout(elapsed_time_ns_1_RNIL13KD1_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_7_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_7_16_6 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_7_16_6  (
            .in0(N__21746),
            .in1(N__20876),
            .in2(N__26373),
            .in3(N__31776),
            .lcout(elapsed_time_ns_1_RNIS5ND11_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_7_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_7_16_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_7_16_7  (
            .in0(N__31570),
            .in1(N__22120),
            .in2(N__22099),
            .in3(N__22035),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_7_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_7_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_7_17_0  (
            .in0(N__23275),
            .in1(N__20893),
            .in2(N__23465),
            .in3(N__23224),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_7_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_7_17_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_7_17_1  (
            .in0(N__25537),
            .in1(N__22061),
            .in2(_gnd_net_),
            .in3(N__24805),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_7_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_7_17_2 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_7_17_2  (
            .in0(N__22036),
            .in1(N__20711),
            .in2(N__20675),
            .in3(N__20740),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_7_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_7_17_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_7_17_3  (
            .in0(N__23527),
            .in1(N__23554),
            .in2(_gnd_net_),
            .in3(N__23497),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_7_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_7_17_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_7_17_4  (
            .in0(N__20872),
            .in1(N__23590),
            .in2(N__20672),
            .in3(N__20669),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_7_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_7_17_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_7_17_5  (
            .in0(N__20794),
            .in1(N__20818),
            .in2(N__20773),
            .in3(N__20839),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_7_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_7_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_7_17_6  (
            .in0(N__24804),
            .in1(N__25536),
            .in2(N__20705),
            .in3(N__20739),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_7_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_7_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_7_18_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(N__22242),
            .in2(N__23696),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_7_18_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__44886),
            .ce(N__23653),
            .sr(N__44219));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_7_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_7_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_7_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(N__22218),
            .in2(N__23675),
            .in3(N__20702),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__44886),
            .ce(N__23653),
            .sr(N__44219));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_7_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_7_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_7_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_7_18_2  (
            .in0(_gnd_net_),
            .in1(N__22194),
            .in2(N__22247),
            .in3(N__20699),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__44886),
            .ce(N__23653),
            .sr(N__44219));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_7_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_7_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_7_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(N__22563),
            .in2(N__22223),
            .in3(N__20696),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__44886),
            .ce(N__23653),
            .sr(N__44219));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_7_18_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_7_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_7_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(N__22542),
            .in2(N__22199),
            .in3(N__20693),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__44886),
            .ce(N__23653),
            .sr(N__44219));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_7_18_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_7_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_7_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(N__22524),
            .in2(N__22568),
            .in3(N__20690),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__44886),
            .ce(N__23653),
            .sr(N__44219));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_7_18_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_7_18_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_7_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(N__22543),
            .in2(N__22508),
            .in3(N__20687),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__44886),
            .ce(N__23653),
            .sr(N__44219));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_7_18_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_7_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_7_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_7_18_7  (
            .in0(_gnd_net_),
            .in1(N__22525),
            .in2(N__22475),
            .in3(N__20828),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__44886),
            .ce(N__23653),
            .sr(N__44219));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_7_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_7_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_7_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__22440),
            .in2(N__22504),
            .in3(N__20801),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__44878),
            .ce(N__23652),
            .sr(N__44225));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_7_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_7_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_7_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__22416),
            .in2(N__22474),
            .in3(N__20777),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__44878),
            .ce(N__23652),
            .sr(N__44225));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_7_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_7_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_7_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__22392),
            .in2(N__22445),
            .in3(N__20750),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__44878),
            .ce(N__23652),
            .sr(N__44225));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_7_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_7_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_7_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__22755),
            .in2(N__22421),
            .in3(N__20747),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__44878),
            .ce(N__23652),
            .sr(N__44225));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_7_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_7_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_7_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__22734),
            .in2(N__22397),
            .in3(N__20723),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__44878),
            .ce(N__23652),
            .sr(N__44225));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_7_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_7_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__22716),
            .in2(N__22760),
            .in3(N__20720),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__44878),
            .ce(N__23652),
            .sr(N__44225));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_7_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_7_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__22735),
            .in2(N__22700),
            .in3(N__20717),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__44878),
            .ce(N__23652),
            .sr(N__44225));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_7_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_7_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_7_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__22717),
            .in2(N__22670),
            .in3(N__20714),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__44878),
            .ce(N__23652),
            .sr(N__44225));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_7_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_7_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_7_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__22635),
            .in2(N__22699),
            .in3(N__20912),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__44872),
            .ce(N__23651),
            .sr(N__44230));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_7_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_7_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_7_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__22611),
            .in2(N__22669),
            .in3(N__20909),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__44872),
            .ce(N__23651),
            .sr(N__44230));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_7_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_7_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_7_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(N__22587),
            .in2(N__22640),
            .in3(N__20906),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__44872),
            .ce(N__23651),
            .sr(N__44230));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_7_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_7_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_7_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(N__22953),
            .in2(N__22616),
            .in3(N__20903),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__44872),
            .ce(N__23651),
            .sr(N__44230));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_7_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_7_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(N__22932),
            .in2(N__22592),
            .in3(N__20879),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__44872),
            .ce(N__23651),
            .sr(N__44230));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_7_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_7_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(N__22914),
            .in2(N__22958),
            .in3(N__20858),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__44872),
            .ce(N__23651),
            .sr(N__44230));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_7_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_7_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(N__22933),
            .in2(N__22898),
            .in3(N__20855),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__44872),
            .ce(N__23651),
            .sr(N__44230));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_7_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_7_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(N__22915),
            .in2(N__22868),
            .in3(N__20852),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__44872),
            .ce(N__23651),
            .sr(N__44230));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_7_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_7_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_7_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__22833),
            .in2(N__22897),
            .in3(N__20849),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__44865),
            .ce(N__23650),
            .sr(N__44233));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_7_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_7_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_7_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__22809),
            .in2(N__22867),
            .in3(N__20990),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__44865),
            .ce(N__23650),
            .sr(N__44233));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_7_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_7_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_7_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(N__22789),
            .in2(N__22838),
            .in3(N__20987),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__44865),
            .ce(N__23650),
            .sr(N__44233));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_7_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_7_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_7_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(N__22771),
            .in2(N__22814),
            .in3(N__20984),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__44865),
            .ce(N__23650),
            .sr(N__44233));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_7_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_7_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_7_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_7_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20981),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44865),
            .ce(N__23650),
            .sr(N__44233));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_7_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_7_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_8_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20978),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44937),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_8_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_8_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__23069),
            .in2(N__32414),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__44921),
            .ce(),
            .sr(N__44152));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_8_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_8_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_8_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__25028),
            .in2(N__32345),
            .in3(N__20933),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__44921),
            .ce(),
            .sr(N__44152));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_8_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_8_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__34490),
            .in2(N__23108),
            .in3(N__20915),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__44921),
            .ce(),
            .sr(N__44152));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_8_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_8_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__23090),
            .in2(N__32255),
            .in3(N__21242),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__44921),
            .ce(),
            .sr(N__44152));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_8_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_8_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__30302),
            .in2(N__23099),
            .in3(N__21203),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__44921),
            .ce(),
            .sr(N__44152));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_8_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_8_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__31268),
            .in2(N__23084),
            .in3(N__21167),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__44921),
            .ce(),
            .sr(N__44152));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_8_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_8_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__23882),
            .in2(N__34649),
            .in3(N__21131),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__44921),
            .ce(),
            .sr(N__44152));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_8_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_8_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_8_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__23075),
            .in2(N__30647),
            .in3(N__21098),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__44921),
            .ce(),
            .sr(N__44152));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_8_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_8_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__25274),
            .in2(N__30443),
            .in3(N__21056),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__44915),
            .ce(),
            .sr(N__44159));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_8_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_8_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__23873),
            .in2(N__31100),
            .in3(N__21023),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__44915),
            .ce(),
            .sr(N__44159));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_8_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_8_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__25265),
            .in2(N__35333),
            .in3(N__21011),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__44915),
            .ce(),
            .sr(N__44159));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_8_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_8_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__23063),
            .in2(N__34232),
            .in3(N__20993),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__44915),
            .ce(),
            .sr(N__44159));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_8_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_8_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__22994),
            .in2(N__30536),
            .in3(N__21398),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__44915),
            .ce(),
            .sr(N__44159));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_8_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_8_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__30907),
            .in2(N__23035),
            .in3(N__21386),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__44915),
            .ce(),
            .sr(N__44159));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_8_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_8_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__22998),
            .in2(N__34397),
            .in3(N__21368),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__44915),
            .ce(),
            .sr(N__44159));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_8_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_8_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__30383),
            .in2(N__23036),
            .in3(N__21347),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__44915),
            .ce(),
            .sr(N__44159));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_8_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_8_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__30809),
            .in2(N__23037),
            .in3(N__21326),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__44912),
            .ce(),
            .sr(N__44164));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_8_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_8_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__23005),
            .in2(N__31013),
            .in3(N__21311),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__44912),
            .ce(),
            .sr(N__44164));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_8_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_8_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_8_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__30707),
            .in2(N__23038),
            .in3(N__21290),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__44912),
            .ce(),
            .sr(N__44164));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_8_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_8_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__23009),
            .in2(N__34346),
            .in3(N__21278),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__44912),
            .ce(),
            .sr(N__44164));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_8_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_8_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_8_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__32618),
            .in2(N__23039),
            .in3(N__21569),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__44912),
            .ce(),
            .sr(N__44164));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_8_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_8_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__23013),
            .in2(N__32564),
            .in3(N__21548),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__44912),
            .ce(),
            .sr(N__44164));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_8_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_8_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_8_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__32510),
            .in2(N__23040),
            .in3(N__21530),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__44912),
            .ce(),
            .sr(N__44164));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_8_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_8_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_8_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__23017),
            .in2(N__35228),
            .in3(N__21518),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__44912),
            .ce(),
            .sr(N__44164));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_8_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_8_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__23041),
            .in2(N__35171),
            .in3(N__21500),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__44908),
            .ce(),
            .sr(N__44174));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_8_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_8_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__35111),
            .in2(N__23055),
            .in3(N__21485),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__44908),
            .ce(),
            .sr(N__44174));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_8_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_8_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__23045),
            .in2(N__35054),
            .in3(N__21464),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__44908),
            .ce(),
            .sr(N__44174));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_8_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_8_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__28664),
            .in2(N__23056),
            .in3(N__21440),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__44908),
            .ce(),
            .sr(N__44174));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_8_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_8_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__23049),
            .in2(N__34595),
            .in3(N__21419),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__44908),
            .ce(),
            .sr(N__44174));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_8_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_8_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__34532),
            .in2(N__23057),
            .in3(N__21707),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__44908),
            .ce(),
            .sr(N__44174));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_8_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_8_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__23053),
            .in2(N__35885),
            .in3(N__21683),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__44908),
            .ce(),
            .sr(N__44174));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_8_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_8_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_8_13_7  (
            .in0(N__23054),
            .in1(N__35834),
            .in2(_gnd_net_),
            .in3(N__21680),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44908),
            .ce(),
            .sr(N__44174));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_14_LC_8_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_14_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_14_LC_8_14_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_14_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__24891),
            .in2(_gnd_net_),
            .in3(N__24404),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__25256),
            .in2(_gnd_net_),
            .in3(N__25202),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_1_9_LC_8_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_1_9_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_1_9_LC_8_14_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_i_1_9_LC_8_14_5  (
            .in0(N__21895),
            .in1(N__24701),
            .in2(_gnd_net_),
            .in3(N__21816),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_8_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_8_14_6 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_8_14_6  (
            .in0(N__31854),
            .in1(N__23416),
            .in2(N__31650),
            .in3(N__22151),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_8_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_8_14_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_8_14_7  (
            .in0(N__24542),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25464),
            .lcout(elapsed_time_ns_1_RNI62CED1_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_14_LC_8_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_14_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_14_LC_8_15_0 .LUT_INIT=16'b0000000011111011;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_14_LC_8_15_0  (
            .in0(N__21934),
            .in1(N__21589),
            .in2(N__24727),
            .in3(N__26010),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44897),
            .ce(N__31527),
            .sr(N__44184));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_9_LC_8_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_9_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_9_LC_8_15_1 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_9_LC_8_15_1  (
            .in0(N__26011),
            .in1(N__21868),
            .in2(N__24439),
            .in3(N__24699),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44897),
            .ce(N__31527),
            .sr(N__44184));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_15_LC_8_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_15_LC_8_15_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_15_LC_8_15_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_15_LC_8_15_2  (
            .in0(N__24881),
            .in1(N__26015),
            .in2(N__24726),
            .in3(N__24409),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44897),
            .ce(N__31527),
            .sr(N__44184));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_18_LC_8_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_18_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_18_LC_8_15_3 .LUT_INIT=16'b0000111000001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_18_LC_8_15_3  (
            .in0(N__23375),
            .in1(N__24691),
            .in2(N__26037),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44897),
            .ce(N__31527),
            .sr(N__44184));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_17_LC_8_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_17_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_17_LC_8_15_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_17_LC_8_15_4  (
            .in0(N__24688),
            .in1(N__26008),
            .in2(_gnd_net_),
            .in3(N__23411),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44897),
            .ce(N__31527),
            .sr(N__44184));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_16_LC_8_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_16_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_16_LC_8_15_5 .LUT_INIT=16'b0000111000001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_16_LC_8_15_5  (
            .in0(N__23341),
            .in1(N__24690),
            .in2(N__26036),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44897),
            .ce(N__31527),
            .sr(N__44184));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_10_LC_8_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_10_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_10_LC_8_15_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_10_LC_8_15_6  (
            .in0(N__24689),
            .in1(N__26009),
            .in2(N__21857),
            .in3(N__21826),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44897),
            .ce(N__31527),
            .sr(N__44184));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_11_LC_8_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_11_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_11_LC_8_15_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_11_LC_8_15_7  (
            .in0(N__21825),
            .in1(N__24692),
            .in2(N__26035),
            .in3(N__21781),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44897),
            .ce(N__31527),
            .sr(N__44184));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_0_15_LC_8_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_0_15_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_0_15_LC_8_16_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_i_o5_0_15_LC_8_16_0  (
            .in0(N__21757),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21745),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_i_o5_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_8_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_8_16_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_8_16_1  (
            .in0(N__44321),
            .in1(N__22340),
            .in2(N__22325),
            .in3(N__23739),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_8_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_8_16_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_8_16_2  (
            .in0(N__44326),
            .in1(N__24522),
            .in2(N__21977),
            .in3(N__21986),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_8_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_8_16_3 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_8_16_3  (
            .in0(N__21974),
            .in1(_gnd_net_),
            .in2(N__21965),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNI40CED1_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1_6_LC_8_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1_6_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1_6_LC_8_16_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1_6_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__21922),
            .in2(_gnd_net_),
            .in3(N__24868),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_f0_i_o2_a1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_8_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_8_16_5 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_8_16_5  (
            .in0(N__24523),
            .in1(N__22276),
            .in2(N__44338),
            .in3(N__23771),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_8_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_8_16_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_8_16_6  (
            .in0(N__23740),
            .in1(N__44322),
            .in2(N__21962),
            .in3(N__22175),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_8_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_8_16_7 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_8_16_7  (
            .in0(N__26120),
            .in1(N__31808),
            .in2(N__21959),
            .in3(N__22361),
            .lcout(elapsed_time_ns_1_RNIB4DJ11_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_8_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_8_17_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__23712),
            .in2(_gnd_net_),
            .in3(N__26248),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_8_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_8_17_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__25448),
            .in2(_gnd_net_),
            .in3(N__21950),
            .lcout(elapsed_time_ns_1_RNI1TBED1_0_14),
            .ltout(elapsed_time_ns_1_RNI1TBED1_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_9_LC_8_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_9_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_9_LC_8_17_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_9_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__24864),
            .in2(N__21899),
            .in3(N__21887),
            .lcout(\phase_controller_inst1.stoper_hc.N_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_8_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_8_17_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_8_17_3  (
            .in0(N__44331),
            .in1(N__24526),
            .in2(_gnd_net_),
            .in3(N__22294),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_8_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_8_17_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_8_17_4  (
            .in0(N__24571),
            .in1(N__22150),
            .in2(N__22169),
            .in3(N__22160),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_8_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_8_17_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22154),
            .in3(N__23752),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_382_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_8_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_8_17_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_8_17_6  (
            .in0(N__23299),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23197),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_8_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_8_17_7 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_8_17_7  (
            .in0(N__25368),
            .in1(N__31809),
            .in2(N__26394),
            .in3(N__22373),
            .lcout(elapsed_time_ns_1_RNIA3DJ11_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_18_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_18_0  (
            .in0(N__22137),
            .in1(N__22114),
            .in2(N__22098),
            .in3(N__24564),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_8_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_8_18_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_8_18_1  (
            .in0(N__22065),
            .in1(N__22034),
            .in2(N__22010),
            .in3(N__31566),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_8_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_8_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_8_18_2  (
            .in0(N__22317),
            .in1(N__44333),
            .in2(N__22007),
            .in3(N__22003),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_8_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_8_18_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_8_18_3  (
            .in0(N__22339),
            .in1(_gnd_net_),
            .in2(N__21989),
            .in3(N__23766),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_8_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_8_18_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__22372),
            .in2(_gnd_net_),
            .in3(N__22357),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_8_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_8_18_5 .LUT_INIT=16'b0011001000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_8_18_5  (
            .in0(N__22298),
            .in1(N__24525),
            .in2(N__22280),
            .in3(N__23767),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_8_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_8_18_6 .LUT_INIT=16'b1110111111001111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_8_18_6  (
            .in0(N__22346),
            .in1(N__22338),
            .in2(N__22324),
            .in3(N__22304),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_8_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_8_18_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__24524),
            .in2(N__22283),
            .in3(N__22269),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_19_0  (
            .in0(N__29030),
            .in1(N__23691),
            .in2(_gnd_net_),
            .in3(N__22253),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__44873),
            .ce(N__25595),
            .sr(N__44220));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_19_1  (
            .in0(N__29003),
            .in1(N__23670),
            .in2(_gnd_net_),
            .in3(N__22250),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__44873),
            .ce(N__25595),
            .sr(N__44220));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_19_2  (
            .in0(N__29031),
            .in1(N__22243),
            .in2(_gnd_net_),
            .in3(N__22226),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__44873),
            .ce(N__25595),
            .sr(N__44220));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_19_3  (
            .in0(N__29004),
            .in1(N__22219),
            .in2(_gnd_net_),
            .in3(N__22202),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__44873),
            .ce(N__25595),
            .sr(N__44220));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_19_4  (
            .in0(N__29032),
            .in1(N__22195),
            .in2(_gnd_net_),
            .in3(N__22178),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__44873),
            .ce(N__25595),
            .sr(N__44220));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_19_5  (
            .in0(N__29005),
            .in1(N__22564),
            .in2(_gnd_net_),
            .in3(N__22547),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__44873),
            .ce(N__25595),
            .sr(N__44220));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_19_6  (
            .in0(N__29033),
            .in1(N__22544),
            .in2(_gnd_net_),
            .in3(N__22529),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__44873),
            .ce(N__25595),
            .sr(N__44220));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_19_7  (
            .in0(N__29006),
            .in1(N__22526),
            .in2(_gnd_net_),
            .in3(N__22511),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__44873),
            .ce(N__25595),
            .sr(N__44220));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_20_0  (
            .in0(N__28977),
            .in1(N__22497),
            .in2(_gnd_net_),
            .in3(N__22478),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__44866),
            .ce(N__25596),
            .sr(N__44226));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_20_1  (
            .in0(N__29002),
            .in1(N__22467),
            .in2(_gnd_net_),
            .in3(N__22448),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__44866),
            .ce(N__25596),
            .sr(N__44226));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_20_2  (
            .in0(N__28974),
            .in1(N__22441),
            .in2(_gnd_net_),
            .in3(N__22424),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__44866),
            .ce(N__25596),
            .sr(N__44226));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_20_3  (
            .in0(N__28999),
            .in1(N__22417),
            .in2(_gnd_net_),
            .in3(N__22400),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__44866),
            .ce(N__25596),
            .sr(N__44226));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_20_4  (
            .in0(N__28975),
            .in1(N__22393),
            .in2(_gnd_net_),
            .in3(N__22376),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__44866),
            .ce(N__25596),
            .sr(N__44226));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_20_5  (
            .in0(N__29000),
            .in1(N__22756),
            .in2(_gnd_net_),
            .in3(N__22739),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__44866),
            .ce(N__25596),
            .sr(N__44226));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_20_6  (
            .in0(N__28976),
            .in1(N__22736),
            .in2(_gnd_net_),
            .in3(N__22721),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__44866),
            .ce(N__25596),
            .sr(N__44226));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_20_7  (
            .in0(N__29001),
            .in1(N__22718),
            .in2(_gnd_net_),
            .in3(N__22703),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__44866),
            .ce(N__25596),
            .sr(N__44226));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_21_0  (
            .in0(N__29007),
            .in1(N__22692),
            .in2(_gnd_net_),
            .in3(N__22673),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__44859),
            .ce(N__25607),
            .sr(N__44231));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_21_1  (
            .in0(N__29013),
            .in1(N__22662),
            .in2(_gnd_net_),
            .in3(N__22643),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__44859),
            .ce(N__25607),
            .sr(N__44231));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_21_2  (
            .in0(N__29008),
            .in1(N__22636),
            .in2(_gnd_net_),
            .in3(N__22619),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__44859),
            .ce(N__25607),
            .sr(N__44231));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_21_3  (
            .in0(N__29014),
            .in1(N__22612),
            .in2(_gnd_net_),
            .in3(N__22595),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__44859),
            .ce(N__25607),
            .sr(N__44231));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_21_4  (
            .in0(N__29009),
            .in1(N__22588),
            .in2(_gnd_net_),
            .in3(N__22571),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__44859),
            .ce(N__25607),
            .sr(N__44231));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_21_5  (
            .in0(N__29015),
            .in1(N__22954),
            .in2(_gnd_net_),
            .in3(N__22937),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__44859),
            .ce(N__25607),
            .sr(N__44231));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_21_6  (
            .in0(N__29010),
            .in1(N__22934),
            .in2(_gnd_net_),
            .in3(N__22919),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__44859),
            .ce(N__25607),
            .sr(N__44231));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_21_7  (
            .in0(N__29016),
            .in1(N__22916),
            .in2(_gnd_net_),
            .in3(N__22901),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__44859),
            .ce(N__25607),
            .sr(N__44231));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_22_0  (
            .in0(N__29017),
            .in1(N__22890),
            .in2(_gnd_net_),
            .in3(N__22871),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__44856),
            .ce(N__25606),
            .sr(N__44234));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_22_1  (
            .in0(N__29011),
            .in1(N__22860),
            .in2(_gnd_net_),
            .in3(N__22841),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__44856),
            .ce(N__25606),
            .sr(N__44234));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_22_2  (
            .in0(N__29018),
            .in1(N__22834),
            .in2(_gnd_net_),
            .in3(N__22817),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__44856),
            .ce(N__25606),
            .sr(N__44234));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_22_3  (
            .in0(N__29012),
            .in1(N__22810),
            .in2(_gnd_net_),
            .in3(N__22793),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__44856),
            .ce(N__25606),
            .sr(N__44234));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_22_4  (
            .in0(N__29019),
            .in1(N__22790),
            .in2(_gnd_net_),
            .in3(N__22778),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__44856),
            .ce(N__25606),
            .sr(N__44234));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_22_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_22_5  (
            .in0(N__22772),
            .in1(N__29020),
            .in2(_gnd_net_),
            .in3(N__22775),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44856),
            .ce(N__25606),
            .sr(N__44234));
    defparam \phase_controller_inst2.S2_LC_8_30_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_8_30_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_8_30_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_8_30_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26603),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44833),
            .ce(),
            .sr(N__44239));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_9_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_9_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28427),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44916),
            .ce(),
            .sr(N__44146));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_9_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_9_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_9_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28277),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44916),
            .ce(),
            .sr(N__44146));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_9_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_9_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28400),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44916),
            .ce(),
            .sr(N__44146));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_9_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_9_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26909),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44916),
            .ce(),
            .sr(N__44146));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_9_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_9_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28298),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44916),
            .ce(),
            .sr(N__44146));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_9_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_9_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28256),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44913),
            .ce(),
            .sr(N__44153));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_9_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_9_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30250),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44913),
            .ce(),
            .sr(N__44153));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_9_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_9_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34942),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44913),
            .ce(),
            .sr(N__44153));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__23144),
            .in2(N__25157),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__23828),
            .in2(_gnd_net_),
            .in3(N__23138),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(N__44904),
            .ce(),
            .sr(N__25130));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__23807),
            .in2(N__25016),
            .in3(N__23135),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(N__44904),
            .ce(),
            .sr(N__25130));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__24134),
            .in2(_gnd_net_),
            .in3(N__23132),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(N__44904),
            .ce(),
            .sr(N__25130));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__24110),
            .in2(_gnd_net_),
            .in3(N__23129),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(N__44904),
            .ce(),
            .sr(N__25130));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__24086),
            .in2(_gnd_net_),
            .in3(N__23126),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(N__44904),
            .ce(),
            .sr(N__25130));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__24050),
            .in2(_gnd_net_),
            .in3(N__23123),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(N__44904),
            .ce(),
            .sr(N__25130));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__24029),
            .in2(_gnd_net_),
            .in3(N__23120),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(N__44904),
            .ce(),
            .sr(N__25130));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_9_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_9_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__23993),
            .in2(_gnd_net_),
            .in3(N__23117),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(N__44898),
            .ce(),
            .sr(N__25126));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_9_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_9_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__23960),
            .in2(_gnd_net_),
            .in3(N__23171),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(N__44898),
            .ce(),
            .sr(N__25126));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__23939),
            .in2(_gnd_net_),
            .in3(N__23168),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(N__44898),
            .ce(),
            .sr(N__25126));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__24374),
            .in2(_gnd_net_),
            .in3(N__23165),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(N__44898),
            .ce(),
            .sr(N__25126));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__24326),
            .in2(_gnd_net_),
            .in3(N__23162),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(N__44898),
            .ce(),
            .sr(N__25126));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__24305),
            .in2(_gnd_net_),
            .in3(N__23159),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(N__44898),
            .ce(),
            .sr(N__25126));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__24263),
            .in2(_gnd_net_),
            .in3(N__23156),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(N__44898),
            .ce(),
            .sr(N__25126));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__24230),
            .in2(_gnd_net_),
            .in3(N__23153),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(N__44898),
            .ce(),
            .sr(N__25126));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__24191),
            .in2(_gnd_net_),
            .in3(N__23150),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(N__44892),
            .ce(),
            .sr(N__25118));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__24155),
            .in2(_gnd_net_),
            .in3(N__23147),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(N__44892),
            .ce(),
            .sr(N__25118));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__24605),
            .in2(_gnd_net_),
            .in3(N__23423),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44892),
            .ce(),
            .sr(N__25118));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3_2_LC_9_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3_2_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3_2_LC_9_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3_2_LC_9_16_0  (
            .in0(N__23401),
            .in1(N__25361),
            .in2(N__26121),
            .in3(N__23377),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_2_LC_9_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_2_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_2_LC_9_16_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_i_a2_1_2_LC_9_16_1  (
            .in0(N__24474),
            .in1(N__23345),
            .in2(N__23315),
            .in3(N__23312),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_9_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_9_16_2 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_9_16_2  (
            .in0(N__31802),
            .in1(N__23252),
            .in2(N__26381),
            .in3(N__23306),
            .lcout(elapsed_time_ns_1_RNIP2ND11_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_9_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_9_16_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_9_16_3  (
            .in0(N__23258),
            .in1(N__26348),
            .in2(N__23285),
            .in3(N__31801),
            .lcout(elapsed_time_ns_1_RNI1BND11_0_29),
            .ltout(elapsed_time_ns_1_RNI1BND11_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_7_15_LC_9_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_7_15_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_7_15_LC_9_16_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_i_o5_7_15_LC_9_16_4  (
            .in0(N__23438),
            .in1(N__23251),
            .in2(N__23243),
            .in3(N__23209),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_7_i_o5_7Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_15_LC_9_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_15_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_15_LC_9_16_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_i_o5_15_LC_9_16_5  (
            .in0(N__23240),
            .in1(N__23179),
            .in2(N__23234),
            .in3(N__23561),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_i_o5Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_9_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_9_16_6 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_9_16_6  (
            .in0(N__31803),
            .in1(N__23210),
            .in2(N__26382),
            .in3(N__23231),
            .lcout(elapsed_time_ns_1_RNIO1ND11_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_9_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_9_16_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_9_16_7  (
            .in0(N__23201),
            .in1(N__23180),
            .in2(N__26398),
            .in3(N__31804),
            .lcout(elapsed_time_ns_1_RNIQ3ND11_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_4_LC_9_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_4_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_4_LC_9_17_0 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_4_LC_9_17_0  (
            .in0(N__25939),
            .in1(N__25799),
            .in2(N__25372),
            .in3(N__25728),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44879),
            .ce(N__31529),
            .sr(N__44189));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_9_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_9_17_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_9_17_1  (
            .in0(N__26333),
            .in1(N__31771),
            .in2(N__23573),
            .in3(N__23594),
            .lcout(elapsed_time_ns_1_RNIT6ND11_0_25),
            .ltout(elapsed_time_ns_1_RNIT6ND11_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_6_15_LC_9_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_6_15_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_o5_6_15_LC_9_17_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_i_o5_6_15_LC_9_17_2  (
            .in0(N__23476),
            .in1(N__23536),
            .in2(N__23564),
            .in3(N__23509),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_i_o5_6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_9_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_9_17_3 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_9_17_3  (
            .in0(N__23537),
            .in1(N__23555),
            .in2(N__26374),
            .in3(N__31774),
            .lcout(elapsed_time_ns_1_RNIV8ND11_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_9_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_9_17_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_9_17_4  (
            .in0(N__31772),
            .in1(N__23528),
            .in2(N__26396),
            .in3(N__23510),
            .lcout(elapsed_time_ns_1_RNIU7ND11_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_9_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_9_17_5 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_9_17_5  (
            .in0(N__26334),
            .in1(N__23501),
            .in2(N__23480),
            .in3(N__31773),
            .lcout(elapsed_time_ns_1_RNI0AND11_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_5_LC_9_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_5_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_5_LC_9_17_6 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_5_LC_9_17_6  (
            .in0(N__25940),
            .in1(N__25800),
            .in2(N__26125),
            .in3(N__25729),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44879),
            .ce(N__31529),
            .sr(N__44189));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_9_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_9_18_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_9_18_0  (
            .in0(N__31799),
            .in1(N__23464),
            .in2(N__26395),
            .in3(N__23437),
            .lcout(elapsed_time_ns_1_RNIP3OD11_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_9_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_9_18_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_9_18_1  (
            .in0(N__23785),
            .in1(N__25486),
            .in2(N__23723),
            .in3(N__26244),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_9_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_9_18_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_9_18_4  (
            .in0(N__44332),
            .in1(N__23753),
            .in2(_gnd_net_),
            .in3(N__23741),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_9_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_9_18_5 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_9_18_5  (
            .in0(N__26204),
            .in1(N__31800),
            .in2(N__23726),
            .in3(N__23722),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_9_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_9_18_6 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23699),
            .in3(N__31608),
            .lcout(elapsed_time_ns_1_RNIQURR91_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23695),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44867),
            .ce(N__23654),
            .sr(N__44210));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23674),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44867),
            .ce(N__23654),
            .sr(N__44210));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_9_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_9_20_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_9_20_1  (
            .in0(N__29065),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29104),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_432_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_9_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_9_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_1_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__27895),
            .in2(_gnd_net_),
            .in3(N__24927),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_9_20_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_9_20_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_9_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_9_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23612),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44860),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S1_LC_9_28_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_28_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_28_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_28_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27907),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44836),
            .ce(),
            .sr(N__44238));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_6_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_6_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_10_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23897),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44928),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_10_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_10_10_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_10_10_4  (
            .in0(N__34453),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44909),
            .ce(),
            .sr(N__44135));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_10_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_10_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_10_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31226),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44905),
            .ce(),
            .sr(N__44143));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_12_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_12_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_10_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23864),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44899),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_10_12_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_10_12_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_10_12_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_10_12_5 (
            .in0(N__23855),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44899),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__25817),
            .in2(N__23837),
            .in3(N__25146),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__25388),
            .in2(N__23816),
            .in3(N__23827),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_13_2  (
            .in0(N__23806),
            .in1(N__25661),
            .in2(N__23795),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_13_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_13_3  (
            .in0(N__24133),
            .in1(N__25340),
            .in2(N__24122),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__26090),
            .in2(N__24098),
            .in3(N__24109),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_13_5  (
            .in0(N__24085),
            .in1(N__25415),
            .in2(N__24074),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__24062),
            .in2(N__24038),
            .in3(N__24049),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__26051),
            .in2(N__24017),
            .in3(N__24028),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__24005),
            .in2(N__23981),
            .in3(N__23992),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__23972),
            .in2(N__23948),
            .in3(N__23959),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_14_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_14_2  (
            .in0(N__23938),
            .in1(N__23927),
            .in2(N__23915),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_14_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_14_3  (
            .in0(N__24373),
            .in1(N__24362),
            .in2(N__24350),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__24341),
            .in2(N__24314),
            .in3(N__24325),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_14_5  (
            .in0(N__24304),
            .in1(N__24281),
            .in2(N__24293),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__24275),
            .in2(N__24251),
            .in3(N__24262),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__24242),
            .in2(N__24218),
            .in3(N__24229),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__24206),
            .in2(N__24179),
            .in3(N__24190),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__24170),
            .in2(N__24143),
            .in3(N__24154),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__24620),
            .in2(N__24593),
            .in3(N__24604),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24584),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_15_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_15_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_15_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_10_15_5 (
            .in0(N__24581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44881),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_10_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_10_16_0 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_10_16_0  (
            .in0(N__31859),
            .in1(N__24482),
            .in2(N__31658),
            .in3(N__24572),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_10_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_10_16_1 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_10_16_1  (
            .in0(N__24530),
            .in1(N__26390),
            .in2(N__26022),
            .in3(N__31858),
            .lcout(elapsed_time_ns_1_RNIQ4OD11_0_31),
            .ltout(elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_19_LC_10_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_19_LC_10_16_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_19_LC_10_16_2 .LUT_INIT=16'b0000111000001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_19_LC_10_16_2  (
            .in0(N__24674),
            .in1(N__24481),
            .in2(N__24443),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44874),
            .ce(N__31526),
            .sr(N__44175));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_3_LC_10_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_3_LC_10_16_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_3_LC_10_16_5 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_3_LC_10_16_5  (
            .in0(N__25785),
            .in1(N__26209),
            .in2(N__25733),
            .in3(N__25673),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44874),
            .ce(N__31526),
            .sr(N__44175));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_0_6_LC_10_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_0_6_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_0_6_LC_10_16_6 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_0_6_LC_10_16_6  (
            .in0(N__24440),
            .in1(N__24413),
            .in2(N__24700),
            .in3(N__24383),
            .lcout(\phase_controller_inst1.stoper_hc.N_325 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_6_LC_10_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_6_LC_10_16_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_6_LC_10_16_7 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_6_LC_10_16_7  (
            .in0(N__25981),
            .in1(N__31683),
            .in2(N__24908),
            .in3(N__25730),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44874),
            .ce(N__31526),
            .sr(N__44175));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0_2_LC_10_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0_2_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0_2_LC_10_17_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_i_a2_0_2_LC_10_17_0  (
            .in0(N__25515),
            .in1(N__31679),
            .in2(N__26077),
            .in3(N__24905),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_7_i_a2_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_6_LC_10_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_6_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_6_LC_10_17_1 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_i_a2_6_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__24892),
            .in2(N__24821),
            .in3(N__24668),
            .lcout(\phase_controller_inst1.stoper_hc.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_0_2_LC_10_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_0_2_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_i_0_2_LC_10_17_2 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_i_0_2_LC_10_17_2  (
            .in0(N__24771),
            .in1(N__26200),
            .in2(N__24791),
            .in3(N__26225),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_i_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_a5_1_LC_10_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_a5_1_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_a5_1_LC_10_17_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_0_a5_1_LC_10_17_3  (
            .in0(N__24786),
            .in1(N__26171),
            .in2(N__24772),
            .in3(N__24669),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.N_307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_1_1_LC_10_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_1_1_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_1_1_LC_10_17_4 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_0_1_1_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__25714),
            .in2(N__24818),
            .in3(N__25845),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_f0_0_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_17_5 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_17_5  (
            .in0(N__31835),
            .in1(N__26399),
            .in2(N__24815),
            .in3(N__26072),
            .lcout(elapsed_time_ns_1_RNIE7DJ11_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_10_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_10_17_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__31547),
            .in2(_gnd_net_),
            .in3(N__25472),
            .lcout(elapsed_time_ns_1_RNIIU2KD1_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_0_3_LC_10_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_0_3_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_0_3_LC_10_17_7 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_0_0_3_LC_10_17_7  (
            .in0(N__24787),
            .in1(N__25911),
            .in2(N__24773),
            .in3(N__24670),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_7_f0_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNI41671_0_1_LC_10_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNI41671_0_1_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNI41671_0_1_LC_10_18_0 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNI41671_0_1_LC_10_18_0  (
            .in0(N__24970),
            .in1(N__44327),
            .in2(N__25248),
            .in3(N__24996),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUB_LC_10_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUB_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUB_LC_10_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUB_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__25234),
            .in2(_gnd_net_),
            .in3(N__25194),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIGEUBZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_10_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_10_18_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_10_18_4 .LUT_INIT=16'b0101000000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_10_18_4  (
            .in0(N__25239),
            .in1(N__25199),
            .in2(N__24977),
            .in3(N__24997),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44861),
            .ce(),
            .sr(N__44185));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNI41671_1_LC_10_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNI41671_1_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNI41671_1_LC_10_18_5 .LUT_INIT=16'b1111000011110110;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNI41671_1_LC_10_18_5  (
            .in0(N__24994),
            .in1(N__24969),
            .in2(N__44339),
            .in3(N__25235),
            .lcout(\phase_controller_inst1.stoper_hc.un1_stoper_state12_1_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_18_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_18_6  (
            .in0(N__24971),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24995),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.N_45_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_10_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_10_18_7 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_10_18_7  (
            .in0(N__36623),
            .in1(N__25240),
            .in2(N__25001),
            .in3(N__25195),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44861),
            .ce(),
            .sr(N__44185));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_10_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_10_19_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_10_19_4  (
            .in0(N__24998),
            .in1(N__25244),
            .in2(N__24976),
            .in3(N__25200),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44857),
            .ce(),
            .sr(N__44199));
    defparam \phase_controller_inst1.start_timer_hc_LC_10_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_10_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_10_20_2 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_10_20_2  (
            .in0(N__26665),
            .in1(N__26135),
            .in2(N__24975),
            .in3(N__36572),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44852),
            .ce(),
            .sr(N__44208));
    defparam \phase_controller_inst2.state_2_LC_10_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_10_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_10_21_0 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst2.state_2_LC_10_21_0  (
            .in0(N__24937),
            .in1(N__28011),
            .in2(N__27905),
            .in3(N__26447),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44848),
            .ce(),
            .sr(N__44214));
    defparam \phase_controller_inst2.state_3_LC_10_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_10_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_10_22_3 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst2.state_3_LC_10_22_3  (
            .in0(N__27891),
            .in1(N__28037),
            .in2(N__24938),
            .in3(N__25051),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44845),
            .ce(),
            .sr(N__44221));
    defparam \phase_controller_inst2.T12_LC_10_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.T12_LC_10_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T12_LC_10_22_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \phase_controller_inst2.T12_LC_10_22_5  (
            .in0(N__26590),
            .in1(N__28015),
            .in2(_gnd_net_),
            .in3(N__25063),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44845),
            .ce(),
            .sr(N__44221));
    defparam \phase_controller_inst1.state_3_LC_10_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_10_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_10_22_7 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst1.state_3_LC_10_22_7  (
            .in0(N__28838),
            .in1(N__25052),
            .in2(N__28895),
            .in3(N__26162),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44845),
            .ce(),
            .sr(N__44221));
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_10_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_10_23_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a3_1_LC_10_23_1  (
            .in0(N__26701),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26650),
            .lcout(state_ns_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_11_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_11_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29135),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25042),
            .ce(),
            .sr(N__44122));
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29136),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25043),
            .ce(),
            .sr(N__44124));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_11_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_11_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_11_9_1  (
            .in0(N__30432),
            .in1(N__34644),
            .in2(N__31096),
            .in3(N__30643),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_11_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_11_9_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_11_9_2  (
            .in0(N__30301),
            .in1(N__32247),
            .in2(N__25031),
            .in3(N__31263),
            .lcout(\current_shift_inst.PI_CTRL.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_11_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_11_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34528),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26797),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44900),
            .ce(),
            .sr(N__44136));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_11_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_11_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28232),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44900),
            .ce(),
            .sr(N__44136));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_11_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_11_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30334),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44900),
            .ce(),
            .sr(N__44136));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_11_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34986),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44900),
            .ce(),
            .sr(N__44136));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_12_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_12_0  (
            .in0(N__25255),
            .in1(N__25201),
            .in2(_gnd_net_),
            .in3(N__25150),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44894),
            .ce(),
            .sr(N__25125));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26483),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_12_4  (
            .in0(N__26824),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26423),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26525),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__28709),
            .in2(N__25562),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__27124),
            .in2(_gnd_net_),
            .in3(N__25079),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(N__44888),
            .ce(),
            .sr(N__31409));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__26924),
            .in2(N__27101),
            .in3(N__25301),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(N__44888),
            .ce(),
            .sr(N__31409));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__27049),
            .in2(_gnd_net_),
            .in3(N__25298),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(N__44888),
            .ce(),
            .sr(N__31409));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__27025),
            .in2(_gnd_net_),
            .in3(N__25295),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(N__44888),
            .ce(),
            .sr(N__31409));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__27445),
            .in2(_gnd_net_),
            .in3(N__25292),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(N__44888),
            .ce(),
            .sr(N__31409));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__27403),
            .in2(_gnd_net_),
            .in3(N__25289),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(N__44888),
            .ce(),
            .sr(N__31409));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__27376),
            .in2(_gnd_net_),
            .in3(N__25286),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(N__44888),
            .ce(),
            .sr(N__31409));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__27325),
            .in2(_gnd_net_),
            .in3(N__25283),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(N__44882),
            .ce(),
            .sr(N__31408));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__27289),
            .in2(_gnd_net_),
            .in3(N__25280),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(N__44882),
            .ce(),
            .sr(N__31408));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__27262),
            .in2(_gnd_net_),
            .in3(N__25277),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(N__44882),
            .ce(),
            .sr(N__31408));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__27211),
            .in2(_gnd_net_),
            .in3(N__25325),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(N__44882),
            .ce(),
            .sr(N__31408));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__27187),
            .in2(_gnd_net_),
            .in3(N__25322),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(N__44882),
            .ce(),
            .sr(N__31408));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__27679),
            .in2(_gnd_net_),
            .in3(N__25319),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(N__44882),
            .ce(),
            .sr(N__31408));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__27628),
            .in2(_gnd_net_),
            .in3(N__25316),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(N__44882),
            .ce(),
            .sr(N__31408));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__27601),
            .in2(_gnd_net_),
            .in3(N__25313),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(N__44882),
            .ce(),
            .sr(N__31408));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__27562),
            .in2(_gnd_net_),
            .in3(N__25310),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(N__44875),
            .ce(),
            .sr(N__31400));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__27526),
            .in2(_gnd_net_),
            .in3(N__25307),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(N__44875),
            .ce(),
            .sr(N__31400));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__27478),
            .in2(_gnd_net_),
            .in3(N__25304),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44875),
            .ce(),
            .sr(N__31400));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_8_LC_11_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_8_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_8_LC_11_16_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_8_LC_11_16_1  (
            .in0(N__25788),
            .in1(N__25931),
            .in2(_gnd_net_),
            .in3(N__26076),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44868),
            .ce(N__31522),
            .sr(N__44168));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_11_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_11_16_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_11_16_2  (
            .in0(N__31855),
            .in1(N__26389),
            .in2(N__25547),
            .in3(N__25519),
            .lcout(elapsed_time_ns_1_RNID6DJ11_0_7),
            .ltout(elapsed_time_ns_1_RNID6DJ11_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_7_LC_11_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_7_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_7_LC_11_16_3 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_7_LC_11_16_3  (
            .in0(N__25787),
            .in1(_gnd_net_),
            .in2(N__25499),
            .in3(N__25932),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44868),
            .ce(N__31522),
            .sr(N__44168));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_11_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_11_16_4 .LUT_INIT=16'b1101111111001110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_11_16_4  (
            .in0(N__31856),
            .in1(N__31645),
            .in2(N__25496),
            .in3(N__25846),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_11_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_11_16_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25475),
            .in3(N__25468),
            .lcout(elapsed_time_ns_1_RNIDP2KD1_0_1),
            .ltout(elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_1_LC_11_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_1_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_1_LC_11_16_6 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_1_LC_11_16_6  (
            .in0(N__25929),
            .in1(N__25789),
            .in2(N__25418),
            .in3(N__25829),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44868),
            .ce(N__31522),
            .sr(N__44168));
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_2_LC_11_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_2_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_time_esr_2_LC_11_16_7 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_esr_2_LC_11_16_7  (
            .in0(N__25786),
            .in1(N__25930),
            .in2(N__25732),
            .in3(N__25402),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44868),
            .ce(N__31522),
            .sr(N__44168));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_6_LC_11_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_6_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_6_LC_11_17_0 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_6_LC_11_17_0  (
            .in0(N__25720),
            .in1(N__25935),
            .in2(N__31687),
            .in3(N__25797),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44862),
            .ce(N__25642),
            .sr(N__44176));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_2_LC_11_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_2_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_2_LC_11_17_1 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_2_LC_11_17_1  (
            .in0(N__25937),
            .in1(N__25790),
            .in2(N__25403),
            .in3(N__25721),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44862),
            .ce(N__25642),
            .sr(N__44176));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_4_LC_11_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_4_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_4_LC_11_17_2 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_4_LC_11_17_2  (
            .in0(N__25719),
            .in1(N__25934),
            .in2(N__25376),
            .in3(N__25796),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44862),
            .ce(N__25642),
            .sr(N__44176));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_5_LC_11_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_5_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_5_LC_11_17_3 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_5_LC_11_17_3  (
            .in0(N__25938),
            .in1(N__25715),
            .in2(N__26129),
            .in3(N__25791),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44862),
            .ce(N__25642),
            .sr(N__44176));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_8_LC_11_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_8_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_8_LC_11_17_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_8_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__25933),
            .in2(N__26078),
            .in3(N__25798),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44862),
            .ce(N__25642),
            .sr(N__44176));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_1_LC_11_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_1_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_1_LC_11_17_5 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_1_LC_11_17_5  (
            .in0(N__25936),
            .in1(N__25850),
            .in2(N__25804),
            .in3(N__25828),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44862),
            .ce(N__25642),
            .sr(N__44176));
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_3_LC_11_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_3_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_time_esr_3_LC_11_17_6 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_esr_3_LC_11_17_6  (
            .in0(N__26210),
            .in1(N__25792),
            .in2(N__25731),
            .in3(N__25672),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44862),
            .ce(N__25642),
            .sr(N__44176));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_17_7  (
            .in0(N__40218),
            .in1(N__38435),
            .in2(_gnd_net_),
            .in3(N__38402),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_18_1 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_18_1  (
            .in0(N__29066),
            .in1(N__29143),
            .in2(_gnd_net_),
            .in3(N__29097),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_433_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_11_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_11_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__28559),
            .in2(_gnd_net_),
            .in3(N__28578),
            .lcout(\phase_controller_inst1.stoper_tr.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_11_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_11_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__31458),
            .in2(_gnd_net_),
            .in3(N__28797),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26411),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_11_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_11_18_5 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_11_18_5  (
            .in0(N__26397),
            .in1(N__31857),
            .in2(N__26255),
            .in3(N__26224),
            .lcout(elapsed_time_ns_1_RNI81DJ11_0_2),
            .ltout(elapsed_time_ns_1_RNI81DJ11_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_o2_1_LC_11_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_o2_1_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_f0_0_o2_1_LC_11_18_6 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_f0_0_o2_1_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26213),
            .in3(N__26205),
            .lcout(\phase_controller_inst1.stoper_hc.N_283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26501),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_19_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__29413),
            .in2(_gnd_net_),
            .in3(N__28761),
            .lcout(),
            .ltout(\phase_controller_inst1.start_timer_tr_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_LC_11_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_11_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_11_19_2 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_11_19_2  (
            .in0(N__28579),
            .in1(N__26666),
            .in2(N__26165),
            .in3(N__26158),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44853),
            .ce(),
            .sr(N__44186));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__28732),
            .in2(_gnd_net_),
            .in3(N__26143),
            .lcout(\phase_controller_inst1.N_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_0_LC_11_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_11_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_11_19_4 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst1.state_0_LC_11_19_4  (
            .in0(N__29414),
            .in1(N__28762),
            .in2(N__26147),
            .in3(N__28733),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44853),
            .ce(),
            .sr(N__44186));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_11_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_11_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__28852),
            .in2(_gnd_net_),
            .in3(N__28890),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_20_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__28009),
            .in2(_gnd_net_),
            .in3(N__26444),
            .lcout(),
            .ltout(\phase_controller_inst2.start_timer_hc_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_LC_11_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_11_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_11_20_2 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_11_20_2  (
            .in0(N__32007),
            .in1(N__26459),
            .in2(N__26450),
            .in3(N__26663),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44849),
            .ce(),
            .sr(N__44200));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_20_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_20_4 .LUT_INIT=16'b1010101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_11_20_4  (
            .in0(N__26445),
            .in1(N__31985),
            .in2(N__28814),
            .in3(N__31472),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44849),
            .ce(),
            .sr(N__44200));
    defparam \phase_controller_inst2.state_1_LC_11_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_11_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_11_20_5 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst2.state_1_LC_11_20_5  (
            .in0(N__26623),
            .in1(N__28010),
            .in2(N__26592),
            .in3(N__26446),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44849),
            .ce(),
            .sr(N__44200));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_11_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_11_20_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__26580),
            .in2(_gnd_net_),
            .in3(N__26622),
            .lcout(),
            .ltout(\phase_controller_inst2.start_timer_tr_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_11_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_11_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_11_20_7 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_11_20_7  (
            .in0(N__26664),
            .in1(N__43759),
            .in2(N__26429),
            .in3(N__28036),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44849),
            .ce(),
            .sr(N__44200));
    defparam \current_shift_inst.control_input_0_LC_11_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_0_LC_11_21_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_0_LC_11_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_0_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__27728),
            .in2(N__39866),
            .in3(N__39864),
            .lcout(\current_shift_inst.control_inputZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\current_shift_inst.control_input_1_cry_0 ),
            .clk(N__44846),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_LC_11_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_1_LC_11_21_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_1_LC_11_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_1_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__27719),
            .in2(_gnd_net_),
            .in3(N__26426),
            .lcout(\current_shift_inst.control_inputZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_0 ),
            .carryout(\current_shift_inst.control_input_1_cry_1 ),
            .clk(N__44846),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_2_LC_11_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_2_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_2_LC_11_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_2_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(N__27710),
            .in2(_gnd_net_),
            .in3(N__26414),
            .lcout(\current_shift_inst.control_inputZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_1 ),
            .carryout(\current_shift_inst.control_input_1_cry_2 ),
            .clk(N__44846),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_3_LC_11_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_3_LC_11_21_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_3_LC_11_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_3_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__27821),
            .in2(_gnd_net_),
            .in3(N__26402),
            .lcout(\current_shift_inst.control_inputZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_2 ),
            .carryout(\current_shift_inst.control_input_1_cry_3 ),
            .clk(N__44846),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_4_LC_11_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_4_LC_11_21_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_4_LC_11_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_4_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__27812),
            .in2(_gnd_net_),
            .in3(N__26510),
            .lcout(\current_shift_inst.control_inputZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_3 ),
            .carryout(\current_shift_inst.control_input_1_cry_4 ),
            .clk(N__44846),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_5_LC_11_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_5_LC_11_21_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_5_LC_11_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_5_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(N__27803),
            .in2(_gnd_net_),
            .in3(N__26507),
            .lcout(\current_shift_inst.control_inputZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_4 ),
            .carryout(\current_shift_inst.control_input_1_cry_5 ),
            .clk(N__44846),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_6_LC_11_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_6_LC_11_21_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_6_LC_11_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_6_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__27794),
            .in2(_gnd_net_),
            .in3(N__26504),
            .lcout(\current_shift_inst.control_inputZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_5 ),
            .carryout(\current_shift_inst.control_input_1_cry_6 ),
            .clk(N__44846),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_7_LC_11_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_7_LC_11_21_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_7_LC_11_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_7_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__27773),
            .in2(_gnd_net_),
            .in3(N__26492),
            .lcout(\current_shift_inst.control_inputZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_6 ),
            .carryout(\current_shift_inst.control_input_1_cry_7 ),
            .clk(N__44846),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_8_LC_11_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_8_LC_11_22_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_8_LC_11_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_8_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__27764),
            .in2(_gnd_net_),
            .in3(N__26489),
            .lcout(\current_shift_inst.control_inputZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\current_shift_inst.control_input_1_cry_8 ),
            .clk(N__44843),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_9_LC_11_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_9_LC_11_22_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_9_LC_11_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_9_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__27755),
            .in2(_gnd_net_),
            .in3(N__26486),
            .lcout(\current_shift_inst.control_inputZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_8 ),
            .carryout(\current_shift_inst.control_input_1_cry_9 ),
            .clk(N__44843),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_10_LC_11_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_10_LC_11_22_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_10_LC_11_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_10_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__26465),
            .in2(_gnd_net_),
            .in3(N__26471),
            .lcout(\current_shift_inst.control_inputZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_9 ),
            .carryout(\current_shift_inst.control_input_1_cry_10 ),
            .clk(N__44843),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_11_LC_11_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_11_LC_11_22_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_11_LC_11_22_3 .LUT_INIT=16'b0001110111100010;
    LogicCell40 \current_shift_inst.control_input_11_LC_11_22_3  (
            .in0(N__40125),
            .in1(N__28046),
            .in2(N__27743),
            .in3(N__26468),
            .lcout(\current_shift_inst.control_inputZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44843),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_c_RNIG7KU_LC_11_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_c_RNIG7KU_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_c_RNIG7KU_LC_11_22_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_c_RNIG7KU_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__28045),
            .in2(_gnd_net_),
            .in3(N__27739),
            .lcout(\current_shift_inst.control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26729),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_4_LC_11_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_11_23_3 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_11_23_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_11_23_3  (
            .in0(N__26700),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26651),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44841),
            .ce(),
            .sr(N__44222));
    defparam \phase_controller_inst2.state_0_LC_11_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_11_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_11_23_5 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \phase_controller_inst2.state_0_LC_11_23_5  (
            .in0(N__26627),
            .in1(N__40814),
            .in2(N__27938),
            .in3(N__26591),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44841),
            .ce(),
            .sr(N__44222));
    defparam \phase_controller_inst2.T23_LC_11_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.T23_LC_11_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T23_LC_11_24_7 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst2.T23_LC_11_24_7  (
            .in0(N__26536),
            .in1(N__26602),
            .in2(_gnd_net_),
            .in3(N__27936),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44839),
            .ce(),
            .sr(N__44227));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_12_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_12_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31253),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_12_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_12_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30808),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_12_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_12_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31002),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_12_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_12_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30529),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_12_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_12_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34875),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_12_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_12_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_12_8_4  (
            .in0(N__35038),
            .in1(N__35099),
            .in2(N__34588),
            .in3(N__28661),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_12_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_12_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_12_8_5  (
            .in0(N__26741),
            .in1(N__30263),
            .in2(N__26744),
            .in3(N__28178),
            .lcout(\current_shift_inst.PI_CTRL.N_74_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_12_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_12_8_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_12_8_6  (
            .in0(N__32508),
            .in1(N__35166),
            .in2(N__32557),
            .in3(N__34342),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_8_7  (
            .in0(N__34874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31341),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_12_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_12_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32246),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_12_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_12_9_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_12_9_3  (
            .in0(N__34882),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_12_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_12_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_12_9_4  (
            .in0(N__30840),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34881),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_12_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_12_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_12_9_5  (
            .in0(N__30703),
            .in1(N__32612),
            .in2(N__31009),
            .in3(N__30382),
            .lcout(\current_shift_inst.PI_CTRL.N_74_16 ),
            .ltout(\current_shift_inst.PI_CTRL.N_74_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_12_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_12_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_12_9_6  (
            .in0(N__28147),
            .in1(N__28165),
            .in2(N__26732),
            .in3(N__34228),
            .lcout(\current_shift_inst.PI_CTRL.N_103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_12_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_12_10_0 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_12_10_0  (
            .in0(N__32338),
            .in1(N__34890),
            .in2(N__28352),
            .in3(N__26902),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_12_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_12_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34486),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34437),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_12_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_12_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32337),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26901),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_12_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_12_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34223),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__26777),
            .in2(_gnd_net_),
            .in3(N__26801),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__26933),
            .in2(_gnd_net_),
            .in3(N__26771),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__44893),
            .ce(),
            .sr(N__44130));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__26768),
            .in2(_gnd_net_),
            .in3(N__26762),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__44893),
            .ce(),
            .sr(N__44130));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__26759),
            .in2(_gnd_net_),
            .in3(N__26747),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__44893),
            .ce(),
            .sr(N__44130));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__26918),
            .in2(_gnd_net_),
            .in3(N__26912),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__44893),
            .ce(),
            .sr(N__44130));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__38327),
            .in2(_gnd_net_),
            .in3(N__26888),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__44893),
            .ce(),
            .sr(N__44130));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__26975),
            .in2(_gnd_net_),
            .in3(N__26885),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__44893),
            .ce(),
            .sr(N__44130));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__26882),
            .in2(_gnd_net_),
            .in3(N__26870),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__44893),
            .ce(),
            .sr(N__44130));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__26951),
            .in2(_gnd_net_),
            .in3(N__26867),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__44887),
            .ce(),
            .sr(N__44137));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__26864),
            .in2(_gnd_net_),
            .in3(N__26849),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__44887),
            .ce(),
            .sr(N__44137));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__26846),
            .in2(_gnd_net_),
            .in3(N__26840),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__44887),
            .ce(),
            .sr(N__44137));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__26837),
            .in2(_gnd_net_),
            .in3(N__26831),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__44887),
            .ce(),
            .sr(N__44137));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__26828),
            .in2(_gnd_net_),
            .in3(N__26804),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44887),
            .ce(),
            .sr(N__44137));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_13_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_13_0  (
            .in0(N__41880),
            .in1(N__43190),
            .in2(_gnd_net_),
            .in3(N__43148),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44880),
            .ce(),
            .sr(N__39651));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26990),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26966),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30330),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31212),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26945),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHE_LC_12_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHE_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHE_LC_12_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHE_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__31470),
            .in2(_gnd_net_),
            .in3(N__28809),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIIGHEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_12_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_12_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_12_14_2  (
            .in0(N__31303),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34864),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_12_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_12_14_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_12_14_3  (
            .in0(N__34867),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31141),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_12_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_12_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_12_14_4  (
            .in0(N__30594),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34865),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_12_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_12_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_12_14_5  (
            .in0(N__34866),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33268),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_12_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_12_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__33526),
            .in2(_gnd_net_),
            .in3(N__34868),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_12_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_12_15_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_12_15_0  (
            .in0(N__28701),
            .in1(N__27149),
            .in2(N__27143),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_12_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_12_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__27110),
            .in2(N__27134),
            .in3(N__27125),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_12_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_12_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_12_15_2  (
            .in0(N__27100),
            .in1(N__27068),
            .in2(N__27083),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_12_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_12_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__27062),
            .in2(N__27035),
            .in3(N__27050),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_12_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_12_15_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_12_15_4  (
            .in0(N__27026),
            .in1(N__27011),
            .in2(N__26999),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_12_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_12_15_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_12_15_5  (
            .in0(N__27449),
            .in1(N__27431),
            .in2(N__27419),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_12_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_12_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__27410),
            .in2(N__27389),
            .in3(N__27404),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_12_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_12_15_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_12_15_7  (
            .in0(N__27377),
            .in1(N__27362),
            .in2(N__27356),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_12_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_12_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__27344),
            .in2(N__27311),
            .in3(N__27332),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_12_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_12_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__27302),
            .in2(N__27275),
            .in3(N__27290),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_12_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_12_16_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_12_16_2  (
            .in0(N__27266),
            .in1(N__27248),
            .in2(N__27236),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_12_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_12_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__27227),
            .in2(N__27197),
            .in3(N__27212),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_12_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_12_16_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_12_16_4  (
            .in0(N__27188),
            .in1(N__27173),
            .in2(N__27158),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_12_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_12_16_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_12_16_5  (
            .in0(N__27680),
            .in1(N__27665),
            .in2(N__27653),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_12_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_12_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__27641),
            .in2(N__27614),
            .in3(N__27629),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_12_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_12_16_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_12_16_7  (
            .in0(N__27602),
            .in1(N__27587),
            .in2(N__27575),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_12_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_12_17_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_12_17_0  (
            .in0(N__27563),
            .in1(N__27548),
            .in2(N__27536),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_12_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_12_17_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_12_17_1  (
            .in0(N__27527),
            .in1(N__27512),
            .in2(N__27500),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_12_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_12_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__27491),
            .in2(N__27464),
            .in3(N__27479),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_12_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_12_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27452),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_c_RNO_LC_12_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_c_RNO_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_c_RNO_LC_12_17_4 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_c_RNO_LC_12_17_4  (
            .in0(N__37976),
            .in1(N__37949),
            .in2(_gnd_net_),
            .in3(N__40184),
            .lcout(\current_shift_inst.un38_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_c_RNO_LC_12_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_c_RNO_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_c_RNO_LC_12_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_c_RNO_LC_12_17_5  (
            .in0(N__40183),
            .in1(N__37259),
            .in2(_gnd_net_),
            .in3(N__37232),
            .lcout(\current_shift_inst.un38_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_c_RNO_LC_12_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_c_RNO_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_c_RNO_LC_12_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_c_RNO_LC_12_17_7  (
            .in0(N__40182),
            .in1(N__37300),
            .in2(_gnd_net_),
            .in3(N__37274),
            .lcout(\current_shift_inst.un38_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_c_THRU_CRY_0_LC_12_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_c_THRU_CRY_0_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_c_THRU_CRY_0_LC_12_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_c_THRU_CRY_0_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__40143),
            .in2(N__40269),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_c_LC_12_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_c_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_c_LC_12_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_c_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__31907),
            .in2(N__39865),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.un38_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_c_LC_12_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_c_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_c_LC_12_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_c_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__29150),
            .in2(N__40270),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_c_LC_12_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_c_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_c_LC_12_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_c_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__32069),
            .in2(N__40219),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_c_LC_12_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_c_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_c_LC_12_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_c_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__27692),
            .in2(N__40271),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_c_LC_12_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_c_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_c_LC_12_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_c_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__27686),
            .in2(N__40220),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_c_LC_12_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_c_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_c_LC_12_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_c_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__32144),
            .in2(N__40272),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_c_LC_12_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_c_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_c_LC_12_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_c_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__31895),
            .in2(N__40221),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_c_LC_12_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_c_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_c_LC_12_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_c_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__27701),
            .in2(N__40222),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_c_LC_12_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_c_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_c_LC_12_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_c_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__40156),
            .in2(N__32126),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_7 ),
            .carryout(\current_shift_inst.un38_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_c_LC_12_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_c_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_c_LC_12_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_c_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__31883),
            .in2(N__40223),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_c_LC_12_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_c_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_c_LC_12_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_c_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__40160),
            .in2(N__32111),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_c_LC_12_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_c_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_c_LC_12_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_c_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__37424),
            .in2(N__40224),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_c_LC_12_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_c_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_c_LC_12_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_c_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__40164),
            .in2(N__32096),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_c_LC_12_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_c_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_c_LC_12_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_c_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__32135),
            .in2(N__40225),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_c_LC_12_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_c_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_c_LC_12_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_c_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(N__40168),
            .in2(N__37991),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_c_LC_12_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_c_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_c_LC_12_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_c_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__32081),
            .in2(N__40273),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_c_LC_12_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_c_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_c_LC_12_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_c_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__38444),
            .in2(N__40226),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_15 ),
            .carryout(\current_shift_inst.un38_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_c_LC_12_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_c_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_c_LC_12_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_c_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__38045),
            .in2(N__40274),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_c_LC_12_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_c_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_c_LC_12_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_c_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__40248),
            .in2(N__38699),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_c_LC_12_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_c_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_c_LC_12_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_c_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__28622),
            .in2(N__40275),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_c_RNIBS3R1_LC_12_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_c_RNIBS3R1_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_c_RNIBS3R1_LC_12_20_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_c_RNIBS3R1_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(N__38759),
            .in2(N__40227),
            .in3(N__27722),
            .lcout(\current_shift_inst.control_input_1_axb_0 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_c_RNITVMS1_LC_12_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_c_RNITVMS1_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_c_RNITVMS1_LC_12_20_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_c_RNITVMS1_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__38222),
            .in2(N__40276),
            .in3(N__27713),
            .lcout(\current_shift_inst.control_input_1_axb_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_c_RNI16PS1_LC_12_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_c_RNI16PS1_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_c_RNI16PS1_LC_12_20_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_c_RNI16PS1_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(N__40255),
            .in2(N__32159),
            .in3(N__27704),
            .lcout(\current_shift_inst.control_input_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_c_RNI5CRS1_LC_12_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_c_RNI5CRS1_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_c_RNI5CRS1_LC_12_21_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_c_RNI5CRS1_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__38852),
            .in2(N__40277),
            .in3(N__27815),
            .lcout(\current_shift_inst.control_input_1_axb_3 ),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_c_RNI9ITS1_LC_12_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_c_RNI9ITS1_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_c_RNI9ITS1_LC_12_21_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_c_RNI9ITS1_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(N__34127),
            .in2(N__40228),
            .in3(N__27806),
            .lcout(\current_shift_inst.control_input_1_axb_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_23 ),
            .carryout(\current_shift_inst.un38_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_c_RNIDOVS1_LC_12_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_c_RNIDOVS1_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_c_RNIDOVS1_LC_12_21_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_c_RNIDOVS1_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(N__34154),
            .in2(N__40278),
            .in3(N__27797),
            .lcout(\current_shift_inst.control_input_1_axb_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_c_RNIHU1T1_LC_12_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_c_RNIHU1T1_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_c_RNIHU1T1_LC_12_21_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_c_RNIHU1T1_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(N__34136),
            .in2(N__40229),
            .in3(N__27788),
            .lcout(\current_shift_inst.control_input_1_axb_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_c_RNIL44T1_LC_12_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_c_RNIL44T1_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_c_RNIL44T1_LC_12_21_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_c_RNIL44T1_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(N__27785),
            .in2(N__40279),
            .in3(N__27767),
            .lcout(\current_shift_inst.control_input_1_axb_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_c_RNIPA6T1_LC_12_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_c_RNIPA6T1_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_c_RNIPA6T1_LC_12_21_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_c_RNIPA6T1_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__40265),
            .in2(N__32192),
            .in3(N__27758),
            .lcout(\current_shift_inst.control_input_1_axb_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_c_RNIB0AT1_LC_12_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_c_RNIB0AT1_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_c_RNIB0AT1_LC_12_21_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_c_RNIB0AT1_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__34145),
            .in2(N__40280),
            .in3(N__27749),
            .lcout(\current_shift_inst.control_input_1_axb_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_THRU_LUT4_0_LC_12_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_THRU_LUT4_0_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_THRU_LUT4_0_LC_12_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_THRU_LUT4_0_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27746),
            .lcout(\current_shift_inst.un38_control_input_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_12_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_12_22_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_12_22_4  (
            .in0(N__40181),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34007),
            .lcout(\current_shift_inst.un38_control_input_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_12_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_12_22_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(N__40813),
            .in2(_gnd_net_),
            .in3(N__27929),
            .lcout(\phase_controller_inst2.time_passed_RNI9M3O ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.T01_LC_12_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.T01_LC_12_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T01_LC_12_23_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst2.T01_LC_12_23_3  (
            .in0(N__27973),
            .in1(N__27906),
            .in2(_gnd_net_),
            .in3(N__28019),
            .lcout(T01_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44838),
            .ce(),
            .sr(N__44215));
    defparam \phase_controller_inst1.S1_LC_12_25_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_12_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_12_25_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.S1_LC_12_25_1  (
            .in0(N__28858),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44834),
            .ce(),
            .sr(N__44228));
    defparam \current_shift_inst.stop_timer_s1_LC_12_25_2 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_12_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_12_25_2 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_12_25_2  (
            .in0(N__27952),
            .in1(N__28857),
            .in2(N__28094),
            .in3(N__28129),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44834),
            .ce(),
            .sr(N__44228));
    defparam \current_shift_inst.timer_s1.running_LC_12_25_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_12_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_12_25_3 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_12_25_3  (
            .in0(N__28130),
            .in1(N__28090),
            .in2(_gnd_net_),
            .in3(N__28112),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44834),
            .ce(),
            .sr(N__44228));
    defparam \current_shift_inst.start_timer_s1_LC_12_25_4 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_12_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_12_25_4 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_12_25_4  (
            .in0(N__27951),
            .in1(N__28128),
            .in2(_gnd_net_),
            .in3(N__28856),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44834),
            .ce(),
            .sr(N__44228));
    defparam \phase_controller_inst2.T45_LC_12_25_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.T45_LC_12_25_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T45_LC_12_25_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \phase_controller_inst2.T45_LC_12_25_7  (
            .in0(N__27937),
            .in1(N__27844),
            .in2(_gnd_net_),
            .in3(N__27908),
            .lcout(T45_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44834),
            .ce(),
            .sr(N__44228));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_12_26_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_12_26_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_12_26_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_12_26_3  (
            .in0(_gnd_net_),
            .in1(N__28109),
            .in2(_gnd_net_),
            .in3(N__28088),
            .lcout(\current_shift_inst.timer_s1.N_166_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_12_26_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_12_26_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_12_26_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_12_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28110),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_26_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_26_7 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_26_7  (
            .in0(N__28127),
            .in1(N__28111),
            .in2(_gnd_net_),
            .in3(N__28089),
            .lcout(\current_shift_inst.timer_s1.N_167_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_6 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_6 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_6  (
            .in0(N__44334),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_13_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_13_6_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_13_6_4 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_13_6_4  (
            .in0(N__35629),
            .in1(N__35828),
            .in2(N__32723),
            .in3(N__35462),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44922),
            .ce(),
            .sr(N__44112));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_13_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_13_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31059),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_13_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_13_6_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_13_6_7 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_13_6_7  (
            .in0(N__35827),
            .in1(N__35630),
            .in2(N__35507),
            .in3(N__33380),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44922),
            .ce(),
            .sr(N__44112));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_13_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_13_7_0 .LUT_INIT=16'b0011001100110111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_13_7_0  (
            .in0(N__34485),
            .in1(N__32245),
            .in2(N__32336),
            .in3(N__32407),
            .lcout(\current_shift_inst.PI_CTRL.N_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_13_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_13_7_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_13_7_1  (
            .in0(N__28640),
            .in1(N__28172),
            .in2(N__35877),
            .in3(N__34283),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_13_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_13_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_13_7_2  (
            .in0(N__28208),
            .in1(N__28214),
            .in2(N__28058),
            .in3(N__28184),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_13_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_13_7_3 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_13_7_3  (
            .in0(N__30287),
            .in1(N__28055),
            .in2(N__28049),
            .in3(N__28190),
            .lcout(\current_shift_inst.PI_CTRL.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_13_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_13_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30286),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_13_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_13_7_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_13_7_5  (
            .in0(N__31241),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30630),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_13_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_13_7_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_13_7_6  (
            .in0(N__30421),
            .in1(N__31085),
            .in2(N__28193),
            .in3(N__34645),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_13_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_13_8_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_13_8_0  (
            .in0(N__34227),
            .in1(N__32507),
            .in2(_gnd_net_),
            .in3(N__28202),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_13_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_13_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_13_8_1  (
            .in0(N__30791),
            .in1(N__35321),
            .in2(N__34527),
            .in3(N__35207),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_13_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_13_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_13_8_2  (
            .in0(N__35156),
            .in1(N__32549),
            .in2(N__35042),
            .in3(N__34340),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_13_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_13_8_3 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_13_8_3  (
            .in0(N__28166),
            .in1(N__28154),
            .in2(N__34172),
            .in3(N__28136),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_13_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_13_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_13_8_4  (
            .in0(N__30463),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34873),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_13_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_13_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30422),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_13_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_13_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_13_8_6  (
            .in0(N__35206),
            .in1(N__30790),
            .in2(N__35328),
            .in3(N__34517),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_13_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_13_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_13_8_7  (
            .in0(N__34381),
            .in1(N__35810),
            .in2(N__30524),
            .in3(N__30893),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_13_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_13_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_13_9_0  (
            .in0(N__30685),
            .in1(N__30994),
            .in2(N__32617),
            .in3(N__30367),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_13_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_13_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_13_9_1  (
            .in0(N__28519),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34877),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_13_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_13_9_2 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_13_9_2  (
            .in0(N__34879),
            .in1(N__30368),
            .in2(N__28196),
            .in3(N__28505),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_13_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_13_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30686),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_13_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_13_9_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_13_9_4  (
            .in0(N__35100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_9_5  (
            .in0(N__30558),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34876),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_13_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_13_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_13_9_6  (
            .in0(N__34878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30739),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_13_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_13_9_7 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_13_9_7  (
            .in0(N__31187),
            .in1(N__32556),
            .in2(N__28478),
            .in3(N__34880),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_13_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_13_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__30967),
            .in2(_gnd_net_),
            .in3(N__34884),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_13_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_13_10_1 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_13_10_1  (
            .in0(N__28291),
            .in1(N__32251),
            .in2(N__34943),
            .in3(N__28325),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28290),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_13_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_13_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__30769),
            .in2(_gnd_net_),
            .in3(N__34885),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_13_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_13_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28269),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_13_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_13_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_13_10_6  (
            .in0(N__30928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34883),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_13_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_13_10_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_13_10_7  (
            .in0(N__34886),
            .in1(N__32443),
            .in2(N__28370),
            .in3(N__28270),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_13_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_13_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__28238),
            .in2(_gnd_net_),
            .in3(N__28252),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_13_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_13_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__28220),
            .in2(_gnd_net_),
            .in3(N__28231),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_13_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_13_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__28406),
            .in2(_gnd_net_),
            .in3(N__28423),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_13_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_13_11_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_13_11_3  (
            .in0(N__28393),
            .in1(N__28382),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_13_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_13_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__28376),
            .in2(_gnd_net_),
            .in3(N__28361),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_13_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_13_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__28358),
            .in2(_gnd_net_),
            .in3(N__28343),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_13_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_13_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__28340),
            .in2(_gnd_net_),
            .in3(N__28334),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_13_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_13_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__28331),
            .in2(_gnd_net_),
            .in3(N__28319),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_13_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_13_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__28316),
            .in2(_gnd_net_),
            .in3(N__28310),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_8 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_13_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_13_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__28307),
            .in2(_gnd_net_),
            .in3(N__28301),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_13_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_13_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__28685),
            .in2(_gnd_net_),
            .in3(N__28454),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_13_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_13_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__28676),
            .in2(_gnd_net_),
            .in3(N__28451),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_13_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_13_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__30464),
            .in2(_gnd_net_),
            .in3(N__28448),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_13_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_13_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__31111),
            .in2(_gnd_net_),
            .in3(N__28445),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_13_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_13_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__31033),
            .in2(_gnd_net_),
            .in3(N__28442),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_13_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_13_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__31348),
            .in2(_gnd_net_),
            .in3(N__28439),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_13_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_13_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__30559),
            .in2(_gnd_net_),
            .in3(N__28436),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_13_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_13_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__30929),
            .in2(_gnd_net_),
            .in3(N__28433),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_13_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_13_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__30847),
            .in2(_gnd_net_),
            .in3(N__28430),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_13_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_13_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__28520),
            .in2(_gnd_net_),
            .in3(N__28496),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_13_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_13_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(N__30770),
            .in2(_gnd_net_),
            .in3(N__28493),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_13_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_13_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(N__30968),
            .in2(_gnd_net_),
            .in3(N__28490),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_13_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_13_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__31936),
            .in2(_gnd_net_),
            .in3(N__28487),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_13_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_13_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(N__30740),
            .in2(_gnd_net_),
            .in3(N__28484),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_13_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_13_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(N__31293),
            .in2(_gnd_net_),
            .in3(N__28481),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ),
            .ltout(),
            .carryin(bfn_13_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_13_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_13_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__31186),
            .in2(_gnd_net_),
            .in3(N__28463),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_13_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_13_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30595),
            .in3(N__28460),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_13_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_13_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__33264),
            .in2(_gnd_net_),
            .in3(N__28457),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_13_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_13_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__31137),
            .in2(_gnd_net_),
            .in3(N__28610),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_13_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_13_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(N__33516),
            .in2(_gnd_net_),
            .in3(N__28607),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_13_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_13_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(N__31957),
            .in2(_gnd_net_),
            .in3(N__28604),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_13_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_13_14_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_13_14_7  (
            .in0(N__34833),
            .in1(N__28663),
            .in2(_gnd_net_),
            .in3(N__28601),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIL7IU_0_1_LC_13_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIL7IU_0_1_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIL7IU_0_1_LC_13_15_0 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIL7IU_0_1_LC_13_15_0  (
            .in0(N__28553),
            .in1(N__44318),
            .in2(N__28597),
            .in3(N__43178),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_15_1 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_15_1  (
            .in0(N__43179),
            .in1(N__28596),
            .in2(N__43143),
            .in3(N__28554),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44876),
            .ce(),
            .sr(N__44150));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_15_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__43174),
            .in2(_gnd_net_),
            .in3(N__43132),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_13_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_13_15_4 .LUT_INIT=16'b0010000001100100;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_13_15_4  (
            .in0(N__28555),
            .in1(N__43181),
            .in2(N__28598),
            .in3(N__43139),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44876),
            .ce(),
            .sr(N__44150));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIL7IU_1_LC_13_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIL7IU_1_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIL7IU_1_LC_13_15_5 .LUT_INIT=16'b1010101110101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIL7IU_1_LC_13_15_5  (
            .in0(N__44319),
            .in1(N__28589),
            .in2(N__43188),
            .in3(N__28552),
            .lcout(\phase_controller_inst1.stoper_tr.un1_stoper_state12_1_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_7 .LUT_INIT=16'b1110111000000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_7  (
            .in0(N__43180),
            .in1(N__28532),
            .in2(N__43144),
            .in3(N__28725),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44876),
            .ce(),
            .sr(N__44150));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_13_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_13_16_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_13_16_0  (
            .in0(N__31462),
            .in1(N__28705),
            .in2(_gnd_net_),
            .in3(N__28808),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44869),
            .ce(),
            .sr(N__31407));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_13_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_13_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34993),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_13_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30249),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35878),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_13_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30908),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_13_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_13_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28662),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_13_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34584),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_c_RNO_LC_13_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_c_RNO_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_c_RNO_LC_13_17_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_c_RNO_LC_13_17_0  (
            .in0(N__40115),
            .in1(_gnd_net_),
            .in2(N__38123),
            .in3(N__38093),
            .lcout(\current_shift_inst.un38_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38118),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_c_RNO_LC_13_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_c_RNO_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_c_RNO_LC_13_17_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_c_RNO_LC_13_17_2  (
            .in0(N__40114),
            .in1(N__33755),
            .in2(_gnd_net_),
            .in3(N__33806),
            .lcout(\current_shift_inst.un38_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_13_17_4 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_13_17_4  (
            .in0(N__29055),
            .in1(N__29144),
            .in2(_gnd_net_),
            .in3(N__29108),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44863),
            .ce(),
            .sr(N__44160));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_17_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_17_6  (
            .in0(N__29054),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_13_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_13_17_7 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_13_17_7  (
            .in0(N__36017),
            .in1(N__36553),
            .in2(N__37180),
            .in3(N__36182),
            .lcout(elapsed_time_ns_1_RNIAE2591_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_2_LC_13_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_13_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_13_18_1 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst1.state_2_LC_13_18_1  (
            .in0(N__28894),
            .in1(N__36588),
            .in2(N__36632),
            .in3(N__28859),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44858),
            .ce(),
            .sr(N__44169));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_13_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_13_18_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_0_LC_13_18_3  (
            .in0(N__32023),
            .in1(N__32050),
            .in2(N__28813),
            .in3(N__31457),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44858),
            .ce(),
            .sr(N__44169));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_13_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_13_18_4 .LUT_INIT=16'b0101001000000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_1_LC_13_18_4  (
            .in0(N__31456),
            .in1(N__28804),
            .in2(N__32057),
            .in3(N__32024),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44858),
            .ce(),
            .sr(N__44169));
    defparam \phase_controller_inst1.state_1_LC_13_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_13_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_13_18_5 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_inst1.state_1_LC_13_18_5  (
            .in0(N__29403),
            .in1(N__36589),
            .in2(N__28769),
            .in3(N__36630),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44858),
            .ce(),
            .sr(N__44169));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__29368),
            .in2(N__33649),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__44854),
            .ce(N__38178),
            .sr(N__44177));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__29343),
            .in2(N__33841),
            .in3(N__29177),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__44854),
            .ce(N__38178),
            .sr(N__44177));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__29369),
            .in2(N__29321),
            .in3(N__29174),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__44854),
            .ce(N__38178),
            .sr(N__44177));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__29287),
            .in2(N__29348),
            .in3(N__29171),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__44854),
            .ce(N__38178),
            .sr(N__44177));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__29320),
            .in2(N__29260),
            .in3(N__29168),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__44854),
            .ce(N__38178),
            .sr(N__44177));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__29644),
            .in2(N__29291),
            .in3(N__29165),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__44854),
            .ce(N__38178),
            .sr(N__44177));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__29614),
            .in2(N__29261),
            .in3(N__29162),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__44854),
            .ce(N__38178),
            .sr(N__44177));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__29645),
            .in2(N__29584),
            .in3(N__29159),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__44854),
            .ce(N__38178),
            .sr(N__44177));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__29551),
            .in2(N__29621),
            .in3(N__29156),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__44850),
            .ce(N__38177),
            .sr(N__44180));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__29527),
            .in2(N__29588),
            .in3(N__29153),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__44850),
            .ce(N__38177),
            .sr(N__44180));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(N__29552),
            .in2(N__29506),
            .in3(N__29204),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__44850),
            .ce(N__38177),
            .sr(N__44180));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__29528),
            .in2(N__29476),
            .in3(N__29201),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__44850),
            .ce(N__38177),
            .sr(N__44180));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__29443),
            .in2(N__29507),
            .in3(N__29198),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__44850),
            .ce(N__38177),
            .sr(N__44180));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__29899),
            .in2(N__29477),
            .in3(N__29195),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__44850),
            .ce(N__38177),
            .sr(N__44180));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(N__29872),
            .in2(N__29447),
            .in3(N__29192),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__44850),
            .ce(N__38177),
            .sr(N__44180));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__29900),
            .in2(N__29842),
            .in3(N__29189),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__44850),
            .ce(N__38177),
            .sr(N__44180));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__29806),
            .in2(N__29876),
            .in3(N__29186),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__44847),
            .ce(N__38176),
            .sr(N__44187));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__29782),
            .in2(N__29843),
            .in3(N__29183),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__44847),
            .ce(N__38176),
            .sr(N__44187));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__29807),
            .in2(N__29761),
            .in3(N__29180),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__44847),
            .ce(N__38176),
            .sr(N__44187));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(N__29783),
            .in2(N__29731),
            .in3(N__29231),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__44847),
            .ce(N__38176),
            .sr(N__44187));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(N__29698),
            .in2(N__29762),
            .in3(N__29228),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__44847),
            .ce(N__38176),
            .sr(N__44187));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__29671),
            .in2(N__29732),
            .in3(N__29225),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__44847),
            .ce(N__38176),
            .sr(N__44187));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(N__30202),
            .in2(N__29702),
            .in3(N__29222),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__44847),
            .ce(N__38176),
            .sr(N__44187));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(N__30175),
            .in2(N__29675),
            .in3(N__29219),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__44847),
            .ce(N__38176),
            .sr(N__44187));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__30148),
            .in2(N__30206),
            .in3(N__29216),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__44844),
            .ce(N__38175),
            .sr(N__44201));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__30124),
            .in2(N__30179),
            .in3(N__29213),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__44844),
            .ce(N__38175),
            .sr(N__44201));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__30149),
            .in2(N__30104),
            .in3(N__29210),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__44844),
            .ce(N__38175),
            .sr(N__44201));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(N__30125),
            .in2(N__29957),
            .in3(N__29207),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__44844),
            .ce(N__38175),
            .sr(N__44201));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29417),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_13_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29412),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44842),
            .ce(),
            .sr(N__44209));
    defparam \current_shift_inst.timer_s1.counter_0_LC_13_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_13_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_13_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_13_24_0  (
            .in0(N__30073),
            .in1(N__33633),
            .in2(_gnd_net_),
            .in3(N__29375),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__44840),
            .ce(N__29936),
            .sr(N__44216));
    defparam \current_shift_inst.timer_s1.counter_1_LC_13_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_13_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_13_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_13_24_1  (
            .in0(N__30069),
            .in1(N__33825),
            .in2(_gnd_net_),
            .in3(N__29372),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__44840),
            .ce(N__29936),
            .sr(N__44216));
    defparam \current_shift_inst.timer_s1.counter_2_LC_13_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_13_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_13_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_13_24_2  (
            .in0(N__30074),
            .in1(N__29367),
            .in2(_gnd_net_),
            .in3(N__29351),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__44840),
            .ce(N__29936),
            .sr(N__44216));
    defparam \current_shift_inst.timer_s1.counter_3_LC_13_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_13_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_13_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_13_24_3  (
            .in0(N__30070),
            .in1(N__29347),
            .in2(_gnd_net_),
            .in3(N__29324),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__44840),
            .ce(N__29936),
            .sr(N__44216));
    defparam \current_shift_inst.timer_s1.counter_4_LC_13_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_13_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_13_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_13_24_4  (
            .in0(N__30075),
            .in1(N__29310),
            .in2(_gnd_net_),
            .in3(N__29294),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__44840),
            .ce(N__29936),
            .sr(N__44216));
    defparam \current_shift_inst.timer_s1.counter_5_LC_13_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_13_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_13_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_13_24_5  (
            .in0(N__30071),
            .in1(N__29280),
            .in2(_gnd_net_),
            .in3(N__29264),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__44840),
            .ce(N__29936),
            .sr(N__44216));
    defparam \current_shift_inst.timer_s1.counter_6_LC_13_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_13_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_13_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_13_24_6  (
            .in0(N__30076),
            .in1(N__29248),
            .in2(_gnd_net_),
            .in3(N__29234),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__44840),
            .ce(N__29936),
            .sr(N__44216));
    defparam \current_shift_inst.timer_s1.counter_7_LC_13_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_13_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_13_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_13_24_7  (
            .in0(N__30072),
            .in1(N__29638),
            .in2(_gnd_net_),
            .in3(N__29624),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__44840),
            .ce(N__29936),
            .sr(N__44216));
    defparam \current_shift_inst.timer_s1.counter_8_LC_13_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_13_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_13_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_13_25_0  (
            .in0(N__30049),
            .in1(N__29613),
            .in2(_gnd_net_),
            .in3(N__29591),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__44837),
            .ce(N__29931),
            .sr(N__44223));
    defparam \current_shift_inst.timer_s1.counter_9_LC_13_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_13_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_13_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_13_25_1  (
            .in0(N__30053),
            .in1(N__29577),
            .in2(_gnd_net_),
            .in3(N__29555),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__44837),
            .ce(N__29931),
            .sr(N__44223));
    defparam \current_shift_inst.timer_s1.counter_10_LC_13_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_13_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_13_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_13_25_2  (
            .in0(N__30046),
            .in1(N__29545),
            .in2(_gnd_net_),
            .in3(N__29531),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__44837),
            .ce(N__29931),
            .sr(N__44223));
    defparam \current_shift_inst.timer_s1.counter_11_LC_13_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_13_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_13_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_13_25_3  (
            .in0(N__30050),
            .in1(N__29526),
            .in2(_gnd_net_),
            .in3(N__29510),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__44837),
            .ce(N__29931),
            .sr(N__44223));
    defparam \current_shift_inst.timer_s1.counter_12_LC_13_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_13_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_13_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_13_25_4  (
            .in0(N__30047),
            .in1(N__29494),
            .in2(_gnd_net_),
            .in3(N__29480),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__44837),
            .ce(N__29931),
            .sr(N__44223));
    defparam \current_shift_inst.timer_s1.counter_13_LC_13_25_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_13_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_13_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_13_25_5  (
            .in0(N__30051),
            .in1(N__29464),
            .in2(_gnd_net_),
            .in3(N__29450),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__44837),
            .ce(N__29931),
            .sr(N__44223));
    defparam \current_shift_inst.timer_s1.counter_14_LC_13_25_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_13_25_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_13_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_13_25_6  (
            .in0(N__30048),
            .in1(N__29436),
            .in2(_gnd_net_),
            .in3(N__29420),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__44837),
            .ce(N__29931),
            .sr(N__44223));
    defparam \current_shift_inst.timer_s1.counter_15_LC_13_25_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_13_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_13_25_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_13_25_7  (
            .in0(N__30052),
            .in1(N__29893),
            .in2(_gnd_net_),
            .in3(N__29879),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__44837),
            .ce(N__29931),
            .sr(N__44223));
    defparam \current_shift_inst.timer_s1.counter_16_LC_13_26_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_13_26_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_13_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_13_26_0  (
            .in0(N__30077),
            .in1(N__29865),
            .in2(_gnd_net_),
            .in3(N__29846),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__44835),
            .ce(N__29930),
            .sr(N__44229));
    defparam \current_shift_inst.timer_s1.counter_17_LC_13_26_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_13_26_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_13_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_13_26_1  (
            .in0(N__30042),
            .in1(N__29829),
            .in2(_gnd_net_),
            .in3(N__29810),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__44835),
            .ce(N__29930),
            .sr(N__44229));
    defparam \current_shift_inst.timer_s1.counter_18_LC_13_26_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_13_26_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_13_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_13_26_2  (
            .in0(N__30078),
            .in1(N__29800),
            .in2(_gnd_net_),
            .in3(N__29786),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__44835),
            .ce(N__29930),
            .sr(N__44229));
    defparam \current_shift_inst.timer_s1.counter_19_LC_13_26_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_13_26_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_13_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_13_26_3  (
            .in0(N__30043),
            .in1(N__29781),
            .in2(_gnd_net_),
            .in3(N__29765),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__44835),
            .ce(N__29930),
            .sr(N__44229));
    defparam \current_shift_inst.timer_s1.counter_20_LC_13_26_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_13_26_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_13_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_13_26_4  (
            .in0(N__30079),
            .in1(N__29749),
            .in2(_gnd_net_),
            .in3(N__29735),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__44835),
            .ce(N__29930),
            .sr(N__44229));
    defparam \current_shift_inst.timer_s1.counter_21_LC_13_26_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_13_26_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_13_26_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_13_26_5  (
            .in0(N__30044),
            .in1(N__29719),
            .in2(_gnd_net_),
            .in3(N__29705),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__44835),
            .ce(N__29930),
            .sr(N__44229));
    defparam \current_shift_inst.timer_s1.counter_22_LC_13_26_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_13_26_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_13_26_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_13_26_6  (
            .in0(N__30080),
            .in1(N__29697),
            .in2(_gnd_net_),
            .in3(N__29678),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__44835),
            .ce(N__29930),
            .sr(N__44229));
    defparam \current_shift_inst.timer_s1.counter_23_LC_13_26_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_13_26_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_13_26_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_13_26_7  (
            .in0(N__30045),
            .in1(N__29664),
            .in2(_gnd_net_),
            .in3(N__29648),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__44835),
            .ce(N__29930),
            .sr(N__44229));
    defparam \current_shift_inst.timer_s1.counter_24_LC_13_27_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_13_27_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_13_27_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_13_27_0  (
            .in0(N__30054),
            .in1(N__30201),
            .in2(_gnd_net_),
            .in3(N__30182),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_27_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__44832),
            .ce(N__29932),
            .sr(N__44232));
    defparam \current_shift_inst.timer_s1.counter_25_LC_13_27_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_13_27_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_13_27_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_13_27_1  (
            .in0(N__30058),
            .in1(N__30168),
            .in2(_gnd_net_),
            .in3(N__30152),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__44832),
            .ce(N__29932),
            .sr(N__44232));
    defparam \current_shift_inst.timer_s1.counter_26_LC_13_27_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_13_27_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_13_27_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_13_27_2  (
            .in0(N__30055),
            .in1(N__30142),
            .in2(_gnd_net_),
            .in3(N__30128),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__44832),
            .ce(N__29932),
            .sr(N__44232));
    defparam \current_shift_inst.timer_s1.counter_27_LC_13_27_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_13_27_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_13_27_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_13_27_3  (
            .in0(N__30059),
            .in1(N__30123),
            .in2(_gnd_net_),
            .in3(N__30107),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__44832),
            .ce(N__29932),
            .sr(N__44232));
    defparam \current_shift_inst.timer_s1.counter_28_LC_13_27_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_13_27_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_13_27_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_13_27_4  (
            .in0(N__30056),
            .in1(N__30097),
            .in2(_gnd_net_),
            .in3(N__30083),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__44832),
            .ce(N__29932),
            .sr(N__44232));
    defparam \current_shift_inst.timer_s1.counter_29_LC_13_27_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_13_27_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_13_27_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_13_27_5  (
            .in0(N__29950),
            .in1(N__30057),
            .in2(_gnd_net_),
            .in3(N__29960),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44832),
            .ce(N__29932),
            .sr(N__44232));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_14_5_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_14_5_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32533),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_14_5_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_14_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32491),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_14_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_14_6_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_14_6_0 .LUT_INIT=16'b0011000111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_14_6_0  (
            .in0(N__35826),
            .in1(N__35632),
            .in2(N__35509),
            .in3(N__32681),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44929),
            .ce(),
            .sr(N__44107));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_14_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_14_6_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_14_6_2 .LUT_INIT=16'b0011000111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_14_6_2  (
            .in0(N__35825),
            .in1(N__35631),
            .in2(N__35508),
            .in3(N__32780),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44929),
            .ce(),
            .sr(N__44107));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_14_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_14_7_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_14_7_0  (
            .in0(N__30294),
            .in1(N__34947),
            .in2(N__30344),
            .in3(N__30314),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_14_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_14_7_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_14_7_2 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_14_7_2  (
            .in0(N__35588),
            .in1(N__35832),
            .in2(N__32822),
            .in3(N__35445),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44923),
            .ce(),
            .sr(N__44113));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_14_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_14_7_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_14_7_3 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_14_7_3  (
            .in0(N__35829),
            .in1(N__35589),
            .in2(N__35494),
            .in3(N__33017),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44923),
            .ce(),
            .sr(N__44113));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_14_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_14_7_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_14_7_4 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_14_7_4  (
            .in0(N__35586),
            .in1(N__35830),
            .in2(N__32987),
            .in3(N__35443),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44923),
            .ce(),
            .sr(N__44113));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_14_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_14_7_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_14_7_6 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_14_7_6  (
            .in0(N__35587),
            .in1(N__35831),
            .in2(N__32966),
            .in3(N__35444),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44923),
            .ce(),
            .sr(N__44113));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_14_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_14_7_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_14_7_7  (
            .in0(N__34386),
            .in1(N__35867),
            .in2(N__30523),
            .in3(N__30892),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_14_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_14_8_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_14_8_0  (
            .in0(N__30626),
            .in1(N__30251),
            .in2(N__34964),
            .in3(N__30218),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_14_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_14_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30625),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_14_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_14_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_14_8_2 .LUT_INIT=16'b0010001110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_14_8_2  (
            .in0(N__35431),
            .in1(N__35635),
            .in2(N__35833),
            .in3(N__32753),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44917),
            .ce(),
            .sr(N__44117));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_14_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_14_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_14_8_3 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_14_8_3  (
            .in0(N__32936),
            .in1(N__35813),
            .in2(N__35672),
            .in3(N__35432),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44917),
            .ce(),
            .sr(N__44117));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_14_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_14_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_14_8_4 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_14_8_4  (
            .in0(N__35811),
            .in1(N__35633),
            .in2(N__35492),
            .in3(N__32906),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44917),
            .ce(),
            .sr(N__44117));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_14_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_14_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_14_8_5 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_14_8_5  (
            .in0(N__32876),
            .in1(N__35814),
            .in2(N__35671),
            .in3(N__35439),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44917),
            .ce(),
            .sr(N__44117));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_14_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_14_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_14_8_6 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_14_8_6  (
            .in0(N__35812),
            .in1(N__35634),
            .in2(N__35493),
            .in3(N__32849),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44917),
            .ce(),
            .sr(N__44117));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_14_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_14_9_0 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_14_9_0  (
            .in0(N__30602),
            .in1(N__32509),
            .in2(N__34961),
            .in3(N__30572),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_14_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_14_9_1 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_14_9_1  (
            .in0(N__30560),
            .in1(N__30528),
            .in2(N__30479),
            .in3(N__34933),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_14_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_14_9_2 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_14_9_2  (
            .in0(N__30462),
            .in1(N__30439),
            .in2(N__34959),
            .in3(N__30392),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_14_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_14_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30369),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_14_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_14_9_5 .LUT_INIT=16'b0011110011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_14_9_5  (
            .in0(N__30995),
            .in1(N__30966),
            .in2(N__30947),
            .in3(N__34938),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_14_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_14_9_6 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_14_9_6  (
            .in0(N__30927),
            .in1(N__30900),
            .in2(N__34960),
            .in3(N__30863),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_14_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_14_9_7 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_14_9_7  (
            .in0(N__34390),
            .in1(N__34937),
            .in2(N__30851),
            .in3(N__30821),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_14_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_14_10_0 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_14_10_0  (
            .in0(N__30804),
            .in1(N__30768),
            .in2(N__34954),
            .in3(N__30749),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_14_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_14_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32406),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_14_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_14_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35043),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_14_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_14_10_4 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_14_10_4  (
            .in0(N__34341),
            .in1(N__30738),
            .in2(N__34955),
            .in3(N__30719),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_14_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_14_10_5 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_14_10_5  (
            .in0(N__31937),
            .in1(N__30702),
            .in2(N__30662),
            .in3(N__34926),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_14_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_14_10_6 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_14_10_6  (
            .in0(N__31267),
            .in1(N__31225),
            .in2(N__34953),
            .in3(N__31196),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_14_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_14_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35217),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_14_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_14_11_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(N__34899),
            .in2(_gnd_net_),
            .in3(N__31185),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_14_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_14_11_1 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_14_11_1  (
            .in0(N__31961),
            .in1(N__35047),
            .in2(N__34949),
            .in3(N__31160),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_14_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_14_11_2 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_14_11_2  (
            .in0(N__35170),
            .in1(N__34905),
            .in2(N__31148),
            .in3(N__31121),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_14_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_14_11_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_14_11_3  (
            .in0(N__34897),
            .in1(N__31112),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_14_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_14_11_4 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_14_11_4  (
            .in0(N__31095),
            .in1(N__34901),
            .in2(N__31043),
            .in3(N__31040),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_14_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_14_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_14_11_5  (
            .in0(N__34898),
            .in1(N__31034),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_14_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_14_11_6 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_14_11_6  (
            .in0(N__35329),
            .in1(N__34900),
            .in2(N__31022),
            .in3(N__31019),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_14_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_14_11_7 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_14_11_7  (
            .in0(N__31349),
            .in1(N__34222),
            .in2(N__34948),
            .in3(N__31319),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_14_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_14_12_0 .LUT_INIT=16'b1111111111100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_14_12_0  (
            .in0(N__36513),
            .in1(N__42488),
            .in2(N__39245),
            .in3(N__36363),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_14_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_14_12_1 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_14_12_1  (
            .in0(N__36309),
            .in1(_gnd_net_),
            .in2(N__31313),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIFG4DM1_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_14_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_14_12_2 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_14_12_2  (
            .in0(N__36509),
            .in1(N__39368),
            .in2(N__33467),
            .in3(N__36152),
            .lcout(elapsed_time_ns_1_RNIRBJF91_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_14_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_14_12_3 .LUT_INIT=16'b1111101111101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_14_12_3  (
            .in0(N__36308),
            .in1(N__36512),
            .in2(N__38660),
            .in3(N__37078),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_14_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_14_12_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31310),
            .in3(N__36362),
            .lcout(elapsed_time_ns_1_RNIRHL2M1_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_14_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_14_12_5 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_14_12_5  (
            .in0(N__34872),
            .in1(N__32608),
            .in2(N__31307),
            .in3(N__31280),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_14_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_14_12_6 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_14_12_6  (
            .in0(N__36511),
            .in1(N__38954),
            .in2(N__42535),
            .in3(N__36153),
            .lcout(elapsed_time_ns_1_RNIQ8HF91_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_14_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_14_12_7 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_14_12_7  (
            .in0(N__39134),
            .in1(N__36510),
            .in2(N__36172),
            .in3(N__33440),
            .lcout(elapsed_time_ns_1_RNIQ9IF91_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_14_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_14_13_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_14_13_0  (
            .in0(N__38975),
            .in1(N__36516),
            .in2(N__36177),
            .in3(N__41517),
            .lcout(elapsed_time_ns_1_RNIP7HF91_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_14_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_14_13_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_14_13_1  (
            .in0(N__36041),
            .in1(N__44313),
            .in2(_gnd_net_),
            .in3(N__33551),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_14_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_14_13_2 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_14_13_2  (
            .in0(N__44314),
            .in1(N__39338),
            .in2(N__31364),
            .in3(N__33557),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_14_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_14_13_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31361),
            .in3(N__31355),
            .lcout(elapsed_time_ns_1_RNIHI4DM1_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_14_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_14_13_4 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_14_13_4  (
            .in0(N__36922),
            .in1(N__36517),
            .in2(N__39011),
            .in3(N__36385),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_14_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_14_13_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31358),
            .in3(N__36310),
            .lcout(elapsed_time_ns_1_RNI1OL2M1_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_14_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_14_13_6 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_14_13_6  (
            .in0(N__33287),
            .in1(_gnd_net_),
            .in2(N__36321),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIUKL2M1_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_13_7 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_13_7  (
            .in0(N__36518),
            .in1(N__39188),
            .in2(N__36396),
            .in3(N__42330),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_14_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_14_14_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__33563),
            .in2(_gnd_net_),
            .in3(N__36314),
            .lcout(elapsed_time_ns_1_RNIIJ4DM1_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_14_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_14_14_1 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_14_14_1  (
            .in0(N__39068),
            .in1(N__36167),
            .in2(N__36867),
            .in3(N__36524),
            .lcout(elapsed_time_ns_1_RNIFJ2591_0_7),
            .ltout(elapsed_time_ns_1_RNIFJ2591_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_2_LC_14_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_2_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_2_LC_14_14_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_2_LC_14_14_2  (
            .in0(N__36794),
            .in1(N__36836),
            .in2(N__31871),
            .in3(N__36898),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_6_LC_14_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_6_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_6_LC_14_14_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_6_LC_14_14_3  (
            .in0(N__42006),
            .in1(_gnd_net_),
            .in2(N__31868),
            .in3(N__37020),
            .lcout(\phase_controller_inst1.stoper_tr.N_250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_14_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_14_14_4 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_14_14_4  (
            .in0(N__31865),
            .in1(N__31691),
            .in2(N__31657),
            .in3(N__31577),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_a5_1_LC_14_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_a5_1_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_a5_1_LC_14_14_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_0_a5_1_LC_14_14_5  (
            .in0(N__42007),
            .in1(N__37112),
            .in2(N__37154),
            .in3(N__31970),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.N_235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_1_1_LC_14_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_1_1_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_1_1_LC_14_14_6 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_0_1_1_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__33690),
            .in2(N__31535),
            .in3(N__36751),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_f0_0_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0_3_LC_14_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0_3_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0_3_LC_14_15_0 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_0_0_3_LC_14_15_0  (
            .in0(N__42069),
            .in1(N__42167),
            .in2(N__37120),
            .in3(N__37146),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_7_f0_0_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_3_LC_14_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_3_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_3_LC_14_15_1 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_3_LC_14_15_1  (
            .in0(N__37086),
            .in1(N__37619),
            .in2(N__31532),
            .in3(N__36770),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44883),
            .ce(N__43743),
            .sr(N__44144));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI74R51_0_1_LC_14_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI74R51_0_1_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI74R51_0_1_LC_14_15_2 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_RNI74R51_0_1_LC_14_15_2  (
            .in0(N__32056),
            .in1(N__44316),
            .in2(N__31471),
            .in3(N__32029),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI74R51_1_LC_14_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI74R51_1_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI74R51_1_LC_14_15_3 .LUT_INIT=16'b1010101010111110;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_RNI74R51_1_LC_14_15_3  (
            .in0(N__44317),
            .in1(N__32055),
            .in2(N__32030),
            .in3(N__31463),
            .lcout(\phase_controller_inst2.stoper_hc.un1_stoper_state12_1_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_14_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_14_15_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_14_15_4  (
            .in0(N__32054),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32025),
            .lcout(\phase_controller_inst2.stoper_hc.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_o2_1_LC_14_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_o2_1_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_0_o2_1_LC_14_16_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_0_o2_1_LC_14_16_1  (
            .in0(N__37079),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37170),
            .lcout(\phase_controller_inst1.stoper_tr.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_16_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_16_2  (
            .in0(N__34916),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31956),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_14_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_14_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__31929),
            .in2(_gnd_net_),
            .in3(N__34915),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_14_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_14_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32613),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_14_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_14_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33612),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_c_RNO_LC_14_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_c_RNO_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_c_RNO_LC_14_16_6 .LUT_INIT=16'b0001110100011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_c_RNO_LC_14_16_6  (
            .in0(N__33613),
            .in1(N__40061),
            .in2(N__31910),
            .in3(N__39857),
            .lcout(\current_shift_inst.un38_control_input_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_c_RNO_LC_14_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_c_RNO_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_c_RNO_LC_14_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_c_RNO_LC_14_17_0  (
            .in0(N__40117),
            .in1(N__37376),
            .in2(_gnd_net_),
            .in3(N__37352),
            .lcout(\current_shift_inst.un38_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_c_RNO_LC_14_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_c_RNO_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_c_RNO_LC_14_17_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_c_RNO_LC_14_17_1  (
            .in0(N__37934),
            .in1(N__40119),
            .in2(_gnd_net_),
            .in3(N__37904),
            .lcout(\current_shift_inst.un38_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_c_RNO_LC_14_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_c_RNO_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_c_RNO_LC_14_17_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_c_RNO_LC_14_17_2  (
            .in0(N__40118),
            .in1(_gnd_net_),
            .in2(N__37339),
            .in3(N__37313),
            .lcout(\current_shift_inst.un38_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_c_RNO_LC_14_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_c_RNO_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_c_RNO_LC_14_17_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_c_RNO_LC_14_17_3  (
            .in0(N__37660),
            .in1(N__40120),
            .in2(_gnd_net_),
            .in3(N__37634),
            .lcout(\current_shift_inst.un38_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_c_RNO_LC_14_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_c_RNO_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_c_RNO_LC_14_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_c_RNO_LC_14_17_4  (
            .in0(N__40121),
            .in1(N__37891),
            .in2(_gnd_net_),
            .in3(N__37865),
            .lcout(\current_shift_inst.un38_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_c_RNO_LC_14_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_c_RNO_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_c_RNO_LC_14_17_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_c_RNO_LC_14_17_5  (
            .in0(N__37835),
            .in1(N__40122),
            .in2(_gnd_net_),
            .in3(N__37847),
            .lcout(\current_shift_inst.un38_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_c_RNO_LC_14_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_c_RNO_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_c_RNO_LC_14_17_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_c_RNO_LC_14_17_6  (
            .in0(N__40116),
            .in1(N__37400),
            .in2(_gnd_net_),
            .in3(N__37412),
            .lcout(\current_shift_inst.un38_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37332),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_14_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_14_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37449),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37920),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_14_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_14_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37387),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37363),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_14_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_14_18_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_14_18_4  (
            .in0(N__40124),
            .in1(N__38263),
            .in2(_gnd_net_),
            .in3(N__38236),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_14_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_14_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37290),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_14_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_14_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37245),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_c_RNO_LC_14_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_c_RNO_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_c_RNO_LC_14_18_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_c_RNO_LC_14_18_7  (
            .in0(N__37450),
            .in1(N__40123),
            .in2(_gnd_net_),
            .in3(N__37436),
            .lcout(\current_shift_inst.un38_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_c_RNO_LC_14_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_c_RNO_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_c_RNO_LC_14_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_c_RNO_LC_14_19_0  (
            .in0(N__40057),
            .in1(N__37762),
            .in2(_gnd_net_),
            .in3(N__37742),
            .lcout(\current_shift_inst.un38_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_14_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_14_19_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_14_19_1  (
            .in0(N__37730),
            .in1(N__38473),
            .in2(_gnd_net_),
            .in3(N__38455),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37650),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38017),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37881),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38472),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37794),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_14_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_14_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38739),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_14_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_14_20_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_14_20_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_14_20_0  (
            .in0(N__43838),
            .in1(N__44378),
            .in2(_gnd_net_),
            .in3(N__43671),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44855),
            .ce(),
            .sr(N__44588));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37962),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38143),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_14_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_14_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37758),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38056),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_1_LC_14_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_1_LC_14_21_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_1_LC_14_21_0 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_1_LC_14_21_0  (
            .in0(N__33698),
            .in1(N__37620),
            .in2(N__42267),
            .in3(N__33671),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44851),
            .ce(N__41941),
            .sr(N__44181));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_4_LC_14_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_4_LC_14_21_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_4_LC_14_21_1 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_4_LC_14_21_1  (
            .in0(N__37622),
            .in1(N__42252),
            .in2(N__37502),
            .in3(N__37540),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44851),
            .ce(N__41941),
            .sr(N__44181));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_3_LC_14_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_3_LC_14_21_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_3_LC_14_21_2 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_3_LC_14_21_2  (
            .in0(N__32168),
            .in1(N__37621),
            .in2(N__36775),
            .in3(N__37091),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44851),
            .ce(N__41941),
            .sr(N__44181));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_14_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_14_21_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_14_21_3  (
            .in0(N__40063),
            .in1(_gnd_net_),
            .in2(N__34037),
            .in3(N__32180),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_14_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_14_21_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_14_21_4  (
            .in0(N__32179),
            .in1(N__40062),
            .in2(_gnd_net_),
            .in3(N__34033),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32178),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_14_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_14_22_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(N__38295),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38830),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_14_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_14_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38536),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_14_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_14_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38373),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38418),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_15_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_15_6_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_15_6_3 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_15_6_3  (
            .in0(N__35818),
            .in1(N__35644),
            .in2(N__35510),
            .in3(N__33227),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44934),
            .ce(),
            .sr(N__44105));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_15_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_15_6_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_15_6_4 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_15_6_4  (
            .in0(N__35642),
            .in1(N__35820),
            .in2(N__33188),
            .in3(N__35475),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44934),
            .ce(),
            .sr(N__44105));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_15_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_15_6_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_15_6_5 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_15_6_5  (
            .in0(N__35819),
            .in1(N__35645),
            .in2(N__35511),
            .in3(N__33146),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44934),
            .ce(),
            .sr(N__44105));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_15_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_15_6_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_15_6_6 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_15_6_6  (
            .in0(N__35643),
            .in1(N__35821),
            .in2(N__33113),
            .in3(N__35476),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44934),
            .ce(),
            .sr(N__44105));
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_15_7_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_15_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(N__32461),
            .in2(N__32465),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_15_7_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_15_7_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_15_7_1 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_15_7_1  (
            .in0(N__35675),
            .in1(N__32444),
            .in2(N__32429),
            .in3(N__32375),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .clk(N__44930),
            .ce(),
            .sr(N__44108));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_15_7_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_15_7_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_15_7_2 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_15_7_2  (
            .in0(N__35677),
            .in1(N__32372),
            .in2(N__32360),
            .in3(N__32300),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .clk(N__44930),
            .ce(),
            .sr(N__44108));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_15_7_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_15_7_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_15_7_3 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_15_7_3  (
            .in0(N__35676),
            .in1(N__32297),
            .in2(N__34409),
            .in3(N__32285),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .clk(N__44930),
            .ce(),
            .sr(N__44108));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_15_7_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_15_7_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_15_7_4 .LUT_INIT=16'b0111110111010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_15_7_4  (
            .in0(N__35678),
            .in1(N__32282),
            .in2(N__32270),
            .in3(N__32204),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .clk(N__44930),
            .ce(),
            .sr(N__44108));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_15_7_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_15_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(N__32201),
            .in2(N__32834),
            .in3(N__32810),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_15_7_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_15_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(N__32807),
            .in2(N__32795),
            .in3(N__32774),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_15_7_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_15_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(N__34265),
            .in2(N__34670),
            .in3(N__32771),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_15_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_15_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__32768),
            .in2(N__32762),
            .in3(N__32744),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_15_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_15_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__32741),
            .in2(N__32732),
            .in3(N__32708),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_15_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_15_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__32705),
            .in2(N__32696),
            .in3(N__32672),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_15_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_15_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__34259),
            .in2(N__32669),
            .in3(N__32654),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_15_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_15_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__32651),
            .in2(N__32636),
            .in3(N__32621),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_15_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_15_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__33038),
            .in2(N__33026),
            .in3(N__33011),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_15_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_15_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(N__33008),
            .in2(N__32996),
            .in3(N__32978),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_15_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_15_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(N__34352),
            .in2(N__32975),
            .in3(N__32957),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_15_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_15_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__32954),
            .in2(N__32948),
            .in3(N__32930),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_15_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_15_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__32927),
            .in2(N__32915),
            .in3(N__32900),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_15_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_15_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__32897),
            .in2(N__32885),
            .in3(N__32870),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_15_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_15_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__32867),
            .in2(N__32858),
            .in3(N__32843),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_15_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_15_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__32840),
            .in2(N__34295),
            .in3(N__33218),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_15_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_15_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__33215),
            .in2(N__33200),
            .in3(N__33176),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_15_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_15_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__33173),
            .in2(N__33161),
            .in3(N__33137),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_15_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_15_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__33134),
            .in2(N__33122),
            .in3(N__33098),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_15_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_15_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__33233),
            .in2(N__33095),
            .in3(N__33086),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_15_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_15_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__34274),
            .in2(N__33083),
            .in3(N__33074),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_15_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_15_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__33071),
            .in2(N__33491),
            .in3(N__33059),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_15_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_15_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__33056),
            .in2(N__33050),
            .in3(N__33041),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_15_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_15_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__33413),
            .in2(N__33398),
            .in3(N__33368),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_15_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_15_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__33330),
            .in2(N__33365),
            .in3(N__33350),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_15_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_15_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__33332),
            .in2(N__33347),
            .in3(N__33335),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_15_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_15_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__33331),
            .in2(N__33311),
            .in3(N__33293),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_15_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_15_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_15_11_0  (
            .in0(N__34914),
            .in1(N__35778),
            .in2(_gnd_net_),
            .in3(N__33290),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_15_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_15_11_1 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_15_11_1  (
            .in0(N__36815),
            .in1(N__36530),
            .in2(N__38582),
            .in3(N__36370),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_15_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_15_11_3 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_15_11_3  (
            .in0(N__39268),
            .in1(N__35243),
            .in2(N__38887),
            .in3(N__35996),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_363_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_15_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_15_11_4 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_15_11_4  (
            .in0(N__39342),
            .in1(N__36249),
            .in2(N__33278),
            .in3(N__36266),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_15_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_15_11_5 .LUT_INIT=16'b0011110011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_15_11_5  (
            .in0(N__35221),
            .in1(N__33275),
            .in2(N__33248),
            .in3(N__34912),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_15_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_15_11_7 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_15_11_7  (
            .in0(N__35110),
            .in1(N__34913),
            .in2(N__33530),
            .in3(N__33503),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_15_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_15_12_0 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_15_12_0  (
            .in0(N__36145),
            .in1(N__33452),
            .in2(N__39116),
            .in3(N__36507),
            .lcout(elapsed_time_ns_1_RNIRAIF91_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_15_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_15_12_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_15_12_1  (
            .in0(N__35914),
            .in1(N__44311),
            .in2(N__36376),
            .in3(N__35273),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_15_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_15_12_2 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_15_12_2  (
            .in0(N__44312),
            .in1(N__39344),
            .in2(N__33479),
            .in3(N__36040),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_15_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_15_12_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_15_12_3  (
            .in0(N__36508),
            .in1(N__38933),
            .in2(N__33476),
            .in3(N__41592),
            .lcout(elapsed_time_ns_1_RNIR9HF91_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_15_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_15_12_4 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_15_12_4  (
            .in0(N__33428),
            .in1(N__36506),
            .in2(N__36171),
            .in3(N__39092),
            .lcout(elapsed_time_ns_1_RNISBIF91_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_15_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_15_12_5 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_15_12_5  (
            .in0(N__39392),
            .in1(N__33473),
            .in2(N__36543),
            .in3(N__36144),
            .lcout(elapsed_time_ns_1_RNI3JIF91_0_29),
            .ltout(elapsed_time_ns_1_RNI3JIF91_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_7_15_LC_15_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_7_15_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_7_15_LC_15_12_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_o5_7_15_LC_15_12_6  (
            .in0(N__33463),
            .in1(N__33451),
            .in2(N__33443),
            .in3(N__33439),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_7_i_o5_7Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_15_LC_15_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_15_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_15_LC_15_12_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_o5_15_LC_15_12_7  (
            .in0(N__35981),
            .in1(N__33427),
            .in2(N__33416),
            .in3(N__36203),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_i_o5_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_15_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_15_13_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_15_13_0  (
            .in0(N__35920),
            .in1(N__36250),
            .in2(N__35960),
            .in3(N__36264),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_359_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_15_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_15_13_1 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_15_13_1  (
            .in0(N__36156),
            .in1(N__36520),
            .in2(N__39044),
            .in3(N__36841),
            .lcout(elapsed_time_ns_1_RNIGK2591_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_15_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_15_13_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_15_13_2  (
            .in0(N__35272),
            .in1(N__36251),
            .in2(N__35924),
            .in3(N__36265),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_381 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_15_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_15_13_3 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_15_13_3  (
            .in0(N__36036),
            .in1(N__33550),
            .in2(N__33539),
            .in3(N__39337),
            .lcout(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ),
            .ltout(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_15_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_15_13_4 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_15_13_4  (
            .in0(N__38912),
            .in1(N__42396),
            .in2(N__33536),
            .in3(N__36154),
            .lcout(elapsed_time_ns_1_RNISAHF91_0_13),
            .ltout(elapsed_time_ns_1_RNISAHF91_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_2_2_LC_15_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_2_2_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_2_2_LC_15_13_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_a2_2_2_LC_15_13_5  (
            .in0(N__41585),
            .in1(N__41511),
            .in2(N__33533),
            .in3(N__42521),
            .lcout(\phase_controller_inst1.stoper_tr.N_244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_15_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_15_13_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_15_13_6  (
            .in0(N__36307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33572),
            .lcout(elapsed_time_ns_1_RNIGH4DM1_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_15_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_15_13_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_15_13_7  (
            .in0(N__36155),
            .in1(N__36519),
            .in2(N__37539),
            .in3(N__38627),
            .lcout(elapsed_time_ns_1_RNICG2591_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_9_LC_15_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_9_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_9_LC_15_14_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_9_LC_15_14_0  (
            .in0(N__42324),
            .in1(N__42498),
            .in2(N__42372),
            .in3(N__42290),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_15_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_15_14_1 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_15_14_1  (
            .in0(N__36515),
            .in1(N__36163),
            .in2(N__37029),
            .in3(N__39272),
            .lcout(elapsed_time_ns_1_RNIUCHF91_0_15),
            .ltout(elapsed_time_ns_1_RNIUCHF91_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_9_LC_15_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_9_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_9_LC_15_14_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_9_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__36917),
            .in2(N__33590),
            .in3(N__41552),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.N_251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_2_LC_15_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_2_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_2_LC_15_14_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_2_LC_15_14_3  (
            .in0(N__42499),
            .in1(N__42365),
            .in2(N__33587),
            .in3(N__33581),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_15_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_15_14_4 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_15_14_4  (
            .in0(N__38606),
            .in1(N__36942),
            .in2(N__36176),
            .in3(N__36514),
            .lcout(elapsed_time_ns_1_RNIDH2591_0_5),
            .ltout(elapsed_time_ns_1_RNIDH2591_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3_2_LC_15_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3_2_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3_2_LC_15_14_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3_2_LC_15_14_5  (
            .in0(N__42289),
            .in1(N__42323),
            .in2(N__33584),
            .in3(N__37523),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_i_a2_1_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_10_LC_15_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_10_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_10_LC_15_14_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_a2_10_LC_15_14_6  (
            .in0(N__37021),
            .in1(N__36968),
            .in2(_gnd_net_),
            .in3(N__41553),
            .lcout(\phase_controller_inst1.stoper_tr.N_241 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_1_9_LC_15_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_1_9_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_1_9_LC_15_14_7 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_i_1_9_LC_15_14_7  (
            .in0(N__36918),
            .in1(_gnd_net_),
            .in2(N__33575),
            .in3(N__42009),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_15_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_15_15_0 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_15_15_0  (
            .in0(N__42303),
            .in1(N__36541),
            .in2(N__36397),
            .in3(N__39212),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_15_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_15_15_2 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_15_15_2  (
            .in0(N__42371),
            .in1(N__36542),
            .in2(N__36398),
            .in3(N__39161),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_15_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_15_15_3 .LUT_INIT=16'b1111111101001110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_15_15_3  (
            .in0(N__36540),
            .in1(N__33691),
            .in2(N__38684),
            .in3(N__36389),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_15_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_15_15_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33701),
            .in3(N__36322),
            .lcout(elapsed_time_ns_1_RNIPFL2M1_0_1),
            .ltout(elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_1_LC_15_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_1_LC_15_15_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_1_LC_15_15_5 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_1_LC_15_15_5  (
            .in0(N__42166),
            .in1(N__37592),
            .in2(N__33674),
            .in3(N__33664),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44889),
            .ce(N__43736),
            .sr(N__44138));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_15_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_15_15_6 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_15_15_6  (
            .in0(N__39343),
            .in1(N__42165),
            .in2(N__36178),
            .in3(N__36539),
            .lcout(elapsed_time_ns_1_RNISCJF91_0_31),
            .ltout(elapsed_time_ns_1_RNISCJF91_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_2_LC_15_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_2_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_a2_2_LC_15_15_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_a2_2_LC_15_15_7  (
            .in0(N__37022),
            .in1(N__37113),
            .in2(N__33653),
            .in3(N__42008),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_i_a2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_15_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_15_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_15_16_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__33650),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44884),
            .ce(N__38180),
            .sr(N__44145));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_15_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_15_16_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_15_16_1  (
            .in0(N__37693),
            .in1(N__33614),
            .in2(_gnd_net_),
            .in3(N__33777),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_16_2  (
            .in0(N__40461),
            .in1(_gnd_net_),
            .in2(N__33599),
            .in3(N__33596),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_16_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_16_3  (
            .in0(N__38210),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44884),
            .ce(N__38180),
            .sr(N__44145));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_15_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_15_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_15_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38209),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44884),
            .ce(N__38180),
            .sr(N__44145));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_16_5 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_16_5  (
            .in0(N__37694),
            .in1(_gnd_net_),
            .in2(N__33754),
            .in3(N__33799),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33842),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44884),
            .ce(N__38180),
            .sr(N__44145));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33798),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_15_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_15_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__33785),
            .in2(N__33778),
            .in3(N__33779),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_15_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_15_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__33737),
            .in2(_gnd_net_),
            .in3(N__33731),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_15_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_15_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__33728),
            .in2(_gnd_net_),
            .in3(N__33722),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_15_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_15_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__33719),
            .in2(_gnd_net_),
            .in3(N__33713),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_15_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_15_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__33710),
            .in2(_gnd_net_),
            .in3(N__33704),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_15_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_15_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__33929),
            .in2(_gnd_net_),
            .in3(N__33923),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_15_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_15_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__33920),
            .in2(_gnd_net_),
            .in3(N__33911),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_15_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_15_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__33908),
            .in2(_gnd_net_),
            .in3(N__33902),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_15_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_15_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__33899),
            .in2(_gnd_net_),
            .in3(N__33893),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_15_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_15_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__33890),
            .in2(_gnd_net_),
            .in3(N__33884),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_15_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_15_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__33881),
            .in2(_gnd_net_),
            .in3(N__33875),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_15_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_15_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__33872),
            .in2(_gnd_net_),
            .in3(N__33866),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_15_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_15_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__33863),
            .in2(_gnd_net_),
            .in3(N__33854),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_15_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_15_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__33851),
            .in2(_gnd_net_),
            .in3(N__33845),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_15_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_15_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__37853),
            .in2(_gnd_net_),
            .in3(N__33992),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_15_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_15_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__33989),
            .in2(_gnd_net_),
            .in3(N__33983),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_15_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_15_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__33980),
            .in2(_gnd_net_),
            .in3(N__33974),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_15_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_15_19_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33971),
            .in3(N__33962),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_15_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_15_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__33959),
            .in2(_gnd_net_),
            .in3(N__33947),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_15_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_15_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__34160),
            .in2(_gnd_net_),
            .in3(N__33944),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_15_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_15_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__33941),
            .in2(_gnd_net_),
            .in3(N__33935),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_15_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_15_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__34118),
            .in2(_gnd_net_),
            .in3(N__33932),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_15_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_15_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(N__34094),
            .in2(_gnd_net_),
            .in3(N__34085),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_15_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_15_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__34082),
            .in2(_gnd_net_),
            .in3(N__34073),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_15_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_15_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__34109),
            .in2(_gnd_net_),
            .in3(N__34070),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_15_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_15_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__34067),
            .in2(_gnd_net_),
            .in3(N__34058),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_15_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_15_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__34055),
            .in2(_gnd_net_),
            .in3(N__34046),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_15_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_15_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__34043),
            .in2(_gnd_net_),
            .in3(N__34025),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_15_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_15_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__34022),
            .in2(_gnd_net_),
            .in3(N__34013),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_15_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_15_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34010),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_20_6 .LUT_INIT=16'b1111001111110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__39980),
            .in2(N__33995),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_15_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_15_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_15_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38793),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_21_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_21_1  (
            .in0(N__38512),
            .in1(N__38489),
            .in2(_gnd_net_),
            .in3(N__40107),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_21_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_21_2  (
            .in0(N__40110),
            .in1(N__38549),
            .in2(_gnd_net_),
            .in3(N__38525),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_15_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_15_21_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_15_21_3  (
            .in0(N__38309),
            .in1(N__40109),
            .in2(_gnd_net_),
            .in3(N__38279),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_21_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_21_5  (
            .in0(N__38383),
            .in1(N__40108),
            .in2(_gnd_net_),
            .in3(N__38357),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_21_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_21_6  (
            .in0(N__38259),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38508),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_22_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_15_22_4  (
            .in0(N__36715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34103),
            .ce(),
            .sr(N__44182));
    defparam \delay_measurement_inst.start_timer_tr_LC_15_22_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_15_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_15_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36714),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34103),
            .ce(),
            .sr(N__44182));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_16_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_16_7_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_16_7_0  (
            .in0(N__34478),
            .in1(N__34454),
            .in2(N__34962),
            .in3(N__34424),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_16_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_16_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_16_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34385),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_16_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_16_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34324),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_16_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_16_7_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(N__34566),
            .in2(_gnd_net_),
            .in3(N__35079),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_16_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_16_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35149),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_16_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_16_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_16_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34631),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_16_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_16_7_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_16_7_7  (
            .in0(N__35306),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_16_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_16_8_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_16_8_1 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_16_8_1  (
            .in0(N__35737),
            .in1(N__35648),
            .in2(N__35512),
            .in3(N__34253),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44931),
            .ce(),
            .sr(N__44109));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_16_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_16_8_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_16_8_3  (
            .in0(N__35736),
            .in1(N__34247),
            .in2(_gnd_net_),
            .in3(N__34193),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_16_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_16_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_16_8_4 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_16_8_4  (
            .in0(N__35646),
            .in1(N__35740),
            .in2(N__35515),
            .in3(N__35237),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44931),
            .ce(),
            .sr(N__44109));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_16_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_16_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_16_8_5 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_16_8_5  (
            .in0(N__35738),
            .in1(N__35649),
            .in2(N__35513),
            .in3(N__35180),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44931),
            .ce(),
            .sr(N__44109));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_16_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_16_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_16_8_6 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_16_8_6  (
            .in0(N__35647),
            .in1(N__35741),
            .in2(N__35516),
            .in3(N__35120),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44931),
            .ce(),
            .sr(N__44109));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_16_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_16_8_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_16_8_7 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_16_8_7  (
            .in0(N__35739),
            .in1(N__35650),
            .in2(N__35514),
            .in3(N__35063),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44931),
            .ce(),
            .sr(N__44109));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_16_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_16_9_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_16_9_0  (
            .in0(N__34630),
            .in1(N__34994),
            .in2(N__34963),
            .in3(N__34682),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_16_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_16_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_16_9_2 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_16_9_2  (
            .in0(N__34658),
            .in1(N__35763),
            .in2(N__35673),
            .in3(N__35506),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44924),
            .ce(),
            .sr(N__44114));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_16_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_16_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_16_9_3 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_16_9_3  (
            .in0(N__35759),
            .in1(N__35653),
            .in2(N__35518),
            .in3(N__34601),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44924),
            .ce(),
            .sr(N__44114));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_16_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_16_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_16_9_4 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_16_9_4  (
            .in0(N__35651),
            .in1(N__35761),
            .in2(N__34544),
            .in3(N__35504),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44924),
            .ce(),
            .sr(N__44114));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_16_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_16_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_16_9_5 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_16_9_5  (
            .in0(N__35760),
            .in1(N__35654),
            .in2(N__35519),
            .in3(N__35900),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44924),
            .ce(),
            .sr(N__44114));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_16_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_16_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_16_9_6 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_16_9_6  (
            .in0(N__35891),
            .in1(N__35762),
            .in2(N__35674),
            .in3(N__35505),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44924),
            .ce(),
            .sr(N__44114));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_16_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_16_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_16_9_7 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_16_9_7  (
            .in0(N__35758),
            .in1(N__35652),
            .in2(N__35517),
            .in3(N__35339),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44924),
            .ce(),
            .sr(N__44114));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_16_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_16_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_16_10_0  (
            .in0(N__36009),
            .in1(N__38671),
            .in2(N__38650),
            .in3(N__35251),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_10_1 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_10_1  (
            .in0(N__38646),
            .in1(N__39157),
            .in2(N__39184),
            .in3(N__36010),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_16_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_16_10_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_16_10_2  (
            .in0(N__39234),
            .in1(N__35258),
            .in2(N__35276),
            .in3(N__35252),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_380 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_16_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_16_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_16_10_3  (
            .in0(N__38873),
            .in1(N__39204),
            .in2(N__39004),
            .in3(N__38571),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_10_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_10_4  (
            .in0(N__38596),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38620),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_10_5  (
            .in0(N__39177),
            .in1(N__39156),
            .in2(N__39238),
            .in3(N__39205),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_367 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_367_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_10_6  (
            .in0(N__38572),
            .in1(N__38874),
            .in2(N__36044),
            .in3(N__38999),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_10_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_10_7  (
            .in0(N__40750),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44918),
            .ce(N__39291),
            .sr(N__44118));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_16_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_16_11_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_16_11_0  (
            .in0(N__39000),
            .in1(N__35933),
            .in2(_gnd_net_),
            .in3(N__35939),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_16_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_16_11_1 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_16_11_1  (
            .in0(N__39452),
            .in1(N__35990),
            .in2(N__36547),
            .in3(N__36124),
            .lcout(elapsed_time_ns_1_RNIVEIF91_0_25),
            .ltout(elapsed_time_ns_1_RNIVEIF91_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_6_15_LC_16_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_6_15_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_6_15_LC_16_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_o5_6_15_LC_16_11_2  (
            .in0(N__35971),
            .in1(N__36193),
            .in2(N__35984),
            .in3(N__36232),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_i_o5_6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_16_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_16_11_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_16_11_3  (
            .in0(N__36529),
            .in1(N__39410),
            .in2(N__35975),
            .in3(N__36125),
            .lcout(elapsed_time_ns_1_RNI2IIF91_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_16_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_16_11_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_16_11_4  (
            .in0(N__39060),
            .in1(N__38570),
            .in2(N__39037),
            .in3(N__35950),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_11_5  (
            .in0(N__38926),
            .in1(N__38947),
            .in2(N__38908),
            .in3(N__38968),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_347 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_16_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_16_11_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_16_11_6  (
            .in0(N__39061),
            .in1(N__39261),
            .in2(N__35927),
            .in3(N__39033),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36698),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_16_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_16_12_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_16_12_0  (
            .in0(N__39451),
            .in1(N__39130),
            .in2(N__39437),
            .in3(N__36221),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_16_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_16_12_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_16_12_1  (
            .in0(N__39361),
            .in1(N__39406),
            .in2(N__39388),
            .in3(N__39421),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_16_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_16_12_2 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_16_12_2  (
            .in0(N__39436),
            .in1(N__36236),
            .in2(N__36554),
            .in3(N__36128),
            .lcout(elapsed_time_ns_1_RNI0GIF91_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_12_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_12_3  (
            .in0(N__39112),
            .in1(N__39478),
            .in2(N__39091),
            .in3(N__39466),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_16_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_16_12_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_16_12_4  (
            .in0(N__39479),
            .in1(N__36126),
            .in2(N__36215),
            .in3(N__36548),
            .lcout(elapsed_time_ns_1_RNITCIF91_0_23),
            .ltout(elapsed_time_ns_1_RNITCIF91_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_15_LC_16_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_15_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_15_LC_16_12_5 .LUT_INIT=16'b1111110011111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_15_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__36055),
            .in2(N__36206),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_i_o5_0_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_16_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_16_12_7 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_16_12_7  (
            .in0(N__36127),
            .in1(N__39422),
            .in2(N__36197),
            .in3(N__36549),
            .lcout(elapsed_time_ns_1_RNI1HIF91_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_13_0 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_13_0  (
            .in0(N__39467),
            .in1(N__36502),
            .in2(N__36059),
            .in3(N__36129),
            .lcout(elapsed_time_ns_1_RNIUDIF91_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_13_2 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_13_2  (
            .in0(N__36696),
            .in1(N__36724),
            .in2(_gnd_net_),
            .in3(N__36673),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_435_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_16_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_16_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_16_13_3 .LUT_INIT=16'b0101010111110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_16_13_3  (
            .in0(N__36674),
            .in1(_gnd_net_),
            .in2(N__36728),
            .in3(N__36697),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44906),
            .ce(),
            .sr(N__44125));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_16_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_16_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__36692),
            .in2(_gnd_net_),
            .in3(N__36672),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_434_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_16_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_16_13_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_16_13_5  (
            .in0(N__36631),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36596),
            .lcout(\phase_controller_inst1.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_14_0 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_14_0  (
            .in0(N__41551),
            .in1(N__36525),
            .in2(N__38888),
            .in3(N__36377),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_16_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_16_14_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36329),
            .in3(N__36326),
            .lcout(elapsed_time_ns_1_RNIDE4DM1_0_14),
            .ltout(elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_6_LC_16_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_6_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_6_LC_16_14_2 .LUT_INIT=16'b0000001100000011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_6_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__37018),
            .in2(N__36269),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a1_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_8_LC_16_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_8_LC_16_14_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_8_LC_16_14_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_8_LC_16_14_3  (
            .in0(N__37586),
            .in1(N__42197),
            .in2(_gnd_net_),
            .in3(N__36837),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44901),
            .ce(N__43745),
            .sr(N__44129));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_7_LC_16_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_7_LC_16_14_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_7_LC_16_14_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_7_LC_16_14_4  (
            .in0(N__42196),
            .in1(N__36871),
            .in2(_gnd_net_),
            .in3(N__37585),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44901),
            .ce(N__43745),
            .sr(N__44129));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a0_6_LC_16_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a0_6_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a0_6_LC_16_14_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_i_o2_a0_6_LC_16_14_5  (
            .in0(N__37019),
            .in1(N__36926),
            .in2(_gnd_net_),
            .in3(N__36899),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_7_f0_i_a5_1_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_0_6_LC_16_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_0_6_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_0_6_LC_16_14_6 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_f0_i_a2_0_6_LC_16_14_6  (
            .in0(N__36969),
            .in1(N__36887),
            .in2(N__36881),
            .in3(N__42025),
            .lcout(\phase_controller_inst1.stoper_tr.N_249 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_249_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_6_LC_16_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_6_LC_16_14_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_6_LC_16_14_7 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_6_LC_16_14_7  (
            .in0(N__36813),
            .in1(N__42198),
            .in2(N__36878),
            .in3(N__36776),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44901),
            .ce(N__43745),
            .sr(N__44129));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_9_LC_16_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_9_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_9_LC_16_15_0 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_9_LC_16_15_0  (
            .in0(N__37195),
            .in1(N__42038),
            .in2(N__37217),
            .in3(N__42194),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44895),
            .ce(N__41934),
            .sr(N__44131));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_12_LC_16_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_12_LC_16_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_12_LC_16_15_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_12_LC_16_15_1  (
            .in0(N__42187),
            .in1(N__42429),
            .in2(N__42074),
            .in3(N__41596),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44895),
            .ce(N__41934),
            .sr(N__44131));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_15_LC_16_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_15_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_15_LC_16_15_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_15_LC_16_15_2  (
            .in0(N__36970),
            .in1(N__42190),
            .in2(N__37033),
            .in3(N__42042),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44895),
            .ce(N__41934),
            .sr(N__44131));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_7_LC_16_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_7_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_7_LC_16_15_3 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_7_LC_16_15_3  (
            .in0(N__42186),
            .in1(_gnd_net_),
            .in2(N__36875),
            .in3(N__37588),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44895),
            .ce(N__41934),
            .sr(N__44131));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_8_LC_16_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_8_LC_16_15_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_8_LC_16_15_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_8_LC_16_15_4  (
            .in0(N__37589),
            .in1(N__42189),
            .in2(_gnd_net_),
            .in3(N__36842),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44895),
            .ce(N__41934),
            .sr(N__44131));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_6_LC_16_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_6_LC_16_15_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_6_LC_16_15_5 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_6_LC_16_15_5  (
            .in0(N__36814),
            .in1(N__37587),
            .in2(N__42227),
            .in3(N__36774),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44895),
            .ce(N__41934),
            .sr(N__44131));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_2_LC_16_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_2_LC_16_15_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_2_LC_16_15_6 .LUT_INIT=16'b0000110000001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_2_LC_16_15_6  (
            .in0(N__37590),
            .in1(N__37488),
            .in2(N__37049),
            .in3(N__42195),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44895),
            .ce(N__41934),
            .sr(N__44131));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_5_LC_16_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_5_LC_16_15_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_5_LC_16_15_7 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_5_LC_16_15_7  (
            .in0(N__42188),
            .in1(N__37591),
            .in2(N__37497),
            .in3(N__36943),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44895),
            .ce(N__41934),
            .sr(N__44131));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_9_LC_16_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_9_LC_16_16_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_9_LC_16_16_0 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_9_LC_16_16_0  (
            .in0(N__42179),
            .in1(N__37216),
            .in2(N__37199),
            .in3(N__42073),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44890),
            .ce(N__43735),
            .sr(N__44139));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_17_LC_16_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_17_LC_16_16_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_17_LC_16_16_1 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_17_LC_16_16_1  (
            .in0(N__42070),
            .in1(N__42304),
            .in2(_gnd_net_),
            .in3(N__42185),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44890),
            .ce(N__43735),
            .sr(N__44139));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_16_LC_16_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_16_LC_16_16_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_16_LC_16_16_2 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_16_LC_16_16_2  (
            .in0(N__42180),
            .in1(N__42500),
            .in2(_gnd_net_),
            .in3(N__42072),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44890),
            .ce(N__43735),
            .sr(N__44139));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0_2_LC_16_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0_2_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0_2_LC_16_16_3 .LUT_INIT=16'b0101010111010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0_2_LC_16_16_3  (
            .in0(N__37181),
            .in1(N__37153),
            .in2(N__37127),
            .in3(N__37087),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_7_i_o2_0_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_2_LC_16_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_2_LC_16_16_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_2_LC_16_16_4 .LUT_INIT=16'b0000110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_2_LC_16_16_4  (
            .in0(N__42181),
            .in1(N__37493),
            .in2(N__37040),
            .in3(N__37616),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44890),
            .ce(N__43735),
            .sr(N__44139));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_15_LC_16_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_15_LC_16_16_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_15_LC_16_16_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_15_LC_16_16_5  (
            .in0(N__42071),
            .in1(N__42183),
            .in2(N__37037),
            .in3(N__36977),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44890),
            .ce(N__43735),
            .sr(N__44139));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_5_LC_16_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_5_LC_16_16_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_5_LC_16_16_6 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_5_LC_16_16_6  (
            .in0(N__42182),
            .in1(N__36947),
            .in2(N__37498),
            .in3(N__37618),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44890),
            .ce(N__43735),
            .sr(N__44139));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_4_LC_16_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_4_LC_16_16_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_4_LC_16_16_7 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_4_LC_16_16_7  (
            .in0(N__37617),
            .in1(N__42184),
            .in2(N__37544),
            .in3(N__37492),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44890),
            .ce(N__43735),
            .sr(N__44139));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_17_0  (
            .in0(N__37698),
            .in1(N__37457),
            .in2(_gnd_net_),
            .in3(N__37435),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_c_RNO_LC_16_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_c_RNO_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_c_RNO_LC_16_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_c_RNO_LC_16_17_1  (
            .in0(N__40003),
            .in1(N__37808),
            .in2(_gnd_net_),
            .in3(N__37778),
            .lcout(\current_shift_inst.un38_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_17_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_17_2  (
            .in0(N__37695),
            .in1(N__37411),
            .in2(_gnd_net_),
            .in3(N__37399),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_17_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_17_3  (
            .in0(N__37375),
            .in1(N__37699),
            .in2(_gnd_net_),
            .in3(N__37351),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_17_4  (
            .in0(N__37701),
            .in1(N__37340),
            .in2(_gnd_net_),
            .in3(N__37312),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_17_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_17_5  (
            .in0(N__37301),
            .in1(N__37696),
            .in2(_gnd_net_),
            .in3(N__37270),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_17_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_17_6  (
            .in0(N__37697),
            .in1(N__37258),
            .in2(_gnd_net_),
            .in3(N__37228),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_17_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_17_7  (
            .in0(N__37975),
            .in1(N__37700),
            .in2(_gnd_net_),
            .in3(N__37945),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_18_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_18_0  (
            .in0(N__37933),
            .in1(N__37720),
            .in2(_gnd_net_),
            .in3(N__37903),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_18_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_18_1  (
            .in0(N__37723),
            .in1(N__37892),
            .in2(_gnd_net_),
            .in3(N__37864),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37833),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_18_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_18_3  (
            .in0(N__37725),
            .in1(N__38029),
            .in2(_gnd_net_),
            .in3(N__38002),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_18_4 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_18_4  (
            .in0(N__37846),
            .in1(N__37726),
            .in2(_gnd_net_),
            .in3(N__37834),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_16_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_16_18_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_16_18_5  (
            .in0(N__37722),
            .in1(N__37807),
            .in2(_gnd_net_),
            .in3(N__37777),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_18_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_18_6  (
            .in0(N__37766),
            .in1(N__37724),
            .in2(_gnd_net_),
            .in3(N__37741),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_18_7  (
            .in0(N__37721),
            .in1(N__37661),
            .in2(_gnd_net_),
            .in3(N__37633),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_19_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_19_0  (
            .in0(N__38156),
            .in1(N__39963),
            .in2(_gnd_net_),
            .in3(N__38132),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38203),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44870),
            .ce(N__38179),
            .sr(N__44157));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_19_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_19_2  (
            .in0(N__38155),
            .in1(N__39961),
            .in2(_gnd_net_),
            .in3(N__38131),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_19_3 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_19_3  (
            .in0(N__39957),
            .in1(N__38074),
            .in2(_gnd_net_),
            .in3(N__38065),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_19_4 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_19_4  (
            .in0(N__38747),
            .in1(N__38710),
            .in2(_gnd_net_),
            .in3(N__39958),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_19_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_19_5  (
            .in0(N__39959),
            .in1(N__38122),
            .in2(_gnd_net_),
            .in3(N__38086),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_19_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_19_6  (
            .in0(N__38800),
            .in1(N__39960),
            .in2(_gnd_net_),
            .in3(N__38770),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_c_RNO_LC_16_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_c_RNO_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_c_RNO_LC_16_19_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_c_RNO_LC_16_19_7  (
            .in0(N__39962),
            .in1(N__38075),
            .in2(_gnd_net_),
            .in3(N__38066),
            .lcout(\current_shift_inst.un38_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_c_RNO_LC_16_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_c_RNO_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_c_RNO_LC_16_20_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_c_RNO_LC_16_20_0  (
            .in0(N__38033),
            .in1(N__39978),
            .in2(_gnd_net_),
            .in3(N__38006),
            .lcout(\current_shift_inst.un38_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_20_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_20_1  (
            .in0(N__39977),
            .in1(N__38548),
            .in2(_gnd_net_),
            .in3(N__38524),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_20_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_20_2  (
            .in0(N__38513),
            .in1(N__39974),
            .in2(_gnd_net_),
            .in3(N__38488),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_c_RNO_LC_16_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_c_RNO_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_c_RNO_LC_16_20_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_c_RNO_LC_16_20_3  (
            .in0(N__39979),
            .in1(N__38477),
            .in2(_gnd_net_),
            .in3(N__38459),
            .lcout(\current_shift_inst.un38_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_20_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_20_4  (
            .in0(N__38431),
            .in1(N__39976),
            .in2(_gnd_net_),
            .in3(N__38395),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_20_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_20_5  (
            .in0(N__39973),
            .in1(N__38384),
            .in2(_gnd_net_),
            .in3(N__38353),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_16_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_16_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38342),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_20_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_20_7  (
            .in0(N__39975),
            .in1(N__38308),
            .in2(_gnd_net_),
            .in3(N__38278),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_22_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_22_1  (
            .in0(N__39995),
            .in1(N__38267),
            .in2(_gnd_net_),
            .in3(N__38237),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_22_3 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_22_3  (
            .in0(N__39999),
            .in1(N__38819),
            .in2(_gnd_net_),
            .in3(N__38840),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_22_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_22_4  (
            .in0(N__38839),
            .in1(N__39996),
            .in2(_gnd_net_),
            .in3(N__38818),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_22_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_22_6  (
            .in0(N__38804),
            .in1(N__39998),
            .in2(_gnd_net_),
            .in3(N__38774),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_c_RNO_LC_16_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_c_RNO_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_c_RNO_LC_16_22_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_c_RNO_LC_16_22_7  (
            .in0(N__39997),
            .in1(N__38746),
            .in2(_gnd_net_),
            .in3(N__38717),
            .lcout(\current_shift_inst.un38_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_17_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_17_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_17_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40778),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44932),
            .ce(N__39292),
            .sr(N__44110));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__40777),
            .in2(N__40720),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__44925),
            .ce(N__39293),
            .sr(N__44115));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__40693),
            .in2(N__40751),
            .in3(N__38609),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__44925),
            .ce(N__39293),
            .sr(N__44115));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__41065),
            .in2(N__40721),
            .in3(N__38585),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__44925),
            .ce(N__39293),
            .sr(N__44115));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__40694),
            .in2(N__41036),
            .in3(N__38552),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__44925),
            .ce(N__39293),
            .sr(N__44115));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__41005),
            .in2(N__41066),
            .in3(N__39047),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__44925),
            .ce(N__39293),
            .sr(N__44115));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__41032),
            .in2(N__40984),
            .in3(N__39014),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__44925),
            .ce(N__39293),
            .sr(N__44115));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(N__41006),
            .in2(N__40957),
            .in3(N__38978),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__44925),
            .ce(N__39293),
            .sr(N__44115));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__40920),
            .in2(N__40985),
            .in3(N__38957),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__44925),
            .ce(N__39293),
            .sr(N__44115));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__40958),
            .in2(N__40894),
            .in3(N__38936),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__44919),
            .ce(N__39294),
            .sr(N__44119));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__40867),
            .in2(N__40928),
            .in3(N__38915),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__44919),
            .ce(N__39294),
            .sr(N__44119));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__40846),
            .in2(N__40895),
            .in3(N__38891),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__44919),
            .ce(N__39294),
            .sr(N__44119));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__40868),
            .in2(N__41285),
            .in3(N__38855),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__44919),
            .ce(N__39294),
            .sr(N__44119));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__41254),
            .in2(N__40847),
            .in3(N__39248),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__44919),
            .ce(N__39294),
            .sr(N__44119));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__41281),
            .in2(N__41233),
            .in3(N__39215),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__44919),
            .ce(N__39294),
            .sr(N__44119));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__41255),
            .in2(N__41206),
            .in3(N__39191),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__44919),
            .ce(N__39294),
            .sr(N__44119));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__41170),
            .in2(N__41234),
            .in3(N__39164),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__44919),
            .ce(N__39294),
            .sr(N__44119));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__41207),
            .in2(N__41143),
            .in3(N__39137),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__44914),
            .ce(N__39295),
            .sr(N__44121));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__41116),
            .in2(N__41177),
            .in3(N__39119),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__44914),
            .ce(N__39295),
            .sr(N__44121));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__41095),
            .in2(N__41144),
            .in3(N__39095),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__44914),
            .ce(N__39295),
            .sr(N__44121));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__41117),
            .in2(N__41495),
            .in3(N__39071),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__44914),
            .ce(N__39295),
            .sr(N__44121));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__41464),
            .in2(N__41096),
            .in3(N__39470),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__44914),
            .ce(N__39295),
            .sr(N__44121));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_12_5  (
            .in0(_gnd_net_),
            .in1(N__41491),
            .in2(N__41443),
            .in3(N__39455),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__44914),
            .ce(N__39295),
            .sr(N__44121));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__41465),
            .in2(N__41416),
            .in3(N__39440),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__44914),
            .ce(N__39295),
            .sr(N__44121));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(N__41379),
            .in2(N__41444),
            .in3(N__39425),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__44914),
            .ce(N__39295),
            .sr(N__44121));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__41417),
            .in2(N__41353),
            .in3(N__39413),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__44910),
            .ce(N__39296),
            .sr(N__44123));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__41326),
            .in2(N__41387),
            .in3(N__39395),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__44910),
            .ce(N__39296),
            .sr(N__44123));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__41306),
            .in2(N__41354),
            .in3(N__39371),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__44910),
            .ce(N__39296),
            .sr(N__44123));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__41327),
            .in2(N__41678),
            .in3(N__39350),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__44910),
            .ce(N__39296),
            .sr(N__44123));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39347),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44910),
            .ce(N__39296),
            .sr(N__44123));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_17_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_17_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__41888),
            .in2(N__39518),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__41849),
            .in2(_gnd_net_),
            .in3(N__39503),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(N__44907),
            .ce(),
            .sr(N__39664));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_14_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__43106),
            .in2(N__42764),
            .in3(N__39500),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(N__44907),
            .ce(),
            .sr(N__39664));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_14_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_14_3  (
            .in0(_gnd_net_),
            .in1(N__42728),
            .in2(_gnd_net_),
            .in3(N__39497),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(N__44907),
            .ce(),
            .sr(N__39664));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_14_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(N__42695),
            .in2(_gnd_net_),
            .in3(N__39494),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(N__44907),
            .ce(),
            .sr(N__39664));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_14_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(N__42662),
            .in2(_gnd_net_),
            .in3(N__39491),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(N__44907),
            .ce(),
            .sr(N__39664));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_14_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(N__42629),
            .in2(_gnd_net_),
            .in3(N__39488),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(N__44907),
            .ce(),
            .sr(N__39664));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_14_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(N__42605),
            .in2(_gnd_net_),
            .in3(N__39485),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(N__44907),
            .ce(),
            .sr(N__39664));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__42560),
            .in2(_gnd_net_),
            .in3(N__39482),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(N__44902),
            .ce(),
            .sr(N__39657));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__43031),
            .in2(_gnd_net_),
            .in3(N__39545),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(N__44902),
            .ce(),
            .sr(N__39657));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_15_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__42992),
            .in2(_gnd_net_),
            .in3(N__39542),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(N__44902),
            .ce(),
            .sr(N__39657));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_15_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__42959),
            .in2(_gnd_net_),
            .in3(N__39539),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(N__44902),
            .ce(),
            .sr(N__39657));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_15_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__42926),
            .in2(_gnd_net_),
            .in3(N__39536),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(N__44902),
            .ce(),
            .sr(N__39657));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_15_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__42896),
            .in2(_gnd_net_),
            .in3(N__39533),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(N__44902),
            .ce(),
            .sr(N__39657));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_15_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__42860),
            .in2(_gnd_net_),
            .in3(N__39530),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(N__44902),
            .ce(),
            .sr(N__39657));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_15_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__42842),
            .in2(_gnd_net_),
            .in3(N__39527),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(N__44902),
            .ce(),
            .sr(N__39657));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_16_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__42800),
            .in2(_gnd_net_),
            .in3(N__39524),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(N__44896),
            .ce(),
            .sr(N__39665));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_16_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__43253),
            .in2(_gnd_net_),
            .in3(N__39521),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(N__44896),
            .ce(),
            .sr(N__39665));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_16_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_16_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__43214),
            .in2(_gnd_net_),
            .in3(N__39668),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44896),
            .ce(),
            .sr(N__39665));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_17_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_17_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__39623),
            .in2(N__39611),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_17_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_17_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__40594),
            .in2(N__39596),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_17_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_17_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__39581),
            .in2(N__40620),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_17_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_17_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__40598),
            .in2(N__39575),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_17_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_17_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__39566),
            .in2(N__40621),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_17_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_17_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__40602),
            .in2(N__39560),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_17_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_17_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__39551),
            .in2(N__40622),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_17_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_17_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__40606),
            .in2(N__39740),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_17_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_17_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__40590),
            .in2(N__39728),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_17_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_17_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__39719),
            .in2(N__40619),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_17_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_17_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__40578),
            .in2(N__39713),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_17_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_17_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__39704),
            .in2(N__40616),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_17_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_17_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__40582),
            .in2(N__39698),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_17_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_17_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(N__39689),
            .in2(N__40617),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_17_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_17_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_17_18_6  (
            .in0(_gnd_net_),
            .in1(N__40586),
            .in2(N__39683),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_17_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_17_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(N__39674),
            .in2(N__40618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_17_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_17_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__39809),
            .in2(N__40574),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_17_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_17_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__40502),
            .in2(N__39800),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_17_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_17_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(N__39791),
            .in2(N__40575),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_17_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_17_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__40506),
            .in2(N__39785),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_17_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_17_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(N__39776),
            .in2(N__40576),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_17_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_17_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__40510),
            .in2(N__39770),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_17_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_17_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__39761),
            .in2(N__40577),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_17_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_17_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(N__40514),
            .in2(N__39752),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_17_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_17_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__40486),
            .in2(N__40673),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_17_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_17_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(N__40664),
            .in2(N__40571),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_17_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_17_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(N__40490),
            .in2(N__40658),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_17_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_17_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__40649),
            .in2(N__40572),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_17_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_17_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(N__40494),
            .in2(N__40643),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_17_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_17_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(N__40628),
            .in2(N__40573),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_17_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_17_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__40498),
            .in2(N__40292),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(N__39991),
            .in2(_gnd_net_),
            .in3(N__39869),
            .lcout(\current_shift_inst.N_1310_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIOA7T_1_LC_17_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIOA7T_1_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIOA7T_1_LC_17_21_0 .LUT_INIT=16'b1010101110101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_RNIOA7T_1_LC_17_21_0  (
            .in0(N__44320),
            .in1(N__43778),
            .in2(N__43832),
            .in3(N__43856),
            .lcout(\phase_controller_inst2.stoper_tr.un1_stoper_state12_1_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_17_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_17_21_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_17_21_1 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_0_LC_17_21_1  (
            .in0(N__43779),
            .in1(N__43819),
            .in2(N__43864),
            .in3(N__44380),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44864),
            .ce(),
            .sr(N__44161));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_17_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_17_21_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(N__43855),
            .in2(_gnd_net_),
            .in3(N__43777),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_tr.N_45_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_17_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_17_21_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_17_21_5 .LUT_INIT=16'b1100100011001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_17_21_5  (
            .in0(N__43826),
            .in1(N__40800),
            .in2(N__40817),
            .in3(N__44381),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44864),
            .ce(),
            .sr(N__44161));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_17_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_17_21_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_17_21_6 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_1_LC_17_21_6  (
            .in0(N__44379),
            .in1(N__43780),
            .in2(N__43833),
            .in3(N__43860),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44864),
            .ce(),
            .sr(N__44161));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_18_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_18_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_18_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_18_7_0  (
            .in0(N__41814),
            .in1(N__40765),
            .in2(_gnd_net_),
            .in3(N__40754),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__44941),
            .ce(N__41657),
            .sr(N__44103));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_18_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_18_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_18_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_18_7_1  (
            .in0(N__41809),
            .in1(N__40740),
            .in2(_gnd_net_),
            .in3(N__40724),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__44941),
            .ce(N__41657),
            .sr(N__44103));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_18_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_18_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_18_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_18_7_2  (
            .in0(N__41815),
            .in1(N__40713),
            .in2(_gnd_net_),
            .in3(N__40697),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__44941),
            .ce(N__41657),
            .sr(N__44103));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_18_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_18_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_18_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_18_7_3  (
            .in0(N__41810),
            .in1(N__40692),
            .in2(_gnd_net_),
            .in3(N__40676),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__44941),
            .ce(N__41657),
            .sr(N__44103));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_18_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_18_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_18_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_18_7_4  (
            .in0(N__41816),
            .in1(N__41058),
            .in2(_gnd_net_),
            .in3(N__41039),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__44941),
            .ce(N__41657),
            .sr(N__44103));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_18_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_18_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_18_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_18_7_5  (
            .in0(N__41811),
            .in1(N__41028),
            .in2(_gnd_net_),
            .in3(N__41009),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__44941),
            .ce(N__41657),
            .sr(N__44103));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_18_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_18_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_18_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_18_7_6  (
            .in0(N__41813),
            .in1(N__41004),
            .in2(_gnd_net_),
            .in3(N__40988),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__44941),
            .ce(N__41657),
            .sr(N__44103));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_18_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_18_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_18_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_18_7_7  (
            .in0(N__41812),
            .in1(N__40977),
            .in2(_gnd_net_),
            .in3(N__40961),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__44941),
            .ce(N__41657),
            .sr(N__44103));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_18_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_18_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_18_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_18_8_0  (
            .in0(N__41798),
            .in1(N__40950),
            .in2(_gnd_net_),
            .in3(N__40931),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__44938),
            .ce(N__41656),
            .sr(N__44104));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_18_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_18_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_18_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_18_8_1  (
            .in0(N__41794),
            .in1(N__40924),
            .in2(_gnd_net_),
            .in3(N__40898),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__44938),
            .ce(N__41656),
            .sr(N__44104));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_18_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_18_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_18_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_18_8_2  (
            .in0(N__41795),
            .in1(N__40887),
            .in2(_gnd_net_),
            .in3(N__40871),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__44938),
            .ce(N__41656),
            .sr(N__44104));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_18_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_18_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_18_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_18_8_3  (
            .in0(N__41791),
            .in1(N__40866),
            .in2(_gnd_net_),
            .in3(N__40850),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__44938),
            .ce(N__41656),
            .sr(N__44104));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_18_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_18_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_18_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_18_8_4  (
            .in0(N__41796),
            .in1(N__40839),
            .in2(_gnd_net_),
            .in3(N__40820),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__44938),
            .ce(N__41656),
            .sr(N__44104));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_18_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_18_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_18_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_18_8_5  (
            .in0(N__41792),
            .in1(N__41277),
            .in2(_gnd_net_),
            .in3(N__41258),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__44938),
            .ce(N__41656),
            .sr(N__44104));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_18_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_18_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_18_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_18_8_6  (
            .in0(N__41797),
            .in1(N__41253),
            .in2(_gnd_net_),
            .in3(N__41237),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__44938),
            .ce(N__41656),
            .sr(N__44104));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_18_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_18_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_18_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_18_8_7  (
            .in0(N__41793),
            .in1(N__41226),
            .in2(_gnd_net_),
            .in3(N__41210),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__44938),
            .ce(N__41656),
            .sr(N__44104));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_18_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_18_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_18_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_18_9_0  (
            .in0(N__41787),
            .in1(N__41199),
            .in2(_gnd_net_),
            .in3(N__41180),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_18_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__44935),
            .ce(N__41655),
            .sr(N__44106));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_18_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_18_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_18_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_18_9_1  (
            .in0(N__41803),
            .in1(N__41169),
            .in2(_gnd_net_),
            .in3(N__41147),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__44935),
            .ce(N__41655),
            .sr(N__44106));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_18_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_18_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_18_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_18_9_2  (
            .in0(N__41788),
            .in1(N__41136),
            .in2(_gnd_net_),
            .in3(N__41120),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__44935),
            .ce(N__41655),
            .sr(N__44106));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_18_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_18_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_18_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_18_9_3  (
            .in0(N__41804),
            .in1(N__41115),
            .in2(_gnd_net_),
            .in3(N__41099),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__44935),
            .ce(N__41655),
            .sr(N__44106));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_18_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_18_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_18_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_18_9_4  (
            .in0(N__41789),
            .in1(N__41088),
            .in2(_gnd_net_),
            .in3(N__41069),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__44935),
            .ce(N__41655),
            .sr(N__44106));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_18_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_18_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_18_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_18_9_5  (
            .in0(N__41805),
            .in1(N__41487),
            .in2(_gnd_net_),
            .in3(N__41468),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__44935),
            .ce(N__41655),
            .sr(N__44106));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_18_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_18_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_18_9_6  (
            .in0(N__41790),
            .in1(N__41463),
            .in2(_gnd_net_),
            .in3(N__41447),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__44935),
            .ce(N__41655),
            .sr(N__44106));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_18_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_18_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_18_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_18_9_7  (
            .in0(N__41806),
            .in1(N__41436),
            .in2(_gnd_net_),
            .in3(N__41420),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__44935),
            .ce(N__41655),
            .sr(N__44106));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_18_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_18_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_18_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_18_10_0  (
            .in0(N__41799),
            .in1(N__41409),
            .in2(_gnd_net_),
            .in3(N__41390),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__44933),
            .ce(N__41645),
            .sr(N__44111));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_18_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_18_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_18_10_1  (
            .in0(N__41807),
            .in1(N__41383),
            .in2(_gnd_net_),
            .in3(N__41357),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__44933),
            .ce(N__41645),
            .sr(N__44111));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_18_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_18_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_18_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_18_10_2  (
            .in0(N__41800),
            .in1(N__41346),
            .in2(_gnd_net_),
            .in3(N__41330),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__44933),
            .ce(N__41645),
            .sr(N__44111));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_18_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_18_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_18_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_18_10_3  (
            .in0(N__41808),
            .in1(N__41325),
            .in2(_gnd_net_),
            .in3(N__41309),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__44933),
            .ce(N__41645),
            .sr(N__44111));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_18_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_18_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_18_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_18_10_4  (
            .in0(N__41801),
            .in1(N__41302),
            .in2(_gnd_net_),
            .in3(N__41288),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__44933),
            .ce(N__41645),
            .sr(N__44111));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_18_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_18_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_18_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_18_10_5  (
            .in0(N__41671),
            .in1(N__41802),
            .in2(_gnd_net_),
            .in3(N__41681),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44933),
            .ce(N__41645),
            .sr(N__44111));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_14_LC_18_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_14_LC_18_11_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_14_LC_18_11_0 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_14_LC_18_11_0  (
            .in0(N__41567),
            .in1(N__42266),
            .in2(N__42089),
            .in3(N__42454),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44926),
            .ce(N__43744),
            .sr(N__44116));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_10_LC_18_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_10_LC_18_11_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_10_LC_18_11_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_10_LC_18_11_1  (
            .in0(N__42450),
            .in1(N__42067),
            .in2(N__42269),
            .in3(N__41527),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44926),
            .ce(N__43744),
            .sr(N__44116));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_11_LC_18_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_11_LC_18_11_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_11_LC_18_11_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_11_LC_18_11_2  (
            .in0(N__42061),
            .in1(N__42264),
            .in2(N__42539),
            .in3(N__42452),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44926),
            .ce(N__43744),
            .sr(N__44116));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_13_LC_18_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_13_LC_18_11_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_13_LC_18_11_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_13_LC_18_11_4  (
            .in0(N__42062),
            .in1(N__42265),
            .in2(N__42413),
            .in3(N__42453),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44926),
            .ce(N__43744),
            .sr(N__44116));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_12_LC_18_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_12_LC_18_11_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_12_LC_18_11_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_12_LC_18_11_5  (
            .in0(N__42451),
            .in1(N__42256),
            .in2(N__41600),
            .in3(N__42068),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44926),
            .ce(N__43744),
            .sr(N__44116));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_19_LC_18_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_19_LC_18_11_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_19_LC_18_11_6 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_19_LC_18_11_6  (
            .in0(N__42060),
            .in1(_gnd_net_),
            .in2(N__42268),
            .in3(N__42380),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44926),
            .ce(N__43744),
            .sr(N__44116));
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_18_LC_18_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_18_LC_18_11_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_time_esr_18_LC_18_11_7 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_esr_18_LC_18_11_7  (
            .in0(N__42260),
            .in1(N__42343),
            .in2(_gnd_net_),
            .in3(N__42066),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44926),
            .ce(N__43744),
            .sr(N__44116));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_14_LC_18_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_14_LC_18_12_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_14_LC_18_12_0 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_14_LC_18_12_0  (
            .in0(N__42457),
            .in1(N__41566),
            .in2(N__42092),
            .in3(N__42248),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44920),
            .ce(N__41945),
            .sr(N__44120));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_10_LC_18_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_10_LC_18_12_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_10_LC_18_12_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_10_LC_18_12_1  (
            .in0(N__42244),
            .in1(N__42458),
            .in2(N__41528),
            .in3(N__42088),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44920),
            .ce(N__41945),
            .sr(N__44120));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_11_LC_18_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_11_LC_18_12_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_11_LC_18_12_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_11_LC_18_12_2  (
            .in0(N__42455),
            .in1(N__42245),
            .in2(N__42090),
            .in3(N__42534),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44920),
            .ce(N__41945),
            .sr(N__44120));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_16_LC_18_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_16_LC_18_12_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_16_LC_18_12_3 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_16_LC_18_12_3  (
            .in0(N__42494),
            .in1(N__42249),
            .in2(_gnd_net_),
            .in3(N__42085),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44920),
            .ce(N__41945),
            .sr(N__44120));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_13_LC_18_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_13_LC_18_12_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_13_LC_18_12_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_13_LC_18_12_4  (
            .in0(N__42456),
            .in1(N__42246),
            .in2(N__42091),
            .in3(N__42412),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44920),
            .ce(N__41945),
            .sr(N__44120));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_19_LC_18_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_19_LC_18_12_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_19_LC_18_12_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_19_LC_18_12_5  (
            .in0(N__42379),
            .in1(N__42251),
            .in2(_gnd_net_),
            .in3(N__42087),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44920),
            .ce(N__41945),
            .sr(N__44120));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_18_LC_18_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_18_LC_18_12_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_18_LC_18_12_6 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_18_LC_18_12_6  (
            .in0(N__42075),
            .in1(N__42344),
            .in2(_gnd_net_),
            .in3(N__42247),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44920),
            .ce(N__41945),
            .sr(N__44120));
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_17_LC_18_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_17_LC_18_12_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_time_esr_17_LC_18_12_7 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_esr_17_LC_18_12_7  (
            .in0(N__42305),
            .in1(N__42250),
            .in2(_gnd_net_),
            .in3(N__42086),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44920),
            .ce(N__41945),
            .sr(N__44120));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_18_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_18_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(N__41906),
            .in2(N__41861),
            .in3(N__41881),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_18_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_18_13_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_18_13_1  (
            .in0(N__41848),
            .in1(N__41837),
            .in2(N__41825),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_18_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_18_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_18_13_2  (
            .in0(_gnd_net_),
            .in1(N__42749),
            .in2(N__42782),
            .in3(N__42760),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_18_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_18_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(N__42743),
            .in2(N__42716),
            .in3(N__42727),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_18_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_18_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(N__42707),
            .in2(N__42683),
            .in3(N__42694),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_18_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_18_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__42674),
            .in2(N__42650),
            .in3(N__42661),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_18_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_18_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(N__42641),
            .in2(N__42617),
            .in3(N__42628),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_18_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_18_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_18_13_7  (
            .in0(N__42604),
            .in1(N__42593),
            .in2(N__42581),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_18_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_18_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__42572),
            .in2(N__42548),
            .in3(N__42559),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_18_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_18_14_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_18_14_1  (
            .in0(N__43030),
            .in1(N__43019),
            .in2(N__43010),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_18_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_18_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__43001),
            .in2(N__42980),
            .in3(N__42991),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_18_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_18_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__42971),
            .in2(N__42947),
            .in3(N__42958),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_18_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_18_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__42914),
            .in2(N__42938),
            .in3(N__42925),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_18_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_18_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__42905),
            .in2(N__42884),
            .in3(N__42895),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_18_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_18_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__42848),
            .in2(N__42875),
            .in3(N__42859),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_18_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_18_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_18_14_7  (
            .in0(N__42841),
            .in1(N__42830),
            .in2(N__42821),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_18_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_18_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__42788),
            .in2(N__42812),
            .in3(N__42799),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_18_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_18_15_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_18_15_1  (
            .in0(N__43252),
            .in1(N__43241),
            .in2(N__43232),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_18_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_18_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__43223),
            .in2(N__43202),
            .in3(N__43213),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43193),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NA_LC_18_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NA_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NA_LC_18_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NA_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__43189),
            .in2(_gnd_net_),
            .in3(N__43131),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNI62NAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_18_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_18_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__43085),
            .in2(N__43100),
            .in3(N__43681),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_18_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_18_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__43079),
            .in2(N__43070),
            .in3(N__43637),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_18_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_18_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__43061),
            .in2(N__43049),
            .in3(N__43607),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_18_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_18_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__43040),
            .in2(N__43406),
            .in3(N__43589),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_18_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_18_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__43385),
            .in2(N__43397),
            .in3(N__44546),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_18_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_18_16_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_18_16_5  (
            .in0(N__44528),
            .in1(N__43379),
            .in2(N__43367),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_18_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_18_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__43358),
            .in2(N__43346),
            .in3(N__44510),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_18_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_18_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(N__43337),
            .in2(N__43325),
            .in3(N__44492),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_18_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_18_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__43313),
            .in2(N__43298),
            .in3(N__44474),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_18_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_18_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__43289),
            .in2(N__43280),
            .in3(N__44456),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_18_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_18_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__43259),
            .in2(N__43271),
            .in3(N__44438),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_18_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_18_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__43571),
            .in2(N__43559),
            .in3(N__44420),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_18_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_18_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__43550),
            .in2(N__43538),
            .in3(N__44402),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_18_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_18_17_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_18_17_5  (
            .in0(N__45059),
            .in1(N__43529),
            .in2(N__43520),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_18_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_18_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__43511),
            .in2(N__43499),
            .in3(N__45041),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_18_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_18_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(N__43475),
            .in2(N__43490),
            .in3(N__45023),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_18_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_18_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__43469),
            .in2(N__43457),
            .in3(N__45005),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_18_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_18_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__43448),
            .in2(N__43439),
            .in3(N__44987),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_18_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_18_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__43427),
            .in2(N__43415),
            .in3(N__44966),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44384),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84AD_LC_18_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84AD_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84AD_LC_18_18_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84AD_LC_18_18_5  (
            .in0(N__43828),
            .in1(_gnd_net_),
            .in2(N__44367),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNI84ADZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_18_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_18_18_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__43827),
            .in2(_gnd_net_),
            .in3(N__44357),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIOA7T_0_1_LC_18_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIOA7T_0_1_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIOA7T_0_1_LC_18_18_7 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_RNIOA7T_0_1_LC_18_18_7  (
            .in0(N__44315),
            .in1(N__43868),
            .in2(N__43837),
            .in3(N__43784),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__43682),
            .in2(N__43646),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_18_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_18_19_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_18_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__43636),
            .in2(_gnd_net_),
            .in3(N__43622),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(N__44885),
            .ce(),
            .sr(N__44587));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_18_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_18_19_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_18_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__43606),
            .in2(N__43619),
            .in3(N__43592),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(N__44885),
            .ce(),
            .sr(N__44587));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_18_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_18_19_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_18_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__43588),
            .in2(_gnd_net_),
            .in3(N__43574),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(N__44885),
            .ce(),
            .sr(N__44587));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_18_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_18_19_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_18_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__44545),
            .in2(_gnd_net_),
            .in3(N__44531),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(N__44885),
            .ce(),
            .sr(N__44587));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_18_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_18_19_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_18_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__44527),
            .in2(_gnd_net_),
            .in3(N__44513),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(N__44885),
            .ce(),
            .sr(N__44587));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_18_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_18_19_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_18_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__44509),
            .in2(_gnd_net_),
            .in3(N__44495),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(N__44885),
            .ce(),
            .sr(N__44587));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_18_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_18_19_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_18_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__44491),
            .in2(_gnd_net_),
            .in3(N__44477),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(N__44885),
            .ce(),
            .sr(N__44587));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_18_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_18_20_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_18_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__44473),
            .in2(_gnd_net_),
            .in3(N__44459),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(N__44877),
            .ce(),
            .sr(N__44577));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_18_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_18_20_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_18_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__44455),
            .in2(_gnd_net_),
            .in3(N__44441),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(N__44877),
            .ce(),
            .sr(N__44577));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_18_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_18_20_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_18_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__44437),
            .in2(_gnd_net_),
            .in3(N__44423),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(N__44877),
            .ce(),
            .sr(N__44577));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_18_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_18_20_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_18_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__44419),
            .in2(_gnd_net_),
            .in3(N__44405),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(N__44877),
            .ce(),
            .sr(N__44577));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_18_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_18_20_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_18_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__44401),
            .in2(_gnd_net_),
            .in3(N__44387),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(N__44877),
            .ce(),
            .sr(N__44577));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_18_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_18_20_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_18_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__45058),
            .in2(_gnd_net_),
            .in3(N__45044),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(N__44877),
            .ce(),
            .sr(N__44577));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_18_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_18_20_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_18_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__45040),
            .in2(_gnd_net_),
            .in3(N__45026),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(N__44877),
            .ce(),
            .sr(N__44577));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_18_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_18_20_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_18_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_18_20_7  (
            .in0(_gnd_net_),
            .in1(N__45022),
            .in2(_gnd_net_),
            .in3(N__45008),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(N__44877),
            .ce(),
            .sr(N__44577));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_18_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_18_21_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_18_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__45004),
            .in2(_gnd_net_),
            .in3(N__44990),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_18_21_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(N__44871),
            .ce(),
            .sr(N__44576));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_18_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_18_21_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_18_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(N__44986),
            .in2(_gnd_net_),
            .in3(N__44972),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(N__44871),
            .ce(),
            .sr(N__44576));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_18_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_18_21_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_18_21_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(N__44965),
            .in2(_gnd_net_),
            .in3(N__44969),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__44871),
            .ce(),
            .sr(N__44576));
endmodule // MAIN
