// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 7 2025 00:28:56

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    start_stop,
    s2_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    input start_stop;
    output s2_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__49354;
    wire N__49353;
    wire N__49352;
    wire N__49343;
    wire N__49342;
    wire N__49341;
    wire N__49334;
    wire N__49333;
    wire N__49332;
    wire N__49325;
    wire N__49324;
    wire N__49323;
    wire N__49316;
    wire N__49315;
    wire N__49314;
    wire N__49307;
    wire N__49306;
    wire N__49305;
    wire N__49298;
    wire N__49297;
    wire N__49296;
    wire N__49289;
    wire N__49288;
    wire N__49287;
    wire N__49280;
    wire N__49279;
    wire N__49278;
    wire N__49271;
    wire N__49270;
    wire N__49269;
    wire N__49262;
    wire N__49261;
    wire N__49260;
    wire N__49253;
    wire N__49252;
    wire N__49251;
    wire N__49244;
    wire N__49243;
    wire N__49242;
    wire N__49225;
    wire N__49224;
    wire N__49221;
    wire N__49218;
    wire N__49213;
    wire N__49212;
    wire N__49211;
    wire N__49208;
    wire N__49205;
    wire N__49202;
    wire N__49197;
    wire N__49192;
    wire N__49189;
    wire N__49186;
    wire N__49183;
    wire N__49180;
    wire N__49177;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49165;
    wire N__49164;
    wire N__49163;
    wire N__49160;
    wire N__49157;
    wire N__49154;
    wire N__49149;
    wire N__49144;
    wire N__49141;
    wire N__49138;
    wire N__49135;
    wire N__49132;
    wire N__49129;
    wire N__49126;
    wire N__49125;
    wire N__49124;
    wire N__49121;
    wire N__49116;
    wire N__49115;
    wire N__49114;
    wire N__49111;
    wire N__49108;
    wire N__49105;
    wire N__49104;
    wire N__49103;
    wire N__49102;
    wire N__49101;
    wire N__49100;
    wire N__49099;
    wire N__49096;
    wire N__49095;
    wire N__49088;
    wire N__49077;
    wire N__49072;
    wire N__49069;
    wire N__49066;
    wire N__49063;
    wire N__49058;
    wire N__49053;
    wire N__49050;
    wire N__49047;
    wire N__49044;
    wire N__49039;
    wire N__49036;
    wire N__49035;
    wire N__49034;
    wire N__49033;
    wire N__49026;
    wire N__49023;
    wire N__49018;
    wire N__49015;
    wire N__49014;
    wire N__49013;
    wire N__49010;
    wire N__49005;
    wire N__49002;
    wire N__48999;
    wire N__48996;
    wire N__48993;
    wire N__48990;
    wire N__48985;
    wire N__48982;
    wire N__48979;
    wire N__48976;
    wire N__48973;
    wire N__48972;
    wire N__48971;
    wire N__48968;
    wire N__48965;
    wire N__48962;
    wire N__48959;
    wire N__48952;
    wire N__48949;
    wire N__48948;
    wire N__48945;
    wire N__48942;
    wire N__48939;
    wire N__48934;
    wire N__48933;
    wire N__48928;
    wire N__48925;
    wire N__48922;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48912;
    wire N__48911;
    wire N__48908;
    wire N__48905;
    wire N__48902;
    wire N__48895;
    wire N__48894;
    wire N__48891;
    wire N__48888;
    wire N__48885;
    wire N__48882;
    wire N__48879;
    wire N__48874;
    wire N__48873;
    wire N__48872;
    wire N__48871;
    wire N__48870;
    wire N__48869;
    wire N__48868;
    wire N__48867;
    wire N__48866;
    wire N__48865;
    wire N__48864;
    wire N__48863;
    wire N__48862;
    wire N__48861;
    wire N__48860;
    wire N__48859;
    wire N__48858;
    wire N__48857;
    wire N__48856;
    wire N__48855;
    wire N__48854;
    wire N__48853;
    wire N__48852;
    wire N__48851;
    wire N__48850;
    wire N__48849;
    wire N__48848;
    wire N__48847;
    wire N__48846;
    wire N__48845;
    wire N__48844;
    wire N__48843;
    wire N__48842;
    wire N__48841;
    wire N__48840;
    wire N__48839;
    wire N__48838;
    wire N__48837;
    wire N__48836;
    wire N__48835;
    wire N__48834;
    wire N__48833;
    wire N__48832;
    wire N__48831;
    wire N__48830;
    wire N__48829;
    wire N__48828;
    wire N__48827;
    wire N__48826;
    wire N__48825;
    wire N__48824;
    wire N__48823;
    wire N__48822;
    wire N__48821;
    wire N__48820;
    wire N__48819;
    wire N__48818;
    wire N__48817;
    wire N__48816;
    wire N__48815;
    wire N__48814;
    wire N__48813;
    wire N__48812;
    wire N__48811;
    wire N__48810;
    wire N__48809;
    wire N__48808;
    wire N__48807;
    wire N__48806;
    wire N__48805;
    wire N__48804;
    wire N__48803;
    wire N__48802;
    wire N__48801;
    wire N__48800;
    wire N__48799;
    wire N__48798;
    wire N__48797;
    wire N__48796;
    wire N__48795;
    wire N__48794;
    wire N__48793;
    wire N__48792;
    wire N__48791;
    wire N__48790;
    wire N__48789;
    wire N__48788;
    wire N__48787;
    wire N__48786;
    wire N__48785;
    wire N__48784;
    wire N__48783;
    wire N__48782;
    wire N__48781;
    wire N__48780;
    wire N__48779;
    wire N__48778;
    wire N__48777;
    wire N__48776;
    wire N__48775;
    wire N__48774;
    wire N__48773;
    wire N__48772;
    wire N__48771;
    wire N__48770;
    wire N__48769;
    wire N__48768;
    wire N__48767;
    wire N__48766;
    wire N__48765;
    wire N__48764;
    wire N__48763;
    wire N__48762;
    wire N__48761;
    wire N__48760;
    wire N__48759;
    wire N__48758;
    wire N__48757;
    wire N__48756;
    wire N__48755;
    wire N__48754;
    wire N__48753;
    wire N__48752;
    wire N__48751;
    wire N__48750;
    wire N__48749;
    wire N__48748;
    wire N__48747;
    wire N__48746;
    wire N__48745;
    wire N__48744;
    wire N__48743;
    wire N__48742;
    wire N__48741;
    wire N__48740;
    wire N__48739;
    wire N__48738;
    wire N__48737;
    wire N__48736;
    wire N__48735;
    wire N__48734;
    wire N__48733;
    wire N__48732;
    wire N__48731;
    wire N__48730;
    wire N__48729;
    wire N__48728;
    wire N__48727;
    wire N__48726;
    wire N__48725;
    wire N__48724;
    wire N__48723;
    wire N__48722;
    wire N__48721;
    wire N__48720;
    wire N__48719;
    wire N__48718;
    wire N__48717;
    wire N__48716;
    wire N__48715;
    wire N__48714;
    wire N__48713;
    wire N__48712;
    wire N__48711;
    wire N__48710;
    wire N__48709;
    wire N__48708;
    wire N__48707;
    wire N__48706;
    wire N__48705;
    wire N__48704;
    wire N__48703;
    wire N__48702;
    wire N__48701;
    wire N__48700;
    wire N__48349;
    wire N__48346;
    wire N__48345;
    wire N__48344;
    wire N__48343;
    wire N__48340;
    wire N__48339;
    wire N__48338;
    wire N__48335;
    wire N__48332;
    wire N__48329;
    wire N__48326;
    wire N__48323;
    wire N__48320;
    wire N__48317;
    wire N__48312;
    wire N__48309;
    wire N__48306;
    wire N__48303;
    wire N__48300;
    wire N__48297;
    wire N__48292;
    wire N__48289;
    wire N__48280;
    wire N__48279;
    wire N__48278;
    wire N__48277;
    wire N__48276;
    wire N__48275;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48263;
    wire N__48260;
    wire N__48257;
    wire N__48254;
    wire N__48251;
    wire N__48248;
    wire N__48245;
    wire N__48242;
    wire N__48241;
    wire N__48240;
    wire N__48239;
    wire N__48238;
    wire N__48237;
    wire N__48236;
    wire N__48235;
    wire N__48234;
    wire N__48233;
    wire N__48232;
    wire N__48231;
    wire N__48230;
    wire N__48229;
    wire N__48228;
    wire N__48227;
    wire N__48226;
    wire N__48225;
    wire N__48224;
    wire N__48223;
    wire N__48222;
    wire N__48221;
    wire N__48220;
    wire N__48219;
    wire N__48218;
    wire N__48217;
    wire N__48216;
    wire N__48215;
    wire N__48214;
    wire N__48213;
    wire N__48212;
    wire N__48211;
    wire N__48210;
    wire N__48209;
    wire N__48208;
    wire N__48207;
    wire N__48206;
    wire N__48205;
    wire N__48204;
    wire N__48203;
    wire N__48202;
    wire N__48201;
    wire N__48200;
    wire N__48199;
    wire N__48198;
    wire N__48197;
    wire N__48196;
    wire N__48195;
    wire N__48194;
    wire N__48193;
    wire N__48192;
    wire N__48191;
    wire N__48190;
    wire N__48189;
    wire N__48188;
    wire N__48187;
    wire N__48186;
    wire N__48185;
    wire N__48184;
    wire N__48183;
    wire N__48182;
    wire N__48181;
    wire N__48180;
    wire N__48179;
    wire N__48178;
    wire N__48177;
    wire N__48176;
    wire N__48175;
    wire N__48174;
    wire N__48173;
    wire N__48172;
    wire N__48171;
    wire N__48170;
    wire N__48167;
    wire N__48166;
    wire N__48165;
    wire N__48164;
    wire N__48163;
    wire N__48162;
    wire N__48161;
    wire N__48160;
    wire N__48159;
    wire N__48158;
    wire N__48157;
    wire N__48156;
    wire N__48155;
    wire N__48154;
    wire N__48153;
    wire N__48152;
    wire N__48151;
    wire N__48150;
    wire N__48149;
    wire N__48148;
    wire N__48147;
    wire N__48146;
    wire N__48145;
    wire N__48144;
    wire N__48143;
    wire N__48142;
    wire N__48141;
    wire N__48140;
    wire N__48139;
    wire N__48138;
    wire N__48137;
    wire N__48136;
    wire N__48135;
    wire N__48134;
    wire N__48133;
    wire N__48132;
    wire N__48131;
    wire N__48130;
    wire N__48129;
    wire N__48128;
    wire N__48127;
    wire N__48126;
    wire N__48125;
    wire N__48124;
    wire N__48123;
    wire N__48122;
    wire N__48121;
    wire N__48120;
    wire N__48119;
    wire N__48118;
    wire N__48117;
    wire N__48114;
    wire N__48113;
    wire N__48112;
    wire N__48111;
    wire N__48110;
    wire N__48109;
    wire N__48108;
    wire N__48107;
    wire N__48106;
    wire N__48105;
    wire N__48104;
    wire N__48103;
    wire N__48102;
    wire N__48101;
    wire N__48100;
    wire N__48099;
    wire N__48098;
    wire N__48097;
    wire N__48096;
    wire N__48095;
    wire N__48094;
    wire N__48093;
    wire N__48092;
    wire N__48091;
    wire N__48090;
    wire N__48089;
    wire N__48088;
    wire N__47779;
    wire N__47776;
    wire N__47773;
    wire N__47772;
    wire N__47771;
    wire N__47768;
    wire N__47765;
    wire N__47762;
    wire N__47757;
    wire N__47752;
    wire N__47749;
    wire N__47746;
    wire N__47743;
    wire N__47740;
    wire N__47737;
    wire N__47736;
    wire N__47735;
    wire N__47732;
    wire N__47729;
    wire N__47726;
    wire N__47721;
    wire N__47716;
    wire N__47713;
    wire N__47710;
    wire N__47707;
    wire N__47704;
    wire N__47701;
    wire N__47700;
    wire N__47699;
    wire N__47696;
    wire N__47691;
    wire N__47686;
    wire N__47683;
    wire N__47680;
    wire N__47677;
    wire N__47674;
    wire N__47671;
    wire N__47670;
    wire N__47669;
    wire N__47666;
    wire N__47661;
    wire N__47656;
    wire N__47653;
    wire N__47650;
    wire N__47647;
    wire N__47644;
    wire N__47641;
    wire N__47638;
    wire N__47637;
    wire N__47636;
    wire N__47633;
    wire N__47630;
    wire N__47627;
    wire N__47622;
    wire N__47617;
    wire N__47614;
    wire N__47611;
    wire N__47608;
    wire N__47605;
    wire N__47602;
    wire N__47601;
    wire N__47600;
    wire N__47597;
    wire N__47594;
    wire N__47591;
    wire N__47586;
    wire N__47581;
    wire N__47578;
    wire N__47575;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47565;
    wire N__47564;
    wire N__47561;
    wire N__47558;
    wire N__47555;
    wire N__47548;
    wire N__47545;
    wire N__47542;
    wire N__47539;
    wire N__47536;
    wire N__47535;
    wire N__47534;
    wire N__47531;
    wire N__47528;
    wire N__47525;
    wire N__47518;
    wire N__47515;
    wire N__47512;
    wire N__47509;
    wire N__47506;
    wire N__47503;
    wire N__47502;
    wire N__47501;
    wire N__47498;
    wire N__47495;
    wire N__47492;
    wire N__47487;
    wire N__47482;
    wire N__47481;
    wire N__47478;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47452;
    wire N__47449;
    wire N__47448;
    wire N__47447;
    wire N__47444;
    wire N__47441;
    wire N__47438;
    wire N__47433;
    wire N__47428;
    wire N__47427;
    wire N__47426;
    wire N__47425;
    wire N__47422;
    wire N__47419;
    wire N__47418;
    wire N__47413;
    wire N__47410;
    wire N__47407;
    wire N__47404;
    wire N__47399;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47383;
    wire N__47380;
    wire N__47379;
    wire N__47378;
    wire N__47375;
    wire N__47370;
    wire N__47365;
    wire N__47364;
    wire N__47363;
    wire N__47362;
    wire N__47361;
    wire N__47358;
    wire N__47355;
    wire N__47354;
    wire N__47351;
    wire N__47348;
    wire N__47345;
    wire N__47342;
    wire N__47339;
    wire N__47336;
    wire N__47333;
    wire N__47328;
    wire N__47319;
    wire N__47314;
    wire N__47311;
    wire N__47308;
    wire N__47307;
    wire N__47306;
    wire N__47303;
    wire N__47298;
    wire N__47293;
    wire N__47290;
    wire N__47289;
    wire N__47286;
    wire N__47283;
    wire N__47282;
    wire N__47279;
    wire N__47276;
    wire N__47273;
    wire N__47268;
    wire N__47265;
    wire N__47262;
    wire N__47257;
    wire N__47254;
    wire N__47253;
    wire N__47252;
    wire N__47249;
    wire N__47246;
    wire N__47243;
    wire N__47238;
    wire N__47233;
    wire N__47232;
    wire N__47229;
    wire N__47228;
    wire N__47225;
    wire N__47222;
    wire N__47219;
    wire N__47216;
    wire N__47211;
    wire N__47208;
    wire N__47203;
    wire N__47200;
    wire N__47199;
    wire N__47198;
    wire N__47195;
    wire N__47192;
    wire N__47189;
    wire N__47184;
    wire N__47179;
    wire N__47176;
    wire N__47173;
    wire N__47172;
    wire N__47169;
    wire N__47168;
    wire N__47165;
    wire N__47162;
    wire N__47159;
    wire N__47156;
    wire N__47151;
    wire N__47148;
    wire N__47143;
    wire N__47140;
    wire N__47139;
    wire N__47138;
    wire N__47135;
    wire N__47132;
    wire N__47129;
    wire N__47122;
    wire N__47119;
    wire N__47118;
    wire N__47117;
    wire N__47114;
    wire N__47111;
    wire N__47108;
    wire N__47105;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47087;
    wire N__47082;
    wire N__47077;
    wire N__47074;
    wire N__47073;
    wire N__47072;
    wire N__47069;
    wire N__47066;
    wire N__47063;
    wire N__47056;
    wire N__47053;
    wire N__47050;
    wire N__47047;
    wire N__47044;
    wire N__47041;
    wire N__47040;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47030;
    wire N__47025;
    wire N__47020;
    wire N__47019;
    wire N__47018;
    wire N__47015;
    wire N__47012;
    wire N__47009;
    wire N__47002;
    wire N__46999;
    wire N__46996;
    wire N__46993;
    wire N__46992;
    wire N__46991;
    wire N__46988;
    wire N__46983;
    wire N__46978;
    wire N__46975;
    wire N__46972;
    wire N__46971;
    wire N__46970;
    wire N__46967;
    wire N__46964;
    wire N__46961;
    wire N__46958;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46942;
    wire N__46939;
    wire N__46938;
    wire N__46937;
    wire N__46934;
    wire N__46929;
    wire N__46924;
    wire N__46921;
    wire N__46918;
    wire N__46917;
    wire N__46916;
    wire N__46913;
    wire N__46910;
    wire N__46907;
    wire N__46904;
    wire N__46899;
    wire N__46896;
    wire N__46893;
    wire N__46888;
    wire N__46885;
    wire N__46884;
    wire N__46883;
    wire N__46880;
    wire N__46877;
    wire N__46874;
    wire N__46869;
    wire N__46864;
    wire N__46861;
    wire N__46860;
    wire N__46857;
    wire N__46856;
    wire N__46853;
    wire N__46852;
    wire N__46849;
    wire N__46846;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46834;
    wire N__46831;
    wire N__46828;
    wire N__46825;
    wire N__46818;
    wire N__46813;
    wire N__46810;
    wire N__46809;
    wire N__46808;
    wire N__46805;
    wire N__46802;
    wire N__46799;
    wire N__46794;
    wire N__46789;
    wire N__46788;
    wire N__46785;
    wire N__46782;
    wire N__46779;
    wire N__46776;
    wire N__46773;
    wire N__46770;
    wire N__46765;
    wire N__46762;
    wire N__46761;
    wire N__46760;
    wire N__46757;
    wire N__46754;
    wire N__46751;
    wire N__46744;
    wire N__46741;
    wire N__46740;
    wire N__46737;
    wire N__46734;
    wire N__46731;
    wire N__46728;
    wire N__46725;
    wire N__46722;
    wire N__46717;
    wire N__46714;
    wire N__46713;
    wire N__46712;
    wire N__46709;
    wire N__46706;
    wire N__46703;
    wire N__46696;
    wire N__46693;
    wire N__46692;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46674;
    wire N__46669;
    wire N__46666;
    wire N__46663;
    wire N__46660;
    wire N__46657;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46645;
    wire N__46644;
    wire N__46643;
    wire N__46642;
    wire N__46641;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46629;
    wire N__46628;
    wire N__46625;
    wire N__46622;
    wire N__46619;
    wire N__46616;
    wire N__46613;
    wire N__46610;
    wire N__46607;
    wire N__46604;
    wire N__46601;
    wire N__46598;
    wire N__46593;
    wire N__46590;
    wire N__46583;
    wire N__46580;
    wire N__46577;
    wire N__46570;
    wire N__46569;
    wire N__46566;
    wire N__46563;
    wire N__46560;
    wire N__46559;
    wire N__46556;
    wire N__46553;
    wire N__46550;
    wire N__46547;
    wire N__46544;
    wire N__46541;
    wire N__46538;
    wire N__46531;
    wire N__46528;
    wire N__46527;
    wire N__46526;
    wire N__46523;
    wire N__46520;
    wire N__46517;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46507;
    wire N__46504;
    wire N__46503;
    wire N__46502;
    wire N__46501;
    wire N__46498;
    wire N__46491;
    wire N__46486;
    wire N__46483;
    wire N__46474;
    wire N__46473;
    wire N__46470;
    wire N__46467;
    wire N__46464;
    wire N__46463;
    wire N__46460;
    wire N__46457;
    wire N__46454;
    wire N__46447;
    wire N__46446;
    wire N__46443;
    wire N__46440;
    wire N__46439;
    wire N__46438;
    wire N__46433;
    wire N__46430;
    wire N__46427;
    wire N__46424;
    wire N__46419;
    wire N__46418;
    wire N__46417;
    wire N__46416;
    wire N__46415;
    wire N__46412;
    wire N__46409;
    wire N__46402;
    wire N__46399;
    wire N__46390;
    wire N__46387;
    wire N__46386;
    wire N__46383;
    wire N__46382;
    wire N__46379;
    wire N__46376;
    wire N__46373;
    wire N__46370;
    wire N__46367;
    wire N__46364;
    wire N__46361;
    wire N__46354;
    wire N__46351;
    wire N__46350;
    wire N__46349;
    wire N__46346;
    wire N__46345;
    wire N__46344;
    wire N__46343;
    wire N__46340;
    wire N__46337;
    wire N__46334;
    wire N__46331;
    wire N__46328;
    wire N__46325;
    wire N__46322;
    wire N__46319;
    wire N__46314;
    wire N__46311;
    wire N__46308;
    wire N__46305;
    wire N__46302;
    wire N__46297;
    wire N__46294;
    wire N__46285;
    wire N__46284;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46270;
    wire N__46269;
    wire N__46268;
    wire N__46265;
    wire N__46262;
    wire N__46259;
    wire N__46252;
    wire N__46251;
    wire N__46250;
    wire N__46245;
    wire N__46242;
    wire N__46241;
    wire N__46240;
    wire N__46239;
    wire N__46238;
    wire N__46235;
    wire N__46232;
    wire N__46229;
    wire N__46226;
    wire N__46221;
    wire N__46220;
    wire N__46219;
    wire N__46216;
    wire N__46213;
    wire N__46210;
    wire N__46205;
    wire N__46202;
    wire N__46199;
    wire N__46196;
    wire N__46191;
    wire N__46184;
    wire N__46177;
    wire N__46174;
    wire N__46171;
    wire N__46168;
    wire N__46167;
    wire N__46166;
    wire N__46165;
    wire N__46162;
    wire N__46159;
    wire N__46156;
    wire N__46155;
    wire N__46154;
    wire N__46153;
    wire N__46148;
    wire N__46145;
    wire N__46142;
    wire N__46139;
    wire N__46136;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46108;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46094;
    wire N__46087;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46079;
    wire N__46076;
    wire N__46073;
    wire N__46070;
    wire N__46065;
    wire N__46062;
    wire N__46059;
    wire N__46056;
    wire N__46051;
    wire N__46048;
    wire N__46047;
    wire N__46046;
    wire N__46043;
    wire N__46040;
    wire N__46037;
    wire N__46030;
    wire N__46029;
    wire N__46028;
    wire N__46025;
    wire N__46022;
    wire N__46019;
    wire N__46016;
    wire N__46013;
    wire N__46010;
    wire N__46007;
    wire N__46004;
    wire N__45997;
    wire N__45994;
    wire N__45993;
    wire N__45992;
    wire N__45989;
    wire N__45986;
    wire N__45983;
    wire N__45978;
    wire N__45973;
    wire N__45970;
    wire N__45969;
    wire N__45968;
    wire N__45965;
    wire N__45962;
    wire N__45959;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45940;
    wire N__45937;
    wire N__45934;
    wire N__45931;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45923;
    wire N__45922;
    wire N__45917;
    wire N__45914;
    wire N__45911;
    wire N__45904;
    wire N__45901;
    wire N__45900;
    wire N__45897;
    wire N__45896;
    wire N__45893;
    wire N__45890;
    wire N__45887;
    wire N__45884;
    wire N__45877;
    wire N__45874;
    wire N__45873;
    wire N__45872;
    wire N__45871;
    wire N__45870;
    wire N__45867;
    wire N__45862;
    wire N__45861;
    wire N__45858;
    wire N__45855;
    wire N__45852;
    wire N__45849;
    wire N__45846;
    wire N__45841;
    wire N__45838;
    wire N__45833;
    wire N__45830;
    wire N__45823;
    wire N__45822;
    wire N__45819;
    wire N__45818;
    wire N__45815;
    wire N__45812;
    wire N__45809;
    wire N__45802;
    wire N__45799;
    wire N__45796;
    wire N__45793;
    wire N__45790;
    wire N__45787;
    wire N__45784;
    wire N__45781;
    wire N__45778;
    wire N__45775;
    wire N__45774;
    wire N__45771;
    wire N__45768;
    wire N__45763;
    wire N__45760;
    wire N__45759;
    wire N__45758;
    wire N__45757;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45747;
    wire N__45744;
    wire N__45741;
    wire N__45736;
    wire N__45727;
    wire N__45726;
    wire N__45723;
    wire N__45720;
    wire N__45715;
    wire N__45714;
    wire N__45713;
    wire N__45710;
    wire N__45707;
    wire N__45704;
    wire N__45701;
    wire N__45696;
    wire N__45691;
    wire N__45688;
    wire N__45685;
    wire N__45684;
    wire N__45681;
    wire N__45678;
    wire N__45673;
    wire N__45670;
    wire N__45667;
    wire N__45666;
    wire N__45663;
    wire N__45660;
    wire N__45655;
    wire N__45654;
    wire N__45653;
    wire N__45652;
    wire N__45651;
    wire N__45650;
    wire N__45649;
    wire N__45648;
    wire N__45647;
    wire N__45644;
    wire N__45643;
    wire N__45640;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45630;
    wire N__45629;
    wire N__45628;
    wire N__45627;
    wire N__45626;
    wire N__45625;
    wire N__45622;
    wire N__45621;
    wire N__45620;
    wire N__45619;
    wire N__45618;
    wire N__45615;
    wire N__45612;
    wire N__45609;
    wire N__45604;
    wire N__45603;
    wire N__45586;
    wire N__45581;
    wire N__45564;
    wire N__45561;
    wire N__45560;
    wire N__45557;
    wire N__45556;
    wire N__45555;
    wire N__45552;
    wire N__45547;
    wire N__45544;
    wire N__45541;
    wire N__45538;
    wire N__45533;
    wire N__45528;
    wire N__45523;
    wire N__45514;
    wire N__45513;
    wire N__45512;
    wire N__45511;
    wire N__45510;
    wire N__45509;
    wire N__45508;
    wire N__45507;
    wire N__45506;
    wire N__45505;
    wire N__45504;
    wire N__45503;
    wire N__45502;
    wire N__45501;
    wire N__45500;
    wire N__45499;
    wire N__45498;
    wire N__45481;
    wire N__45464;
    wire N__45461;
    wire N__45460;
    wire N__45459;
    wire N__45458;
    wire N__45457;
    wire N__45456;
    wire N__45451;
    wire N__45446;
    wire N__45443;
    wire N__45438;
    wire N__45435;
    wire N__45434;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45424;
    wire N__45419;
    wire N__45414;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45394;
    wire N__45393;
    wire N__45392;
    wire N__45391;
    wire N__45390;
    wire N__45389;
    wire N__45388;
    wire N__45387;
    wire N__45386;
    wire N__45385;
    wire N__45384;
    wire N__45383;
    wire N__45382;
    wire N__45381;
    wire N__45380;
    wire N__45379;
    wire N__45378;
    wire N__45377;
    wire N__45376;
    wire N__45375;
    wire N__45374;
    wire N__45371;
    wire N__45366;
    wire N__45365;
    wire N__45362;
    wire N__45361;
    wire N__45344;
    wire N__45327;
    wire N__45326;
    wire N__45323;
    wire N__45320;
    wire N__45317;
    wire N__45314;
    wire N__45309;
    wire N__45304;
    wire N__45301;
    wire N__45292;
    wire N__45287;
    wire N__45284;
    wire N__45281;
    wire N__45274;
    wire N__45271;
    wire N__45270;
    wire N__45267;
    wire N__45264;
    wire N__45263;
    wire N__45260;
    wire N__45257;
    wire N__45254;
    wire N__45253;
    wire N__45250;
    wire N__45245;
    wire N__45242;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45226;
    wire N__45223;
    wire N__45220;
    wire N__45219;
    wire N__45216;
    wire N__45213;
    wire N__45212;
    wire N__45211;
    wire N__45206;
    wire N__45203;
    wire N__45200;
    wire N__45197;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45176;
    wire N__45173;
    wire N__45166;
    wire N__45165;
    wire N__45164;
    wire N__45161;
    wire N__45158;
    wire N__45157;
    wire N__45156;
    wire N__45155;
    wire N__45154;
    wire N__45153;
    wire N__45142;
    wire N__45141;
    wire N__45138;
    wire N__45137;
    wire N__45136;
    wire N__45135;
    wire N__45134;
    wire N__45133;
    wire N__45132;
    wire N__45131;
    wire N__45128;
    wire N__45125;
    wire N__45122;
    wire N__45119;
    wire N__45116;
    wire N__45113;
    wire N__45106;
    wire N__45099;
    wire N__45094;
    wire N__45089;
    wire N__45084;
    wire N__45079;
    wire N__45076;
    wire N__45071;
    wire N__45068;
    wire N__45065;
    wire N__45058;
    wire N__45057;
    wire N__45054;
    wire N__45053;
    wire N__45052;
    wire N__45049;
    wire N__45044;
    wire N__45041;
    wire N__45038;
    wire N__45035;
    wire N__45034;
    wire N__45033;
    wire N__45030;
    wire N__45027;
    wire N__45024;
    wire N__45019;
    wire N__45014;
    wire N__45007;
    wire N__45006;
    wire N__45005;
    wire N__45004;
    wire N__44995;
    wire N__44994;
    wire N__44993;
    wire N__44990;
    wire N__44987;
    wire N__44984;
    wire N__44979;
    wire N__44976;
    wire N__44975;
    wire N__44974;
    wire N__44973;
    wire N__44972;
    wire N__44969;
    wire N__44966;
    wire N__44963;
    wire N__44956;
    wire N__44953;
    wire N__44944;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44932;
    wire N__44929;
    wire N__44926;
    wire N__44923;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44913;
    wire N__44910;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44896;
    wire N__44893;
    wire N__44890;
    wire N__44889;
    wire N__44886;
    wire N__44883;
    wire N__44878;
    wire N__44875;
    wire N__44872;
    wire N__44869;
    wire N__44866;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44854;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44839;
    wire N__44836;
    wire N__44833;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44823;
    wire N__44822;
    wire N__44821;
    wire N__44818;
    wire N__44811;
    wire N__44806;
    wire N__44805;
    wire N__44802;
    wire N__44799;
    wire N__44798;
    wire N__44795;
    wire N__44790;
    wire N__44785;
    wire N__44782;
    wire N__44779;
    wire N__44776;
    wire N__44773;
    wire N__44770;
    wire N__44767;
    wire N__44766;
    wire N__44763;
    wire N__44760;
    wire N__44757;
    wire N__44754;
    wire N__44749;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44737;
    wire N__44734;
    wire N__44731;
    wire N__44728;
    wire N__44725;
    wire N__44722;
    wire N__44721;
    wire N__44718;
    wire N__44715;
    wire N__44710;
    wire N__44707;
    wire N__44704;
    wire N__44701;
    wire N__44698;
    wire N__44695;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44683;
    wire N__44680;
    wire N__44677;
    wire N__44674;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44662;
    wire N__44659;
    wire N__44656;
    wire N__44653;
    wire N__44652;
    wire N__44649;
    wire N__44646;
    wire N__44641;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44620;
    wire N__44617;
    wire N__44614;
    wire N__44611;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44589;
    wire N__44586;
    wire N__44583;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44569;
    wire N__44568;
    wire N__44567;
    wire N__44566;
    wire N__44565;
    wire N__44564;
    wire N__44563;
    wire N__44562;
    wire N__44561;
    wire N__44560;
    wire N__44559;
    wire N__44558;
    wire N__44557;
    wire N__44556;
    wire N__44555;
    wire N__44554;
    wire N__44553;
    wire N__44552;
    wire N__44551;
    wire N__44550;
    wire N__44549;
    wire N__44548;
    wire N__44547;
    wire N__44546;
    wire N__44545;
    wire N__44544;
    wire N__44543;
    wire N__44542;
    wire N__44541;
    wire N__44540;
    wire N__44531;
    wire N__44526;
    wire N__44517;
    wire N__44508;
    wire N__44499;
    wire N__44490;
    wire N__44481;
    wire N__44472;
    wire N__44461;
    wire N__44458;
    wire N__44451;
    wire N__44446;
    wire N__44443;
    wire N__44442;
    wire N__44441;
    wire N__44440;
    wire N__44437;
    wire N__44434;
    wire N__44431;
    wire N__44428;
    wire N__44425;
    wire N__44422;
    wire N__44417;
    wire N__44410;
    wire N__44407;
    wire N__44404;
    wire N__44401;
    wire N__44398;
    wire N__44397;
    wire N__44394;
    wire N__44393;
    wire N__44390;
    wire N__44387;
    wire N__44384;
    wire N__44377;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44353;
    wire N__44350;
    wire N__44347;
    wire N__44344;
    wire N__44341;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44329;
    wire N__44326;
    wire N__44323;
    wire N__44320;
    wire N__44319;
    wire N__44316;
    wire N__44313;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44296;
    wire N__44293;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44281;
    wire N__44278;
    wire N__44275;
    wire N__44272;
    wire N__44269;
    wire N__44268;
    wire N__44265;
    wire N__44262;
    wire N__44257;
    wire N__44254;
    wire N__44251;
    wire N__44248;
    wire N__44245;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44218;
    wire N__44215;
    wire N__44212;
    wire N__44209;
    wire N__44206;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44179;
    wire N__44176;
    wire N__44173;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44161;
    wire N__44158;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44143;
    wire N__44140;
    wire N__44137;
    wire N__44134;
    wire N__44131;
    wire N__44128;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44116;
    wire N__44115;
    wire N__44114;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44098;
    wire N__44097;
    wire N__44094;
    wire N__44091;
    wire N__44086;
    wire N__44083;
    wire N__44082;
    wire N__44081;
    wire N__44080;
    wire N__44079;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44059;
    wire N__44058;
    wire N__44057;
    wire N__44056;
    wire N__44053;
    wire N__44050;
    wire N__44045;
    wire N__44042;
    wire N__44035;
    wire N__44032;
    wire N__44029;
    wire N__44026;
    wire N__44023;
    wire N__44020;
    wire N__44017;
    wire N__44014;
    wire N__44011;
    wire N__44010;
    wire N__44007;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43987;
    wire N__43986;
    wire N__43985;
    wire N__43982;
    wire N__43981;
    wire N__43976;
    wire N__43973;
    wire N__43970;
    wire N__43967;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43951;
    wire N__43948;
    wire N__43947;
    wire N__43944;
    wire N__43943;
    wire N__43940;
    wire N__43937;
    wire N__43934;
    wire N__43931;
    wire N__43924;
    wire N__43921;
    wire N__43918;
    wire N__43915;
    wire N__43912;
    wire N__43909;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43878;
    wire N__43877;
    wire N__43876;
    wire N__43873;
    wire N__43870;
    wire N__43865;
    wire N__43860;
    wire N__43857;
    wire N__43852;
    wire N__43851;
    wire N__43848;
    wire N__43845;
    wire N__43840;
    wire N__43837;
    wire N__43836;
    wire N__43833;
    wire N__43830;
    wire N__43827;
    wire N__43826;
    wire N__43821;
    wire N__43818;
    wire N__43815;
    wire N__43810;
    wire N__43807;
    wire N__43806;
    wire N__43803;
    wire N__43800;
    wire N__43799;
    wire N__43794;
    wire N__43791;
    wire N__43788;
    wire N__43783;
    wire N__43780;
    wire N__43777;
    wire N__43776;
    wire N__43773;
    wire N__43772;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43758;
    wire N__43753;
    wire N__43750;
    wire N__43747;
    wire N__43744;
    wire N__43743;
    wire N__43740;
    wire N__43737;
    wire N__43734;
    wire N__43729;
    wire N__43726;
    wire N__43725;
    wire N__43724;
    wire N__43723;
    wire N__43722;
    wire N__43721;
    wire N__43720;
    wire N__43719;
    wire N__43718;
    wire N__43717;
    wire N__43716;
    wire N__43715;
    wire N__43714;
    wire N__43713;
    wire N__43712;
    wire N__43711;
    wire N__43710;
    wire N__43709;
    wire N__43708;
    wire N__43707;
    wire N__43706;
    wire N__43705;
    wire N__43704;
    wire N__43703;
    wire N__43694;
    wire N__43685;
    wire N__43676;
    wire N__43667;
    wire N__43658;
    wire N__43649;
    wire N__43648;
    wire N__43647;
    wire N__43646;
    wire N__43645;
    wire N__43644;
    wire N__43643;
    wire N__43634;
    wire N__43629;
    wire N__43624;
    wire N__43615;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43590;
    wire N__43587;
    wire N__43584;
    wire N__43581;
    wire N__43576;
    wire N__43573;
    wire N__43572;
    wire N__43571;
    wire N__43568;
    wire N__43565;
    wire N__43562;
    wire N__43561;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43545;
    wire N__43542;
    wire N__43539;
    wire N__43536;
    wire N__43531;
    wire N__43528;
    wire N__43525;
    wire N__43522;
    wire N__43519;
    wire N__43516;
    wire N__43513;
    wire N__43510;
    wire N__43507;
    wire N__43504;
    wire N__43501;
    wire N__43500;
    wire N__43499;
    wire N__43498;
    wire N__43497;
    wire N__43496;
    wire N__43495;
    wire N__43494;
    wire N__43493;
    wire N__43490;
    wire N__43483;
    wire N__43474;
    wire N__43473;
    wire N__43472;
    wire N__43471;
    wire N__43470;
    wire N__43469;
    wire N__43468;
    wire N__43467;
    wire N__43466;
    wire N__43465;
    wire N__43464;
    wire N__43463;
    wire N__43462;
    wire N__43461;
    wire N__43460;
    wire N__43459;
    wire N__43458;
    wire N__43457;
    wire N__43456;
    wire N__43455;
    wire N__43454;
    wire N__43453;
    wire N__43452;
    wire N__43451;
    wire N__43450;
    wire N__43449;
    wire N__43446;
    wire N__43443;
    wire N__43438;
    wire N__43435;
    wire N__43434;
    wire N__43431;
    wire N__43430;
    wire N__43427;
    wire N__43424;
    wire N__43421;
    wire N__43418;
    wire N__43415;
    wire N__43412;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43394;
    wire N__43391;
    wire N__43388;
    wire N__43385;
    wire N__43382;
    wire N__43379;
    wire N__43376;
    wire N__43373;
    wire N__43370;
    wire N__43367;
    wire N__43364;
    wire N__43363;
    wire N__43362;
    wire N__43361;
    wire N__43360;
    wire N__43359;
    wire N__43358;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43350;
    wire N__43345;
    wire N__43342;
    wire N__43341;
    wire N__43340;
    wire N__43339;
    wire N__43338;
    wire N__43337;
    wire N__43336;
    wire N__43335;
    wire N__43334;
    wire N__43331;
    wire N__43326;
    wire N__43317;
    wire N__43308;
    wire N__43301;
    wire N__43294;
    wire N__43285;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43267;
    wire N__43264;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43250;
    wire N__43247;
    wire N__43242;
    wire N__43235;
    wire N__43226;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43212;
    wire N__43203;
    wire N__43196;
    wire N__43187;
    wire N__43182;
    wire N__43179;
    wire N__43174;
    wire N__43171;
    wire N__43166;
    wire N__43163;
    wire N__43156;
    wire N__43153;
    wire N__43148;
    wire N__43145;
    wire N__43142;
    wire N__43137;
    wire N__43134;
    wire N__43131;
    wire N__43126;
    wire N__43123;
    wire N__43114;
    wire N__43113;
    wire N__43110;
    wire N__43107;
    wire N__43104;
    wire N__43103;
    wire N__43098;
    wire N__43095;
    wire N__43092;
    wire N__43087;
    wire N__43084;
    wire N__43083;
    wire N__43080;
    wire N__43077;
    wire N__43074;
    wire N__43073;
    wire N__43068;
    wire N__43065;
    wire N__43062;
    wire N__43057;
    wire N__43054;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43046;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43023;
    wire N__43020;
    wire N__43019;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43005;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42993;
    wire N__42988;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42973;
    wire N__42970;
    wire N__42969;
    wire N__42966;
    wire N__42963;
    wire N__42958;
    wire N__42957;
    wire N__42954;
    wire N__42951;
    wire N__42948;
    wire N__42943;
    wire N__42940;
    wire N__42939;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42929;
    wire N__42924;
    wire N__42921;
    wire N__42918;
    wire N__42913;
    wire N__42910;
    wire N__42909;
    wire N__42904;
    wire N__42903;
    wire N__42900;
    wire N__42897;
    wire N__42894;
    wire N__42889;
    wire N__42886;
    wire N__42885;
    wire N__42882;
    wire N__42879;
    wire N__42876;
    wire N__42875;
    wire N__42870;
    wire N__42867;
    wire N__42864;
    wire N__42859;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42848;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42832;
    wire N__42829;
    wire N__42828;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42816;
    wire N__42815;
    wire N__42810;
    wire N__42807;
    wire N__42804;
    wire N__42799;
    wire N__42796;
    wire N__42795;
    wire N__42792;
    wire N__42791;
    wire N__42788;
    wire N__42785;
    wire N__42782;
    wire N__42777;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42765;
    wire N__42764;
    wire N__42759;
    wire N__42756;
    wire N__42753;
    wire N__42748;
    wire N__42745;
    wire N__42742;
    wire N__42741;
    wire N__42738;
    wire N__42735;
    wire N__42730;
    wire N__42729;
    wire N__42726;
    wire N__42723;
    wire N__42720;
    wire N__42715;
    wire N__42712;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42700;
    wire N__42699;
    wire N__42696;
    wire N__42693;
    wire N__42690;
    wire N__42685;
    wire N__42682;
    wire N__42681;
    wire N__42676;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42661;
    wire N__42658;
    wire N__42657;
    wire N__42652;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42637;
    wire N__42634;
    wire N__42631;
    wire N__42630;
    wire N__42629;
    wire N__42628;
    wire N__42623;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42609;
    wire N__42606;
    wire N__42601;
    wire N__42600;
    wire N__42595;
    wire N__42592;
    wire N__42591;
    wire N__42590;
    wire N__42589;
    wire N__42588;
    wire N__42585;
    wire N__42580;
    wire N__42575;
    wire N__42568;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42554;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42538;
    wire N__42535;
    wire N__42532;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42519;
    wire N__42518;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42502;
    wire N__42499;
    wire N__42498;
    wire N__42497;
    wire N__42492;
    wire N__42489;
    wire N__42486;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42474;
    wire N__42469;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42454;
    wire N__42451;
    wire N__42450;
    wire N__42447;
    wire N__42444;
    wire N__42439;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42424;
    wire N__42421;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42409;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42394;
    wire N__42391;
    wire N__42390;
    wire N__42385;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42370;
    wire N__42367;
    wire N__42366;
    wire N__42361;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42351;
    wire N__42346;
    wire N__42343;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42333;
    wire N__42332;
    wire N__42331;
    wire N__42328;
    wire N__42325;
    wire N__42322;
    wire N__42319;
    wire N__42318;
    wire N__42317;
    wire N__42316;
    wire N__42315;
    wire N__42314;
    wire N__42313;
    wire N__42312;
    wire N__42311;
    wire N__42310;
    wire N__42309;
    wire N__42308;
    wire N__42307;
    wire N__42306;
    wire N__42305;
    wire N__42296;
    wire N__42287;
    wire N__42272;
    wire N__42271;
    wire N__42270;
    wire N__42267;
    wire N__42264;
    wire N__42261;
    wire N__42254;
    wire N__42251;
    wire N__42250;
    wire N__42247;
    wire N__42242;
    wire N__42237;
    wire N__42232;
    wire N__42231;
    wire N__42230;
    wire N__42227;
    wire N__42220;
    wire N__42219;
    wire N__42214;
    wire N__42211;
    wire N__42208;
    wire N__42205;
    wire N__42196;
    wire N__42195;
    wire N__42192;
    wire N__42191;
    wire N__42190;
    wire N__42189;
    wire N__42188;
    wire N__42187;
    wire N__42184;
    wire N__42179;
    wire N__42178;
    wire N__42177;
    wire N__42176;
    wire N__42175;
    wire N__42174;
    wire N__42173;
    wire N__42172;
    wire N__42169;
    wire N__42166;
    wire N__42163;
    wire N__42160;
    wire N__42157;
    wire N__42154;
    wire N__42153;
    wire N__42152;
    wire N__42151;
    wire N__42150;
    wire N__42147;
    wire N__42144;
    wire N__42141;
    wire N__42138;
    wire N__42137;
    wire N__42136;
    wire N__42135;
    wire N__42134;
    wire N__42133;
    wire N__42132;
    wire N__42117;
    wire N__42114;
    wire N__42111;
    wire N__42102;
    wire N__42085;
    wire N__42080;
    wire N__42077;
    wire N__42070;
    wire N__42061;
    wire N__42058;
    wire N__42057;
    wire N__42056;
    wire N__42055;
    wire N__42054;
    wire N__42053;
    wire N__42052;
    wire N__42051;
    wire N__42050;
    wire N__42049;
    wire N__42048;
    wire N__42047;
    wire N__42046;
    wire N__42045;
    wire N__42044;
    wire N__42043;
    wire N__42042;
    wire N__42039;
    wire N__42024;
    wire N__42007;
    wire N__42006;
    wire N__42005;
    wire N__42004;
    wire N__42003;
    wire N__42002;
    wire N__41999;
    wire N__41994;
    wire N__41991;
    wire N__41982;
    wire N__41979;
    wire N__41978;
    wire N__41975;
    wire N__41968;
    wire N__41967;
    wire N__41962;
    wire N__41959;
    wire N__41956;
    wire N__41953;
    wire N__41944;
    wire N__41941;
    wire N__41938;
    wire N__41935;
    wire N__41932;
    wire N__41931;
    wire N__41928;
    wire N__41927;
    wire N__41924;
    wire N__41921;
    wire N__41918;
    wire N__41913;
    wire N__41908;
    wire N__41905;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41895;
    wire N__41890;
    wire N__41887;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41873;
    wire N__41870;
    wire N__41867;
    wire N__41864;
    wire N__41857;
    wire N__41854;
    wire N__41851;
    wire N__41848;
    wire N__41847;
    wire N__41844;
    wire N__41841;
    wire N__41838;
    wire N__41835;
    wire N__41832;
    wire N__41829;
    wire N__41824;
    wire N__41821;
    wire N__41820;
    wire N__41819;
    wire N__41818;
    wire N__41817;
    wire N__41806;
    wire N__41803;
    wire N__41800;
    wire N__41797;
    wire N__41794;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41782;
    wire N__41779;
    wire N__41776;
    wire N__41773;
    wire N__41770;
    wire N__41767;
    wire N__41764;
    wire N__41761;
    wire N__41758;
    wire N__41755;
    wire N__41752;
    wire N__41751;
    wire N__41750;
    wire N__41747;
    wire N__41744;
    wire N__41741;
    wire N__41738;
    wire N__41731;
    wire N__41728;
    wire N__41727;
    wire N__41722;
    wire N__41721;
    wire N__41718;
    wire N__41715;
    wire N__41712;
    wire N__41709;
    wire N__41706;
    wire N__41705;
    wire N__41702;
    wire N__41699;
    wire N__41696;
    wire N__41689;
    wire N__41686;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41678;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41662;
    wire N__41661;
    wire N__41658;
    wire N__41655;
    wire N__41654;
    wire N__41651;
    wire N__41648;
    wire N__41645;
    wire N__41642;
    wire N__41639;
    wire N__41638;
    wire N__41635;
    wire N__41632;
    wire N__41629;
    wire N__41626;
    wire N__41617;
    wire N__41614;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41606;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41590;
    wire N__41587;
    wire N__41584;
    wire N__41581;
    wire N__41580;
    wire N__41579;
    wire N__41576;
    wire N__41571;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41561;
    wire N__41554;
    wire N__41551;
    wire N__41548;
    wire N__41547;
    wire N__41546;
    wire N__41543;
    wire N__41540;
    wire N__41537;
    wire N__41532;
    wire N__41527;
    wire N__41526;
    wire N__41521;
    wire N__41520;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41510;
    wire N__41507;
    wire N__41504;
    wire N__41501;
    wire N__41494;
    wire N__41491;
    wire N__41490;
    wire N__41485;
    wire N__41484;
    wire N__41481;
    wire N__41478;
    wire N__41475;
    wire N__41470;
    wire N__41469;
    wire N__41468;
    wire N__41465;
    wire N__41460;
    wire N__41457;
    wire N__41454;
    wire N__41451;
    wire N__41450;
    wire N__41447;
    wire N__41444;
    wire N__41441;
    wire N__41434;
    wire N__41431;
    wire N__41430;
    wire N__41427;
    wire N__41426;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41412;
    wire N__41407;
    wire N__41406;
    wire N__41405;
    wire N__41402;
    wire N__41397;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41384;
    wire N__41381;
    wire N__41378;
    wire N__41375;
    wire N__41368;
    wire N__41365;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41355;
    wire N__41354;
    wire N__41349;
    wire N__41346;
    wire N__41343;
    wire N__41338;
    wire N__41337;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41290;
    wire N__41287;
    wire N__41286;
    wire N__41283;
    wire N__41280;
    wire N__41277;
    wire N__41272;
    wire N__41271;
    wire N__41270;
    wire N__41267;
    wire N__41264;
    wire N__41261;
    wire N__41256;
    wire N__41251;
    wire N__41248;
    wire N__41247;
    wire N__41244;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41231;
    wire N__41228;
    wire N__41225;
    wire N__41222;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41208;
    wire N__41207;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41191;
    wire N__41190;
    wire N__41187;
    wire N__41184;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41143;
    wire N__41140;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41132;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41116;
    wire N__41115;
    wire N__41112;
    wire N__41111;
    wire N__41108;
    wire N__41105;
    wire N__41102;
    wire N__41099;
    wire N__41094;
    wire N__41091;
    wire N__41090;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41074;
    wire N__41071;
    wire N__41070;
    wire N__41067;
    wire N__41064;
    wire N__41063;
    wire N__41058;
    wire N__41055;
    wire N__41052;
    wire N__41047;
    wire N__41044;
    wire N__41043;
    wire N__41040;
    wire N__41037;
    wire N__41036;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41005;
    wire N__41002;
    wire N__41001;
    wire N__41000;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40984;
    wire N__40983;
    wire N__40982;
    wire N__40979;
    wire N__40974;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40949;
    wire N__40942;
    wire N__40939;
    wire N__40938;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40928;
    wire N__40923;
    wire N__40920;
    wire N__40917;
    wire N__40912;
    wire N__40911;
    wire N__40906;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40894;
    wire N__40891;
    wire N__40888;
    wire N__40887;
    wire N__40884;
    wire N__40881;
    wire N__40876;
    wire N__40873;
    wire N__40870;
    wire N__40867;
    wire N__40866;
    wire N__40863;
    wire N__40862;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40848;
    wire N__40843;
    wire N__40842;
    wire N__40839;
    wire N__40838;
    wire N__40835;
    wire N__40832;
    wire N__40829;
    wire N__40826;
    wire N__40821;
    wire N__40818;
    wire N__40815;
    wire N__40814;
    wire N__40811;
    wire N__40808;
    wire N__40805;
    wire N__40798;
    wire N__40795;
    wire N__40794;
    wire N__40793;
    wire N__40790;
    wire N__40787;
    wire N__40784;
    wire N__40781;
    wire N__40774;
    wire N__40771;
    wire N__40770;
    wire N__40765;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40752;
    wire N__40749;
    wire N__40748;
    wire N__40745;
    wire N__40742;
    wire N__40739;
    wire N__40732;
    wire N__40729;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40721;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40705;
    wire N__40702;
    wire N__40701;
    wire N__40698;
    wire N__40697;
    wire N__40694;
    wire N__40691;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40679;
    wire N__40676;
    wire N__40673;
    wire N__40670;
    wire N__40663;
    wire N__40660;
    wire N__40659;
    wire N__40656;
    wire N__40653;
    wire N__40652;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40636;
    wire N__40633;
    wire N__40632;
    wire N__40629;
    wire N__40628;
    wire N__40625;
    wire N__40622;
    wire N__40619;
    wire N__40616;
    wire N__40613;
    wire N__40610;
    wire N__40607;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40585;
    wire N__40582;
    wire N__40581;
    wire N__40580;
    wire N__40575;
    wire N__40572;
    wire N__40569;
    wire N__40564;
    wire N__40563;
    wire N__40562;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40541;
    wire N__40538;
    wire N__40535;
    wire N__40532;
    wire N__40525;
    wire N__40522;
    wire N__40521;
    wire N__40520;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40504;
    wire N__40503;
    wire N__40502;
    wire N__40499;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40478;
    wire N__40473;
    wire N__40472;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40456;
    wire N__40453;
    wire N__40450;
    wire N__40447;
    wire N__40446;
    wire N__40443;
    wire N__40442;
    wire N__40439;
    wire N__40436;
    wire N__40433;
    wire N__40428;
    wire N__40423;
    wire N__40420;
    wire N__40419;
    wire N__40416;
    wire N__40413;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40394;
    wire N__40393;
    wire N__40390;
    wire N__40387;
    wire N__40384;
    wire N__40381;
    wire N__40372;
    wire N__40369;
    wire N__40368;
    wire N__40365;
    wire N__40362;
    wire N__40359;
    wire N__40358;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40342;
    wire N__40341;
    wire N__40340;
    wire N__40337;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40319;
    wire N__40316;
    wire N__40313;
    wire N__40310;
    wire N__40303;
    wire N__40300;
    wire N__40299;
    wire N__40298;
    wire N__40295;
    wire N__40292;
    wire N__40289;
    wire N__40284;
    wire N__40279;
    wire N__40276;
    wire N__40273;
    wire N__40270;
    wire N__40269;
    wire N__40266;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40247;
    wire N__40244;
    wire N__40243;
    wire N__40240;
    wire N__40237;
    wire N__40234;
    wire N__40231;
    wire N__40222;
    wire N__40219;
    wire N__40218;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40198;
    wire N__40195;
    wire N__40194;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40154;
    wire N__40147;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40118;
    wire N__40115;
    wire N__40112;
    wire N__40109;
    wire N__40102;
    wire N__40101;
    wire N__40096;
    wire N__40095;
    wire N__40092;
    wire N__40089;
    wire N__40084;
    wire N__40083;
    wire N__40082;
    wire N__40079;
    wire N__40076;
    wire N__40073;
    wire N__40070;
    wire N__40065;
    wire N__40060;
    wire N__40059;
    wire N__40058;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40044;
    wire N__40041;
    wire N__40038;
    wire N__40037;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40021;
    wire N__40018;
    wire N__40017;
    wire N__40016;
    wire N__40013;
    wire N__40010;
    wire N__40007;
    wire N__40004;
    wire N__39997;
    wire N__39994;
    wire N__39991;
    wire N__39990;
    wire N__39989;
    wire N__39986;
    wire N__39983;
    wire N__39980;
    wire N__39975;
    wire N__39972;
    wire N__39971;
    wire N__39966;
    wire N__39963;
    wire N__39958;
    wire N__39955;
    wire N__39954;
    wire N__39953;
    wire N__39950;
    wire N__39947;
    wire N__39944;
    wire N__39941;
    wire N__39934;
    wire N__39931;
    wire N__39930;
    wire N__39929;
    wire N__39926;
    wire N__39921;
    wire N__39918;
    wire N__39917;
    wire N__39914;
    wire N__39911;
    wire N__39908;
    wire N__39901;
    wire N__39898;
    wire N__39895;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39879;
    wire N__39878;
    wire N__39877;
    wire N__39876;
    wire N__39875;
    wire N__39862;
    wire N__39859;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39831;
    wire N__39828;
    wire N__39825;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39815;
    wire N__39814;
    wire N__39811;
    wire N__39806;
    wire N__39803;
    wire N__39800;
    wire N__39797;
    wire N__39794;
    wire N__39787;
    wire N__39786;
    wire N__39783;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39764;
    wire N__39763;
    wire N__39760;
    wire N__39755;
    wire N__39752;
    wire N__39745;
    wire N__39742;
    wire N__39741;
    wire N__39740;
    wire N__39737;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39712;
    wire N__39709;
    wire N__39706;
    wire N__39701;
    wire N__39694;
    wire N__39691;
    wire N__39690;
    wire N__39687;
    wire N__39684;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39666;
    wire N__39663;
    wire N__39660;
    wire N__39655;
    wire N__39652;
    wire N__39643;
    wire N__39642;
    wire N__39639;
    wire N__39636;
    wire N__39635;
    wire N__39632;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39611;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39597;
    wire N__39594;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39584;
    wire N__39583;
    wire N__39580;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39567;
    wire N__39564;
    wire N__39553;
    wire N__39550;
    wire N__39549;
    wire N__39546;
    wire N__39545;
    wire N__39542;
    wire N__39539;
    wire N__39536;
    wire N__39533;
    wire N__39530;
    wire N__39525;
    wire N__39520;
    wire N__39517;
    wire N__39514;
    wire N__39511;
    wire N__39508;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39490;
    wire N__39487;
    wire N__39484;
    wire N__39481;
    wire N__39478;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39451;
    wire N__39448;
    wire N__39445;
    wire N__39442;
    wire N__39439;
    wire N__39436;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39424;
    wire N__39421;
    wire N__39418;
    wire N__39415;
    wire N__39412;
    wire N__39409;
    wire N__39406;
    wire N__39403;
    wire N__39400;
    wire N__39397;
    wire N__39394;
    wire N__39391;
    wire N__39388;
    wire N__39385;
    wire N__39382;
    wire N__39379;
    wire N__39376;
    wire N__39373;
    wire N__39370;
    wire N__39367;
    wire N__39364;
    wire N__39361;
    wire N__39358;
    wire N__39355;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39340;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39313;
    wire N__39310;
    wire N__39307;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39289;
    wire N__39286;
    wire N__39283;
    wire N__39280;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39268;
    wire N__39265;
    wire N__39262;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39244;
    wire N__39241;
    wire N__39238;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39226;
    wire N__39223;
    wire N__39220;
    wire N__39219;
    wire N__39216;
    wire N__39215;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39200;
    wire N__39197;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39181;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39165;
    wire N__39164;
    wire N__39161;
    wire N__39156;
    wire N__39151;
    wire N__39150;
    wire N__39147;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39135;
    wire N__39130;
    wire N__39129;
    wire N__39124;
    wire N__39123;
    wire N__39122;
    wire N__39119;
    wire N__39116;
    wire N__39113;
    wire N__39112;
    wire N__39107;
    wire N__39102;
    wire N__39099;
    wire N__39094;
    wire N__39091;
    wire N__39090;
    wire N__39089;
    wire N__39082;
    wire N__39081;
    wire N__39080;
    wire N__39079;
    wire N__39076;
    wire N__39069;
    wire N__39066;
    wire N__39063;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39045;
    wire N__39042;
    wire N__39039;
    wire N__39038;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39028;
    wire N__39025;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39011;
    wire N__39004;
    wire N__39003;
    wire N__39002;
    wire N__38999;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38969;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38955;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38913;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38903;
    wire N__38898;
    wire N__38897;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38885;
    wire N__38884;
    wire N__38883;
    wire N__38876;
    wire N__38873;
    wire N__38870;
    wire N__38869;
    wire N__38868;
    wire N__38867;
    wire N__38864;
    wire N__38861;
    wire N__38858;
    wire N__38851;
    wire N__38848;
    wire N__38845;
    wire N__38836;
    wire N__38833;
    wire N__38830;
    wire N__38827;
    wire N__38826;
    wire N__38825;
    wire N__38824;
    wire N__38823;
    wire N__38820;
    wire N__38815;
    wire N__38810;
    wire N__38805;
    wire N__38800;
    wire N__38799;
    wire N__38798;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38761;
    wire N__38758;
    wire N__38755;
    wire N__38752;
    wire N__38749;
    wire N__38746;
    wire N__38743;
    wire N__38740;
    wire N__38737;
    wire N__38734;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38701;
    wire N__38698;
    wire N__38695;
    wire N__38692;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38680;
    wire N__38677;
    wire N__38674;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38626;
    wire N__38623;
    wire N__38620;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38581;
    wire N__38578;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38560;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38523;
    wire N__38520;
    wire N__38517;
    wire N__38512;
    wire N__38509;
    wire N__38506;
    wire N__38503;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38491;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38458;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38446;
    wire N__38443;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38413;
    wire N__38410;
    wire N__38407;
    wire N__38406;
    wire N__38403;
    wire N__38402;
    wire N__38399;
    wire N__38396;
    wire N__38393;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38368;
    wire N__38365;
    wire N__38362;
    wire N__38359;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38299;
    wire N__38296;
    wire N__38293;
    wire N__38290;
    wire N__38287;
    wire N__38284;
    wire N__38281;
    wire N__38280;
    wire N__38277;
    wire N__38274;
    wire N__38269;
    wire N__38266;
    wire N__38263;
    wire N__38260;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38250;
    wire N__38247;
    wire N__38244;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38218;
    wire N__38217;
    wire N__38214;
    wire N__38211;
    wire N__38206;
    wire N__38203;
    wire N__38200;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38158;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38074;
    wire N__38071;
    wire N__38068;
    wire N__38065;
    wire N__38062;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38032;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38002;
    wire N__37999;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37987;
    wire N__37984;
    wire N__37981;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37936;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37909;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37879;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37831;
    wire N__37828;
    wire N__37825;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37765;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37744;
    wire N__37741;
    wire N__37738;
    wire N__37735;
    wire N__37732;
    wire N__37729;
    wire N__37726;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37702;
    wire N__37699;
    wire N__37696;
    wire N__37693;
    wire N__37690;
    wire N__37687;
    wire N__37684;
    wire N__37681;
    wire N__37678;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37666;
    wire N__37663;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37639;
    wire N__37636;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37624;
    wire N__37621;
    wire N__37618;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37597;
    wire N__37594;
    wire N__37591;
    wire N__37588;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37549;
    wire N__37546;
    wire N__37543;
    wire N__37540;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37522;
    wire N__37519;
    wire N__37516;
    wire N__37513;
    wire N__37510;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37449;
    wire N__37448;
    wire N__37445;
    wire N__37444;
    wire N__37443;
    wire N__37440;
    wire N__37437;
    wire N__37432;
    wire N__37431;
    wire N__37428;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37413;
    wire N__37410;
    wire N__37409;
    wire N__37408;
    wire N__37405;
    wire N__37402;
    wire N__37399;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37381;
    wire N__37376;
    wire N__37373;
    wire N__37368;
    wire N__37363;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37330;
    wire N__37329;
    wire N__37328;
    wire N__37323;
    wire N__37322;
    wire N__37321;
    wire N__37318;
    wire N__37317;
    wire N__37314;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37294;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37286;
    wire N__37285;
    wire N__37282;
    wire N__37277;
    wire N__37274;
    wire N__37267;
    wire N__37264;
    wire N__37261;
    wire N__37258;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37210;
    wire N__37207;
    wire N__37204;
    wire N__37201;
    wire N__37198;
    wire N__37195;
    wire N__37192;
    wire N__37189;
    wire N__37186;
    wire N__37183;
    wire N__37180;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37158;
    wire N__37153;
    wire N__37152;
    wire N__37149;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37134;
    wire N__37129;
    wire N__37128;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37113;
    wire N__37108;
    wire N__37107;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37092;
    wire N__37087;
    wire N__37084;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37066;
    wire N__37063;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37012;
    wire N__37011;
    wire N__37010;
    wire N__37009;
    wire N__37006;
    wire N__37005;
    wire N__37002;
    wire N__36993;
    wire N__36992;
    wire N__36991;
    wire N__36990;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36974;
    wire N__36973;
    wire N__36966;
    wire N__36963;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36949;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36828;
    wire N__36823;
    wire N__36822;
    wire N__36821;
    wire N__36818;
    wire N__36815;
    wire N__36812;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36793;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36757;
    wire N__36754;
    wire N__36751;
    wire N__36748;
    wire N__36745;
    wire N__36742;
    wire N__36739;
    wire N__36736;
    wire N__36733;
    wire N__36730;
    wire N__36727;
    wire N__36724;
    wire N__36721;
    wire N__36718;
    wire N__36715;
    wire N__36712;
    wire N__36709;
    wire N__36706;
    wire N__36703;
    wire N__36700;
    wire N__36697;
    wire N__36694;
    wire N__36691;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36676;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36666;
    wire N__36665;
    wire N__36664;
    wire N__36663;
    wire N__36662;
    wire N__36661;
    wire N__36660;
    wire N__36659;
    wire N__36658;
    wire N__36657;
    wire N__36656;
    wire N__36655;
    wire N__36654;
    wire N__36653;
    wire N__36652;
    wire N__36651;
    wire N__36650;
    wire N__36649;
    wire N__36648;
    wire N__36647;
    wire N__36646;
    wire N__36643;
    wire N__36630;
    wire N__36615;
    wire N__36614;
    wire N__36613;
    wire N__36612;
    wire N__36611;
    wire N__36596;
    wire N__36593;
    wire N__36588;
    wire N__36587;
    wire N__36586;
    wire N__36585;
    wire N__36584;
    wire N__36581;
    wire N__36572;
    wire N__36567;
    wire N__36566;
    wire N__36565;
    wire N__36564;
    wire N__36563;
    wire N__36562;
    wire N__36561;
    wire N__36558;
    wire N__36549;
    wire N__36544;
    wire N__36541;
    wire N__36534;
    wire N__36527;
    wire N__36526;
    wire N__36525;
    wire N__36520;
    wire N__36517;
    wire N__36510;
    wire N__36505;
    wire N__36496;
    wire N__36495;
    wire N__36492;
    wire N__36491;
    wire N__36490;
    wire N__36487;
    wire N__36484;
    wire N__36481;
    wire N__36478;
    wire N__36477;
    wire N__36474;
    wire N__36471;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36451;
    wire N__36450;
    wire N__36449;
    wire N__36446;
    wire N__36445;
    wire N__36444;
    wire N__36443;
    wire N__36442;
    wire N__36441;
    wire N__36440;
    wire N__36439;
    wire N__36438;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36422;
    wire N__36421;
    wire N__36420;
    wire N__36419;
    wire N__36418;
    wire N__36417;
    wire N__36414;
    wire N__36399;
    wire N__36398;
    wire N__36397;
    wire N__36396;
    wire N__36393;
    wire N__36386;
    wire N__36379;
    wire N__36376;
    wire N__36369;
    wire N__36368;
    wire N__36367;
    wire N__36362;
    wire N__36361;
    wire N__36360;
    wire N__36359;
    wire N__36358;
    wire N__36357;
    wire N__36354;
    wire N__36349;
    wire N__36348;
    wire N__36345;
    wire N__36344;
    wire N__36341;
    wire N__36340;
    wire N__36339;
    wire N__36336;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36325;
    wire N__36322;
    wire N__36321;
    wire N__36320;
    wire N__36319;
    wire N__36318;
    wire N__36317;
    wire N__36316;
    wire N__36315;
    wire N__36314;
    wire N__36311;
    wire N__36306;
    wire N__36295;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36271;
    wire N__36268;
    wire N__36255;
    wire N__36250;
    wire N__36235;
    wire N__36232;
    wire N__36231;
    wire N__36228;
    wire N__36227;
    wire N__36226;
    wire N__36223;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36213;
    wire N__36210;
    wire N__36207;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36185;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36166;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36150;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36129;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36114;
    wire N__36111;
    wire N__36108;
    wire N__36101;
    wire N__36094;
    wire N__36091;
    wire N__36088;
    wire N__36087;
    wire N__36086;
    wire N__36085;
    wire N__36082;
    wire N__36079;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36064;
    wire N__36063;
    wire N__36060;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36040;
    wire N__36031;
    wire N__36028;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36020;
    wire N__36019;
    wire N__36018;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36003;
    wire N__35996;
    wire N__35993;
    wire N__35986;
    wire N__35985;
    wire N__35984;
    wire N__35983;
    wire N__35980;
    wire N__35977;
    wire N__35974;
    wire N__35971;
    wire N__35968;
    wire N__35967;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35932;
    wire N__35931;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35910;
    wire N__35905;
    wire N__35900;
    wire N__35897;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35868;
    wire N__35863;
    wire N__35858;
    wire N__35855;
    wire N__35848;
    wire N__35845;
    wire N__35842;
    wire N__35841;
    wire N__35838;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35827;
    wire N__35824;
    wire N__35819;
    wire N__35816;
    wire N__35813;
    wire N__35810;
    wire N__35803;
    wire N__35802;
    wire N__35801;
    wire N__35798;
    wire N__35795;
    wire N__35792;
    wire N__35791;
    wire N__35790;
    wire N__35781;
    wire N__35780;
    wire N__35779;
    wire N__35778;
    wire N__35777;
    wire N__35776;
    wire N__35775;
    wire N__35774;
    wire N__35773;
    wire N__35770;
    wire N__35769;
    wire N__35766;
    wire N__35759;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35737;
    wire N__35734;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35713;
    wire N__35710;
    wire N__35709;
    wire N__35708;
    wire N__35705;
    wire N__35704;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35691;
    wire N__35688;
    wire N__35685;
    wire N__35680;
    wire N__35677;
    wire N__35668;
    wire N__35665;
    wire N__35664;
    wire N__35663;
    wire N__35662;
    wire N__35659;
    wire N__35658;
    wire N__35655;
    wire N__35652;
    wire N__35649;
    wire N__35646;
    wire N__35643;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35628;
    wire N__35625;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35607;
    wire N__35606;
    wire N__35605;
    wire N__35604;
    wire N__35603;
    wire N__35602;
    wire N__35601;
    wire N__35600;
    wire N__35599;
    wire N__35598;
    wire N__35597;
    wire N__35596;
    wire N__35595;
    wire N__35594;
    wire N__35593;
    wire N__35592;
    wire N__35591;
    wire N__35590;
    wire N__35589;
    wire N__35588;
    wire N__35587;
    wire N__35586;
    wire N__35585;
    wire N__35584;
    wire N__35583;
    wire N__35582;
    wire N__35581;
    wire N__35580;
    wire N__35579;
    wire N__35570;
    wire N__35561;
    wire N__35556;
    wire N__35547;
    wire N__35538;
    wire N__35529;
    wire N__35520;
    wire N__35511;
    wire N__35506;
    wire N__35497;
    wire N__35488;
    wire N__35485;
    wire N__35482;
    wire N__35481;
    wire N__35480;
    wire N__35477;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35459;
    wire N__35454;
    wire N__35451;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35425;
    wire N__35424;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35403;
    wire N__35400;
    wire N__35397;
    wire N__35392;
    wire N__35389;
    wire N__35380;
    wire N__35379;
    wire N__35378;
    wire N__35375;
    wire N__35374;
    wire N__35371;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35361;
    wire N__35358;
    wire N__35355;
    wire N__35352;
    wire N__35349;
    wire N__35346;
    wire N__35341;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35323;
    wire N__35320;
    wire N__35319;
    wire N__35316;
    wire N__35315;
    wire N__35314;
    wire N__35313;
    wire N__35310;
    wire N__35307;
    wire N__35304;
    wire N__35301;
    wire N__35298;
    wire N__35295;
    wire N__35290;
    wire N__35287;
    wire N__35284;
    wire N__35281;
    wire N__35278;
    wire N__35275;
    wire N__35266;
    wire N__35265;
    wire N__35262;
    wire N__35259;
    wire N__35256;
    wire N__35255;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35232;
    wire N__35229;
    wire N__35226;
    wire N__35219;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35130;
    wire N__35127;
    wire N__35122;
    wire N__35119;
    wire N__35118;
    wire N__35117;
    wire N__35114;
    wire N__35111;
    wire N__35108;
    wire N__35105;
    wire N__35102;
    wire N__35095;
    wire N__35092;
    wire N__35091;
    wire N__35090;
    wire N__35087;
    wire N__35084;
    wire N__35081;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35056;
    wire N__35055;
    wire N__35054;
    wire N__35051;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35039;
    wire N__35036;
    wire N__35029;
    wire N__35028;
    wire N__35025;
    wire N__35024;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35012;
    wire N__35009;
    wire N__35002;
    wire N__35001;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34986;
    wire N__34985;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34960;
    wire N__34959;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34932;
    wire N__34927;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34913;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34897;
    wire N__34894;
    wire N__34893;
    wire N__34890;
    wire N__34887;
    wire N__34884;
    wire N__34881;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34866;
    wire N__34865;
    wire N__34862;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34843;
    wire N__34834;
    wire N__34833;
    wire N__34830;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34819;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34794;
    wire N__34791;
    wire N__34788;
    wire N__34785;
    wire N__34784;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34759;
    wire N__34756;
    wire N__34755;
    wire N__34750;
    wire N__34749;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34723;
    wire N__34722;
    wire N__34719;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34708;
    wire N__34705;
    wire N__34702;
    wire N__34697;
    wire N__34694;
    wire N__34687;
    wire N__34686;
    wire N__34685;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34660;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34635;
    wire N__34632;
    wire N__34629;
    wire N__34628;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34616;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34600;
    wire N__34597;
    wire N__34596;
    wire N__34595;
    wire N__34594;
    wire N__34591;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34577;
    wire N__34574;
    wire N__34571;
    wire N__34568;
    wire N__34565;
    wire N__34558;
    wire N__34555;
    wire N__34554;
    wire N__34551;
    wire N__34550;
    wire N__34549;
    wire N__34546;
    wire N__34543;
    wire N__34540;
    wire N__34537;
    wire N__34534;
    wire N__34529;
    wire N__34522;
    wire N__34521;
    wire N__34516;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34505;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34479;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34469;
    wire N__34468;
    wire N__34463;
    wire N__34460;
    wire N__34457;
    wire N__34454;
    wire N__34451;
    wire N__34444;
    wire N__34441;
    wire N__34440;
    wire N__34439;
    wire N__34434;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34421;
    wire N__34418;
    wire N__34415;
    wire N__34412;
    wire N__34405;
    wire N__34402;
    wire N__34401;
    wire N__34400;
    wire N__34397;
    wire N__34394;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34373;
    wire N__34370;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34356;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34319;
    wire N__34312;
    wire N__34311;
    wire N__34308;
    wire N__34307;
    wire N__34304;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34276;
    wire N__34275;
    wire N__34272;
    wire N__34269;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34258;
    wire N__34253;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34241;
    wire N__34234;
    wire N__34233;
    wire N__34232;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34219;
    wire N__34216;
    wire N__34211;
    wire N__34208;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34161;
    wire N__34158;
    wire N__34155;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34122;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34107;
    wire N__34104;
    wire N__34101;
    wire N__34096;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34084;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34065;
    wire N__34062;
    wire N__34059;
    wire N__34058;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34033;
    wire N__34032;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34009;
    wire N__34006;
    wire N__34003;
    wire N__34002;
    wire N__34001;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33989;
    wire N__33986;
    wire N__33983;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33964;
    wire N__33961;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33943;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33916;
    wire N__33915;
    wire N__33914;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33898;
    wire N__33897;
    wire N__33894;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33862;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33780;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33766;
    wire N__33761;
    wire N__33758;
    wire N__33755;
    wire N__33752;
    wire N__33749;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33733;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33688;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33651;
    wire N__33650;
    wire N__33649;
    wire N__33648;
    wire N__33647;
    wire N__33646;
    wire N__33645;
    wire N__33640;
    wire N__33635;
    wire N__33634;
    wire N__33633;
    wire N__33632;
    wire N__33629;
    wire N__33628;
    wire N__33627;
    wire N__33626;
    wire N__33623;
    wire N__33622;
    wire N__33621;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33613;
    wire N__33608;
    wire N__33605;
    wire N__33604;
    wire N__33603;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33586;
    wire N__33575;
    wire N__33574;
    wire N__33567;
    wire N__33562;
    wire N__33561;
    wire N__33560;
    wire N__33559;
    wire N__33558;
    wire N__33557;
    wire N__33556;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33546;
    wire N__33545;
    wire N__33544;
    wire N__33541;
    wire N__33534;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33510;
    wire N__33501;
    wire N__33490;
    wire N__33485;
    wire N__33480;
    wire N__33473;
    wire N__33460;
    wire N__33457;
    wire N__33456;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33445;
    wire N__33444;
    wire N__33443;
    wire N__33442;
    wire N__33441;
    wire N__33438;
    wire N__33433;
    wire N__33424;
    wire N__33421;
    wire N__33412;
    wire N__33411;
    wire N__33408;
    wire N__33407;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33393;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33379;
    wire N__33370;
    wire N__33369;
    wire N__33366;
    wire N__33365;
    wire N__33364;
    wire N__33361;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33351;
    wire N__33348;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33327;
    wire N__33324;
    wire N__33319;
    wire N__33310;
    wire N__33309;
    wire N__33308;
    wire N__33307;
    wire N__33306;
    wire N__33303;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33266;
    wire N__33259;
    wire N__33258;
    wire N__33255;
    wire N__33254;
    wire N__33253;
    wire N__33250;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33226;
    wire N__33223;
    wire N__33216;
    wire N__33211;
    wire N__33210;
    wire N__33209;
    wire N__33208;
    wire N__33205;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33178;
    wire N__33175;
    wire N__33170;
    wire N__33163;
    wire N__33160;
    wire N__33159;
    wire N__33156;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33135;
    wire N__33130;
    wire N__33129;
    wire N__33126;
    wire N__33125;
    wire N__33122;
    wire N__33119;
    wire N__33116;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33066;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32947;
    wire N__32944;
    wire N__32941;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32926;
    wire N__32925;
    wire N__32924;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32913;
    wire N__32910;
    wire N__32909;
    wire N__32908;
    wire N__32907;
    wire N__32906;
    wire N__32905;
    wire N__32904;
    wire N__32903;
    wire N__32902;
    wire N__32901;
    wire N__32900;
    wire N__32899;
    wire N__32898;
    wire N__32897;
    wire N__32896;
    wire N__32895;
    wire N__32894;
    wire N__32889;
    wire N__32886;
    wire N__32869;
    wire N__32858;
    wire N__32853;
    wire N__32852;
    wire N__32851;
    wire N__32848;
    wire N__32843;
    wire N__32834;
    wire N__32831;
    wire N__32828;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32814;
    wire N__32811;
    wire N__32810;
    wire N__32805;
    wire N__32800;
    wire N__32797;
    wire N__32794;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32778;
    wire N__32777;
    wire N__32776;
    wire N__32775;
    wire N__32774;
    wire N__32773;
    wire N__32772;
    wire N__32771;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32760;
    wire N__32759;
    wire N__32758;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32737;
    wire N__32734;
    wire N__32733;
    wire N__32732;
    wire N__32731;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32703;
    wire N__32694;
    wire N__32691;
    wire N__32690;
    wire N__32687;
    wire N__32686;
    wire N__32685;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32669;
    wire N__32666;
    wire N__32661;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32630;
    wire N__32627;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32617;
    wire N__32610;
    wire N__32607;
    wire N__32596;
    wire N__32595;
    wire N__32594;
    wire N__32591;
    wire N__32590;
    wire N__32587;
    wire N__32586;
    wire N__32585;
    wire N__32584;
    wire N__32583;
    wire N__32582;
    wire N__32581;
    wire N__32580;
    wire N__32577;
    wire N__32576;
    wire N__32575;
    wire N__32574;
    wire N__32573;
    wire N__32572;
    wire N__32571;
    wire N__32570;
    wire N__32569;
    wire N__32568;
    wire N__32565;
    wire N__32548;
    wire N__32545;
    wire N__32530;
    wire N__32527;
    wire N__32526;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32510;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32499;
    wire N__32492;
    wire N__32489;
    wire N__32484;
    wire N__32481;
    wire N__32478;
    wire N__32473;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32461;
    wire N__32458;
    wire N__32453;
    wire N__32450;
    wire N__32443;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32428;
    wire N__32425;
    wire N__32422;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32407;
    wire N__32406;
    wire N__32403;
    wire N__32402;
    wire N__32401;
    wire N__32398;
    wire N__32395;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32368;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32351;
    wire N__32350;
    wire N__32349;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32331;
    wire N__32320;
    wire N__32317;
    wire N__32316;
    wire N__32315;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32293;
    wire N__32290;
    wire N__32287;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32251;
    wire N__32248;
    wire N__32245;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32188;
    wire N__32185;
    wire N__32182;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32149;
    wire N__32146;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32125;
    wire N__32122;
    wire N__32119;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32107;
    wire N__32104;
    wire N__32101;
    wire N__32098;
    wire N__32095;
    wire N__32092;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32080;
    wire N__32077;
    wire N__32074;
    wire N__32071;
    wire N__32068;
    wire N__32065;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32044;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32011;
    wire N__32008;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31990;
    wire N__31987;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31972;
    wire N__31969;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31948;
    wire N__31945;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31927;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31861;
    wire N__31858;
    wire N__31855;
    wire N__31852;
    wire N__31849;
    wire N__31846;
    wire N__31845;
    wire N__31844;
    wire N__31841;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31831;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31795;
    wire N__31792;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31784;
    wire N__31781;
    wire N__31778;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31762;
    wire N__31761;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31750;
    wire N__31747;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31699;
    wire N__31696;
    wire N__31693;
    wire N__31690;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31678;
    wire N__31675;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31561;
    wire N__31558;
    wire N__31555;
    wire N__31552;
    wire N__31549;
    wire N__31546;
    wire N__31543;
    wire N__31540;
    wire N__31537;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31501;
    wire N__31498;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31445;
    wire N__31444;
    wire N__31441;
    wire N__31436;
    wire N__31433;
    wire N__31432;
    wire N__31431;
    wire N__31424;
    wire N__31421;
    wire N__31418;
    wire N__31413;
    wire N__31412;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31395;
    wire N__31392;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31357;
    wire N__31356;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31341;
    wire N__31336;
    wire N__31333;
    wire N__31332;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31312;
    wire N__31309;
    wire N__31308;
    wire N__31307;
    wire N__31304;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31288;
    wire N__31285;
    wire N__31284;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31274;
    wire N__31269;
    wire N__31264;
    wire N__31261;
    wire N__31260;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31245;
    wire N__31240;
    wire N__31237;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31225;
    wire N__31222;
    wire N__31221;
    wire N__31220;
    wire N__31219;
    wire N__31218;
    wire N__31217;
    wire N__31216;
    wire N__31215;
    wire N__31214;
    wire N__31213;
    wire N__31212;
    wire N__31211;
    wire N__31210;
    wire N__31209;
    wire N__31208;
    wire N__31207;
    wire N__31206;
    wire N__31205;
    wire N__31204;
    wire N__31203;
    wire N__31202;
    wire N__31201;
    wire N__31200;
    wire N__31199;
    wire N__31198;
    wire N__31197;
    wire N__31196;
    wire N__31195;
    wire N__31194;
    wire N__31193;
    wire N__31188;
    wire N__31179;
    wire N__31170;
    wire N__31161;
    wire N__31152;
    wire N__31143;
    wire N__31134;
    wire N__31125;
    wire N__31116;
    wire N__31109;
    wire N__31104;
    wire N__31099;
    wire N__31096;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31084;
    wire N__31083;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31060;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31033;
    wire N__31032;
    wire N__31029;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31012;
    wire N__31009;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30992;
    wire N__30989;
    wire N__30988;
    wire N__30985;
    wire N__30984;
    wire N__30977;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30922;
    wire N__30917;
    wire N__30914;
    wire N__30907;
    wire N__30906;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30891;
    wire N__30886;
    wire N__30883;
    wire N__30882;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30862;
    wire N__30859;
    wire N__30858;
    wire N__30857;
    wire N__30854;
    wire N__30851;
    wire N__30848;
    wire N__30845;
    wire N__30838;
    wire N__30835;
    wire N__30834;
    wire N__30833;
    wire N__30830;
    wire N__30827;
    wire N__30824;
    wire N__30819;
    wire N__30814;
    wire N__30811;
    wire N__30810;
    wire N__30809;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30795;
    wire N__30790;
    wire N__30787;
    wire N__30786;
    wire N__30785;
    wire N__30782;
    wire N__30777;
    wire N__30772;
    wire N__30769;
    wire N__30768;
    wire N__30767;
    wire N__30764;
    wire N__30759;
    wire N__30754;
    wire N__30751;
    wire N__30750;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30735;
    wire N__30730;
    wire N__30727;
    wire N__30726;
    wire N__30725;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30711;
    wire N__30706;
    wire N__30703;
    wire N__30702;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30687;
    wire N__30682;
    wire N__30679;
    wire N__30678;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30658;
    wire N__30655;
    wire N__30654;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30641;
    wire N__30634;
    wire N__30631;
    wire N__30630;
    wire N__30629;
    wire N__30626;
    wire N__30623;
    wire N__30620;
    wire N__30615;
    wire N__30610;
    wire N__30607;
    wire N__30606;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30591;
    wire N__30586;
    wire N__30583;
    wire N__30582;
    wire N__30581;
    wire N__30578;
    wire N__30573;
    wire N__30568;
    wire N__30565;
    wire N__30564;
    wire N__30563;
    wire N__30560;
    wire N__30555;
    wire N__30550;
    wire N__30547;
    wire N__30546;
    wire N__30545;
    wire N__30542;
    wire N__30539;
    wire N__30536;
    wire N__30531;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30519;
    wire N__30516;
    wire N__30515;
    wire N__30512;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30490;
    wire N__30487;
    wire N__30486;
    wire N__30485;
    wire N__30484;
    wire N__30483;
    wire N__30482;
    wire N__30481;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30469;
    wire N__30468;
    wire N__30467;
    wire N__30460;
    wire N__30457;
    wire N__30456;
    wire N__30455;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30441;
    wire N__30438;
    wire N__30437;
    wire N__30434;
    wire N__30429;
    wire N__30428;
    wire N__30427;
    wire N__30426;
    wire N__30425;
    wire N__30424;
    wire N__30423;
    wire N__30422;
    wire N__30421;
    wire N__30420;
    wire N__30419;
    wire N__30418;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30402;
    wire N__30397;
    wire N__30382;
    wire N__30373;
    wire N__30358;
    wire N__30357;
    wire N__30356;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30337;
    wire N__30336;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30319;
    wire N__30316;
    wire N__30315;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30298;
    wire N__30295;
    wire N__30294;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30279;
    wire N__30274;
    wire N__30271;
    wire N__30270;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30255;
    wire N__30250;
    wire N__30247;
    wire N__30246;
    wire N__30245;
    wire N__30242;
    wire N__30237;
    wire N__30232;
    wire N__30229;
    wire N__30228;
    wire N__30227;
    wire N__30224;
    wire N__30219;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30174;
    wire N__30173;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30145;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30043;
    wire N__30040;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30019;
    wire N__30016;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29991;
    wire N__29990;
    wire N__29987;
    wire N__29982;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29970;
    wire N__29969;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29956;
    wire N__29947;
    wire N__29946;
    wire N__29943;
    wire N__29940;
    wire N__29937;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29927;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29905;
    wire N__29904;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29886;
    wire N__29881;
    wire N__29880;
    wire N__29879;
    wire N__29878;
    wire N__29877;
    wire N__29874;
    wire N__29871;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29857;
    wire N__29854;
    wire N__29851;
    wire N__29848;
    wire N__29845;
    wire N__29840;
    wire N__29833;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29822;
    wire N__29819;
    wire N__29816;
    wire N__29815;
    wire N__29812;
    wire N__29807;
    wire N__29804;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29788;
    wire N__29785;
    wire N__29782;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29721;
    wire N__29720;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29695;
    wire N__29694;
    wire N__29693;
    wire N__29692;
    wire N__29691;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29664;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29637;
    wire N__29636;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29620;
    wire N__29617;
    wire N__29616;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29590;
    wire N__29587;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29572;
    wire N__29569;
    wire N__29568;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29553;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29529;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29512;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29500;
    wire N__29497;
    wire N__29496;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29476;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29457;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29442;
    wire N__29439;
    wire N__29438;
    wire N__29435;
    wire N__29432;
    wire N__29429;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29405;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29379;
    wire N__29376;
    wire N__29373;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29356;
    wire N__29353;
    wire N__29352;
    wire N__29349;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29333;
    wire N__29330;
    wire N__29327;
    wire N__29324;
    wire N__29319;
    wire N__29314;
    wire N__29311;
    wire N__29308;
    wire N__29307;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29271;
    wire N__29270;
    wire N__29269;
    wire N__29268;
    wire N__29267;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29255;
    wire N__29252;
    wire N__29247;
    wire N__29240;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29215;
    wire N__29212;
    wire N__29209;
    wire N__29208;
    wire N__29205;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29187;
    wire N__29182;
    wire N__29179;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29162;
    wire N__29159;
    wire N__29152;
    wire N__29149;
    wire N__29148;
    wire N__29145;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29130;
    wire N__29125;
    wire N__29122;
    wire N__29121;
    wire N__29118;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29106;
    wire N__29101;
    wire N__29100;
    wire N__29097;
    wire N__29094;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29073;
    wire N__29070;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28986;
    wire N__28983;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28965;
    wire N__28964;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28950;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28889;
    wire N__28882;
    wire N__28879;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28866;
    wire N__28863;
    wire N__28860;
    wire N__28857;
    wire N__28854;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28804;
    wire N__28801;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28723;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28674;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28647;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28453;
    wire N__28450;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28281;
    wire N__28278;
    wire N__28275;
    wire N__28272;
    wire N__28267;
    wire N__28264;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28147;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27964;
    wire N__27963;
    wire N__27960;
    wire N__27957;
    wire N__27954;
    wire N__27951;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27936;
    wire N__27931;
    wire N__27930;
    wire N__27929;
    wire N__27928;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27916;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27868;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27846;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27792;
    wire N__27791;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27775;
    wire N__27774;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27757;
    wire N__27756;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27739;
    wire N__27738;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27721;
    wire N__27720;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27703;
    wire N__27700;
    wire N__27699;
    wire N__27698;
    wire N__27697;
    wire N__27696;
    wire N__27695;
    wire N__27694;
    wire N__27693;
    wire N__27692;
    wire N__27691;
    wire N__27682;
    wire N__27677;
    wire N__27668;
    wire N__27661;
    wire N__27660;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27650;
    wire N__27643;
    wire N__27642;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27625;
    wire N__27624;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27607;
    wire N__27606;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27589;
    wire N__27586;
    wire N__27585;
    wire N__27584;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27532;
    wire N__27529;
    wire N__27528;
    wire N__27527;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27478;
    wire N__27475;
    wire N__27472;
    wire N__27469;
    wire N__27468;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27453;
    wire N__27452;
    wire N__27449;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27433;
    wire N__27430;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27378;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27345;
    wire N__27344;
    wire N__27343;
    wire N__27342;
    wire N__27341;
    wire N__27338;
    wire N__27337;
    wire N__27334;
    wire N__27333;
    wire N__27330;
    wire N__27327;
    wire N__27312;
    wire N__27309;
    wire N__27306;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27280;
    wire N__27277;
    wire N__27274;
    wire N__27273;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27232;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27115;
    wire N__27112;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27079;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27040;
    wire N__27037;
    wire N__27034;
    wire N__27031;
    wire N__27028;
    wire N__27025;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26881;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26869;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26820;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26810;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26800;
    wire N__26797;
    wire N__26792;
    wire N__26785;
    wire N__26784;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26742;
    wire N__26739;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26704;
    wire N__26701;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26691;
    wire N__26688;
    wire N__26687;
    wire N__26684;
    wire N__26681;
    wire N__26678;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26646;
    wire N__26643;
    wire N__26642;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26617;
    wire N__26614;
    wire N__26613;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26575;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26567;
    wire N__26564;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26527;
    wire N__26526;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26498;
    wire N__26491;
    wire N__26490;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26455;
    wire N__26454;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26444;
    wire N__26441;
    wire N__26440;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26407;
    wire N__26406;
    wire N__26403;
    wire N__26402;
    wire N__26401;
    wire N__26398;
    wire N__26395;
    wire N__26392;
    wire N__26389;
    wire N__26386;
    wire N__26377;
    wire N__26376;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26353;
    wire N__26350;
    wire N__26347;
    wire N__26338;
    wire N__26337;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26302;
    wire N__26301;
    wire N__26298;
    wire N__26295;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26257;
    wire N__26256;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26206;
    wire N__26205;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26190;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26180;
    wire N__26177;
    wire N__26176;
    wire N__26173;
    wire N__26170;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26153;
    wire N__26146;
    wire N__26143;
    wire N__26140;
    wire N__26139;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26121;
    wire N__26118;
    wire N__26115;
    wire N__26110;
    wire N__26107;
    wire N__26104;
    wire N__26101;
    wire N__26098;
    wire N__26095;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26083;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26067;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26050;
    wire N__26047;
    wire N__26044;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26007;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25990;
    wire N__25989;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25972;
    wire N__25971;
    wire N__25970;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25952;
    wire N__25945;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25933;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25918;
    wire N__25917;
    wire N__25914;
    wire N__25911;
    wire N__25906;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25894;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25882;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25870;
    wire N__25869;
    wire N__25866;
    wire N__25863;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25848;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25805;
    wire N__25802;
    wire N__25801;
    wire N__25796;
    wire N__25795;
    wire N__25794;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25779;
    wire N__25776;
    wire N__25765;
    wire N__25762;
    wire N__25761;
    wire N__25758;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25707;
    wire N__25706;
    wire N__25705;
    wire N__25704;
    wire N__25703;
    wire N__25700;
    wire N__25699;
    wire N__25698;
    wire N__25697;
    wire N__25696;
    wire N__25685;
    wire N__25678;
    wire N__25677;
    wire N__25676;
    wire N__25673;
    wire N__25672;
    wire N__25671;
    wire N__25670;
    wire N__25667;
    wire N__25662;
    wire N__25659;
    wire N__25658;
    wire N__25657;
    wire N__25656;
    wire N__25655;
    wire N__25654;
    wire N__25653;
    wire N__25652;
    wire N__25651;
    wire N__25650;
    wire N__25649;
    wire N__25646;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25623;
    wire N__25622;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25614;
    wire N__25607;
    wire N__25600;
    wire N__25595;
    wire N__25586;
    wire N__25575;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25555;
    wire N__25554;
    wire N__25553;
    wire N__25552;
    wire N__25551;
    wire N__25550;
    wire N__25549;
    wire N__25548;
    wire N__25547;
    wire N__25546;
    wire N__25545;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25528;
    wire N__25527;
    wire N__25526;
    wire N__25523;
    wire N__25522;
    wire N__25521;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25510;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25482;
    wire N__25479;
    wire N__25478;
    wire N__25477;
    wire N__25476;
    wire N__25475;
    wire N__25474;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25449;
    wire N__25440;
    wire N__25433;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25421;
    wire N__25418;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25410;
    wire N__25407;
    wire N__25402;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25386;
    wire N__25379;
    wire N__25374;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25351;
    wire N__25336;
    wire N__25335;
    wire N__25334;
    wire N__25333;
    wire N__25332;
    wire N__25331;
    wire N__25330;
    wire N__25329;
    wire N__25328;
    wire N__25327;
    wire N__25326;
    wire N__25325;
    wire N__25324;
    wire N__25323;
    wire N__25322;
    wire N__25321;
    wire N__25318;
    wire N__25307;
    wire N__25300;
    wire N__25295;
    wire N__25294;
    wire N__25293;
    wire N__25292;
    wire N__25291;
    wire N__25290;
    wire N__25289;
    wire N__25286;
    wire N__25277;
    wire N__25274;
    wire N__25267;
    wire N__25264;
    wire N__25253;
    wire N__25252;
    wire N__25251;
    wire N__25250;
    wire N__25249;
    wire N__25248;
    wire N__25247;
    wire N__25242;
    wire N__25235;
    wire N__25232;
    wire N__25219;
    wire N__25210;
    wire N__25209;
    wire N__25208;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25197;
    wire N__25196;
    wire N__25195;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25183;
    wire N__25180;
    wire N__25179;
    wire N__25178;
    wire N__25175;
    wire N__25174;
    wire N__25173;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25156;
    wire N__25155;
    wire N__25154;
    wire N__25153;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25135;
    wire N__25134;
    wire N__25133;
    wire N__25132;
    wire N__25129;
    wire N__25124;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25106;
    wire N__25101;
    wire N__25098;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25081;
    wire N__25078;
    wire N__25077;
    wire N__25074;
    wire N__25065;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25054;
    wire N__25049;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25025;
    wire N__25022;
    wire N__25015;
    wire N__25012;
    wire N__25007;
    wire N__25002;
    wire N__24997;
    wire N__24994;
    wire N__24987;
    wire N__24980;
    wire N__24973;
    wire N__24972;
    wire N__24969;
    wire N__24968;
    wire N__24965;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24923;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24901;
    wire N__24900;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24883;
    wire N__24880;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24859;
    wire N__24858;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24825;
    wire N__24822;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24811;
    wire N__24808;
    wire N__24803;
    wire N__24800;
    wire N__24795;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24673;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24626;
    wire N__24623;
    wire N__24622;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24595;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24587;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24555;
    wire N__24554;
    wire N__24553;
    wire N__24550;
    wire N__24543;
    wire N__24542;
    wire N__24541;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24525;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24451;
    wire N__24448;
    wire N__24445;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24369;
    wire N__24366;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24349;
    wire N__24348;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24331;
    wire N__24330;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24307;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24270;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24255;
    wire N__24250;
    wire N__24245;
    wire N__24242;
    wire N__24235;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24183;
    wire N__24180;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24169;
    wire N__24168;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24109;
    wire N__24106;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24094;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24078;
    wire N__24077;
    wire N__24074;
    wire N__24073;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24054;
    wire N__24051;
    wire N__24046;
    wire N__24043;
    wire N__24040;
    wire N__24037;
    wire N__24034;
    wire N__24033;
    wire N__24032;
    wire N__24029;
    wire N__24024;
    wire N__24021;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23980;
    wire N__23977;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23947;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23930;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23914;
    wire N__23913;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23898;
    wire N__23893;
    wire N__23890;
    wire N__23889;
    wire N__23886;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23871;
    wire N__23866;
    wire N__23863;
    wire N__23862;
    wire N__23861;
    wire N__23860;
    wire N__23857;
    wire N__23850;
    wire N__23845;
    wire N__23844;
    wire N__23843;
    wire N__23842;
    wire N__23839;
    wire N__23834;
    wire N__23831;
    wire N__23826;
    wire N__23821;
    wire N__23818;
    wire N__23817;
    wire N__23816;
    wire N__23813;
    wire N__23808;
    wire N__23805;
    wire N__23800;
    wire N__23797;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23769;
    wire N__23766;
    wire N__23765;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23753;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23734;
    wire N__23731;
    wire N__23730;
    wire N__23729;
    wire N__23726;
    wire N__23721;
    wire N__23720;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23694;
    wire N__23691;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23679;
    wire N__23678;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23662;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23632;
    wire N__23631;
    wire N__23630;
    wire N__23629;
    wire N__23628;
    wire N__23627;
    wire N__23626;
    wire N__23625;
    wire N__23622;
    wire N__23621;
    wire N__23618;
    wire N__23617;
    wire N__23614;
    wire N__23613;
    wire N__23610;
    wire N__23609;
    wire N__23606;
    wire N__23605;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23597;
    wire N__23594;
    wire N__23579;
    wire N__23578;
    wire N__23577;
    wire N__23560;
    wire N__23557;
    wire N__23556;
    wire N__23553;
    wire N__23552;
    wire N__23551;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23541;
    wire N__23532;
    wire N__23531;
    wire N__23530;
    wire N__23529;
    wire N__23524;
    wire N__23517;
    wire N__23510;
    wire N__23503;
    wire N__23502;
    wire N__23501;
    wire N__23500;
    wire N__23499;
    wire N__23498;
    wire N__23497;
    wire N__23496;
    wire N__23495;
    wire N__23494;
    wire N__23493;
    wire N__23492;
    wire N__23489;
    wire N__23488;
    wire N__23485;
    wire N__23484;
    wire N__23483;
    wire N__23466;
    wire N__23465;
    wire N__23464;
    wire N__23461;
    wire N__23448;
    wire N__23445;
    wire N__23444;
    wire N__23443;
    wire N__23442;
    wire N__23441;
    wire N__23440;
    wire N__23439;
    wire N__23438;
    wire N__23433;
    wire N__23428;
    wire N__23425;
    wire N__23420;
    wire N__23411;
    wire N__23408;
    wire N__23395;
    wire N__23394;
    wire N__23393;
    wire N__23392;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23378;
    wire N__23377;
    wire N__23376;
    wire N__23375;
    wire N__23374;
    wire N__23371;
    wire N__23370;
    wire N__23369;
    wire N__23368;
    wire N__23367;
    wire N__23366;
    wire N__23365;
    wire N__23356;
    wire N__23347;
    wire N__23346;
    wire N__23345;
    wire N__23344;
    wire N__23341;
    wire N__23340;
    wire N__23339;
    wire N__23332;
    wire N__23323;
    wire N__23318;
    wire N__23315;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23307;
    wire N__23306;
    wire N__23301;
    wire N__23298;
    wire N__23293;
    wire N__23290;
    wire N__23285;
    wire N__23278;
    wire N__23275;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23241;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23229;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22890;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22819;
    wire N__22816;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22669;
    wire N__22666;
    wire N__22663;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22485;
    wire N__22482;
    wire N__22479;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22306;
    wire N__22303;
    wire N__22300;
    wire N__22297;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22200;
    wire N__22199;
    wire N__22198;
    wire N__22197;
    wire N__22194;
    wire N__22193;
    wire N__22190;
    wire N__22189;
    wire N__22186;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21985;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21955;
    wire N__21952;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21873;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21865;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21847;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21835;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21823;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21808;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21793;
    wire N__21792;
    wire N__21791;
    wire N__21790;
    wire N__21787;
    wire N__21786;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21760;
    wire N__21751;
    wire N__21750;
    wire N__21749;
    wire N__21748;
    wire N__21747;
    wire N__21746;
    wire N__21741;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21721;
    wire N__21720;
    wire N__21719;
    wire N__21718;
    wire N__21717;
    wire N__21716;
    wire N__21711;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21691;
    wire N__21690;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21658;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21594;
    wire N__21591;
    wire N__21588;
    wire N__21583;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21571;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21556;
    wire N__21553;
    wire N__21552;
    wire N__21549;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21532;
    wire N__21529;
    wire N__21528;
    wire N__21527;
    wire N__21526;
    wire N__21523;
    wire N__21522;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21514;
    wire N__21513;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21505;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21399;
    wire N__21396;
    wire N__21393;
    wire N__21388;
    wire N__21385;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21373;
    wire N__21370;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21358;
    wire N__21355;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21340;
    wire N__21337;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21301;
    wire N__21298;
    wire N__21297;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21250;
    wire N__21247;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21211;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21118;
    wire N__21115;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21097;
    wire N__21094;
    wire N__21093;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21078;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21055;
    wire N__21052;
    wire N__21051;
    wire N__21048;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21033;
    wire N__21030;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20994;
    wire N__20991;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20878;
    wire N__20875;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20860;
    wire N__20857;
    wire N__20854;
    wire N__20851;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20839;
    wire N__20836;
    wire N__20835;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20809;
    wire N__20806;
    wire N__20805;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20682;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20660;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20628;
    wire N__20625;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20607;
    wire N__20604;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20590;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20569;
    wire N__20566;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20326;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20316;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20293;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20212;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20136;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20107;
    wire N__20104;
    wire N__20103;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20007;
    wire N__20004;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19987;
    wire N__19986;
    wire N__19985;
    wire N__19982;
    wire N__19977;
    wire N__19974;
    wire N__19969;
    wire N__19968;
    wire N__19967;
    wire N__19964;
    wire N__19959;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19896;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19857;
    wire N__19854;
    wire N__19853;
    wire N__19852;
    wire N__19851;
    wire N__19850;
    wire N__19849;
    wire N__19848;
    wire N__19847;
    wire N__19846;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19828;
    wire N__19825;
    wire N__19818;
    wire N__19811;
    wire N__19810;
    wire N__19807;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19764;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19734;
    wire N__19733;
    wire N__19732;
    wire N__19731;
    wire N__19730;
    wire N__19729;
    wire N__19728;
    wire N__19727;
    wire N__19722;
    wire N__19717;
    wire N__19706;
    wire N__19705;
    wire N__19704;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19672;
    wire N__19671;
    wire N__19670;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19659;
    wire N__19658;
    wire N__19657;
    wire N__19656;
    wire N__19655;
    wire N__19654;
    wire N__19649;
    wire N__19644;
    wire N__19641;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19615;
    wire N__19614;
    wire N__19613;
    wire N__19612;
    wire N__19611;
    wire N__19610;
    wire N__19609;
    wire N__19608;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19587;
    wire N__19582;
    wire N__19581;
    wire N__19574;
    wire N__19569;
    wire N__19564;
    wire N__19561;
    wire N__19556;
    wire N__19553;
    wire N__19548;
    wire N__19545;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19299;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19282;
    wire N__19281;
    wire N__19278;
    wire N__19277;
    wire N__19276;
    wire N__19275;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19259;
    wire N__19258;
    wire N__19251;
    wire N__19248;
    wire N__19243;
    wire N__19240;
    wire N__19239;
    wire N__19236;
    wire N__19235;
    wire N__19234;
    wire N__19233;
    wire N__19232;
    wire N__19229;
    wire N__19218;
    wire N__19217;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19203;
    wire N__19194;
    wire N__19191;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19177;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19077;
    wire N__19076;
    wire N__19075;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19065;
    wire N__19064;
    wire N__19061;
    wire N__19060;
    wire N__19057;
    wire N__19056;
    wire N__19051;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19005;
    wire N__19004;
    wire N__19001;
    wire N__18996;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18981;
    wire N__18976;
    wire N__18975;
    wire N__18974;
    wire N__18971;
    wire N__18966;
    wire N__18965;
    wire N__18960;
    wire N__18957;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18943;
    wire N__18940;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18886;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18862;
    wire N__18859;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18553;
    wire N__18552;
    wire N__18551;
    wire N__18550;
    wire N__18549;
    wire N__18548;
    wire N__18547;
    wire N__18546;
    wire N__18545;
    wire N__18544;
    wire N__18543;
    wire N__18542;
    wire N__18541;
    wire N__18524;
    wire N__18519;
    wire N__18518;
    wire N__18517;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18487;
    wire N__18486;
    wire N__18485;
    wire N__18484;
    wire N__18483;
    wire N__18482;
    wire N__18481;
    wire N__18480;
    wire N__18471;
    wire N__18466;
    wire N__18463;
    wire N__18448;
    wire N__18445;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18423;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18340;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18319;
    wire N__18318;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18297;
    wire N__18292;
    wire N__18289;
    wire N__18288;
    wire N__18285;
    wire N__18282;
    wire N__18277;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18256;
    wire N__18253;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18243;
    wire N__18240;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18213;
    wire N__18212;
    wire N__18209;
    wire N__18204;
    wire N__18199;
    wire N__18196;
    wire N__18193;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18181;
    wire N__18178;
    wire N__18175;
    wire N__18174;
    wire N__18171;
    wire N__18170;
    wire N__18167;
    wire N__18162;
    wire N__18159;
    wire N__18154;
    wire N__18153;
    wire N__18152;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire GNDG0;
    wire VCCG0;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire pwm_duty_input_9;
    wire pwm_duty_input_5;
    wire pwm_duty_input_2;
    wire pwm_duty_input_3;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire \current_shift_inst.PI_CTRL.m14_2 ;
    wire \current_shift_inst.PI_CTRL.N_19_cascade_ ;
    wire pwm_duty_input_4;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire bfn_2_8_0_;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire bfn_2_9_0_;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire pwm_duty_input_8;
    wire pwm_duty_input_10;
    wire \current_shift_inst.PI_CTRL.m7_2 ;
    wire pwm_duty_input_7;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire bfn_2_12_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire bfn_2_13_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire bfn_2_14_0_;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire \current_shift_inst.PI_CTRL.N_98 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \current_shift_inst.PI_CTRL.N_178 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire N_22_i_i;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire pwm_duty_input_6;
    wire i8_mux;
    wire N_28_mux;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_3_9_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_3_10_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire bfn_3_11_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire bfn_3_12_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire bfn_3_13_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire bfn_3_14_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire clk_10khz_RNIIENAZ0Z2;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_4_17_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_4_18_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire bfn_4_19_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_4_20_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire un7_start_stop_0_a3;
    wire bfn_5_7_0_;
    wire un5_counter_cry_1;
    wire counterZ0Z_3;
    wire un5_counter_cry_2;
    wire counterZ0Z_4;
    wire un5_counter_cry_3;
    wire counterZ0Z_5;
    wire un5_counter_cry_4;
    wire counterZ0Z_6;
    wire un5_counter_cry_5;
    wire counter_RNO_0Z0Z_7;
    wire un5_counter_cry_6;
    wire un5_counter_cry_7;
    wire un5_counter_cry_8;
    wire bfn_5_8_0_;
    wire counter_RNO_0Z0Z_10;
    wire un5_counter_cry_9;
    wire un5_counter_cry_10;
    wire un5_counter_cry_11;
    wire counter_RNO_0Z0Z_12;
    wire counterZ0Z_10;
    wire counterZ0Z_7;
    wire counterZ0Z_2;
    wire counterZ0Z_1;
    wire un2_counter_5_cascade_;
    wire counterZ0Z_0;
    wire counterZ0Z_11;
    wire counterZ0Z_9;
    wire counterZ0Z_12;
    wire counterZ0Z_8;
    wire un2_counter_7;
    wire un2_counter_8;
    wire un2_counter_9;
    wire clk_10khz_i;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_5_13_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire bfn_5_14_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire bfn_5_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un1_enablelt3_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_7_13_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire bfn_7_14_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ;
    wire bfn_7_15_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire \current_shift_inst.PI_CTRL.N_47_16_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31 ;
    wire \current_shift_inst.PI_CTRL.N_47_21 ;
    wire \current_shift_inst.PI_CTRL.N_47_16 ;
    wire \current_shift_inst.PI_CTRL.N_47_21_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2 ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_44 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.timer_s1.N_187_i ;
    wire il_max_comp1_c;
    wire il_max_comp1_D1;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ;
    wire \phase_controller_inst1.N_228_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire bfn_8_17_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire bfn_8_18_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire bfn_8_19_0_;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire bfn_8_20_0_;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.N_199 ;
    wire \current_shift_inst.phase_validZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3 ;
    wire measured_delay_hc_21;
    wire measured_delay_hc_20;
    wire measured_delay_hc_22;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt8_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt15 ;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_9_11_0_;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_9_12_0_;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.time_passed11 ;
    wire \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.N_46_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.N_75 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_76 ;
    wire N_717_g;
    wire \current_shift_inst.meas_stateZ0Z_0 ;
    wire \current_shift_inst.S3_riseZ0 ;
    wire \current_shift_inst.S3_syncZ0Z0 ;
    wire \current_shift_inst.S3_syncZ0Z1 ;
    wire \current_shift_inst.S3_sync_prevZ0 ;
    wire il_min_comp2_c;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4 ;
    wire \delay_measurement_inst.prev_hc_sigZ0 ;
    wire \delay_measurement_inst.hc_stateZ0Z_0 ;
    wire delay_hc_d2;
    wire measured_delay_hc_26;
    wire measured_delay_hc_30;
    wire measured_delay_hc_25;
    wire measured_delay_hc_23;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire measured_delay_hc_24;
    wire measured_delay_hc_29;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto13 ;
    wire measured_delay_hc_19;
    wire \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ;
    wire bfn_10_12_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_10_13_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \phase_controller_inst1.N_232_cascade_ ;
    wire il_max_comp1_D2;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_46_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ;
    wire \phase_controller_inst1.stoper_tr.N_21_cascade_ ;
    wire bfn_10_21_0_;
    wire \current_shift_inst.z_i_0_31 ;
    wire \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ;
    wire \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_0 ;
    wire \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_1 ;
    wire \current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_2 ;
    wire \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_3 ;
    wire \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ;
    wire \current_shift_inst.un38_control_input_0_cry_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ;
    wire \current_shift_inst.un38_control_input_0_cry_5 ;
    wire \current_shift_inst.un38_control_input_0_cry_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ;
    wire bfn_10_22_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ;
    wire \current_shift_inst.un38_control_input_0_cry_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ;
    wire \current_shift_inst.un38_control_input_0_cry_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ;
    wire \current_shift_inst.un38_control_input_0_cry_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ;
    wire \current_shift_inst.un38_control_input_0_cry_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNILORI_11 ;
    wire \current_shift_inst.un38_control_input_0_cry_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ;
    wire \current_shift_inst.un38_control_input_0_cry_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ;
    wire \current_shift_inst.un38_control_input_0_cry_13 ;
    wire \current_shift_inst.un38_control_input_0_cry_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ;
    wire bfn_10_23_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI190J_15 ;
    wire \current_shift_inst.un38_control_input_0_cry_15 ;
    wire \current_shift_inst.un38_control_input_0_cry_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ;
    wire \current_shift_inst.un38_control_input_0_cry_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ;
    wire \current_shift_inst.un38_control_input_0_cry_18 ;
    wire \current_shift_inst.un38_control_input_0_cry_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ;
    wire \current_shift_inst.un38_control_input_0_cry_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ;
    wire \current_shift_inst.un38_control_input_0_cry_21 ;
    wire \current_shift_inst.un38_control_input_0_cry_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ;
    wire bfn_10_24_0_;
    wire \current_shift_inst.un38_control_input_0_cry_23 ;
    wire \current_shift_inst.un38_control_input_0_cry_24 ;
    wire \current_shift_inst.un38_control_input_0_cry_25 ;
    wire \current_shift_inst.un38_control_input_0_cry_26 ;
    wire \current_shift_inst.un38_control_input_0_cry_27 ;
    wire \current_shift_inst.un38_control_input_0_cry_28 ;
    wire \current_shift_inst.un38_control_input_0_cry_29 ;
    wire \current_shift_inst.un38_control_input_0_cry_30 ;
    wire bfn_10_25_0_;
    wire \current_shift_inst.control_inputZ0Z_25 ;
    wire il_max_comp2_c;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_336_i ;
    wire measured_delay_hc_27;
    wire measured_delay_hc_28;
    wire il_min_comp1_c;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.un1_counterlto9_2_cascade_ ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.un1_counterlt9 ;
    wire il_min_comp1_D1;
    wire \phase_controller_inst1.N_231 ;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire \current_shift_inst.S1_riseZ0 ;
    wire \current_shift_inst.S1_syncZ0Z0 ;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire \current_shift_inst.S1_syncZ0Z1 ;
    wire \current_shift_inst.S1_sync_prevZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ;
    wire \current_shift_inst.control_input_1_axb_0 ;
    wire \current_shift_inst.control_inputZ0Z_0 ;
    wire bfn_11_20_0_;
    wire \current_shift_inst.control_input_1_axb_1 ;
    wire \current_shift_inst.control_inputZ0Z_1 ;
    wire \current_shift_inst.control_input_1_cry_0 ;
    wire \current_shift_inst.control_input_1_axb_2 ;
    wire \current_shift_inst.control_inputZ0Z_2 ;
    wire \current_shift_inst.control_input_1_cry_1 ;
    wire \current_shift_inst.control_input_1_axb_3 ;
    wire \current_shift_inst.control_inputZ0Z_3 ;
    wire \current_shift_inst.control_input_1_cry_2 ;
    wire \current_shift_inst.control_input_1_axb_4 ;
    wire \current_shift_inst.control_inputZ0Z_4 ;
    wire \current_shift_inst.control_input_1_cry_3 ;
    wire \current_shift_inst.control_input_1_axb_5 ;
    wire \current_shift_inst.control_inputZ0Z_5 ;
    wire \current_shift_inst.control_input_1_cry_4 ;
    wire \current_shift_inst.control_input_1_axb_6 ;
    wire \current_shift_inst.control_inputZ0Z_6 ;
    wire \current_shift_inst.control_input_1_cry_5 ;
    wire \current_shift_inst.control_input_1_axb_7 ;
    wire \current_shift_inst.control_inputZ0Z_7 ;
    wire \current_shift_inst.control_input_1_cry_6 ;
    wire \current_shift_inst.control_input_1_cry_7 ;
    wire \current_shift_inst.control_input_1_axb_8 ;
    wire \current_shift_inst.control_inputZ0Z_8 ;
    wire bfn_11_21_0_;
    wire \current_shift_inst.control_input_1_axb_9 ;
    wire \current_shift_inst.control_inputZ0Z_9 ;
    wire \current_shift_inst.control_input_1_cry_8 ;
    wire \current_shift_inst.control_input_1_axb_10 ;
    wire \current_shift_inst.control_inputZ0Z_10 ;
    wire \current_shift_inst.control_input_1_cry_9 ;
    wire \current_shift_inst.control_input_1_axb_11 ;
    wire \current_shift_inst.control_inputZ0Z_11 ;
    wire \current_shift_inst.control_input_1_cry_10 ;
    wire \current_shift_inst.control_input_1_axb_12 ;
    wire \current_shift_inst.control_inputZ0Z_12 ;
    wire \current_shift_inst.control_input_1_cry_11 ;
    wire \current_shift_inst.control_input_1_axb_13 ;
    wire \current_shift_inst.control_inputZ0Z_13 ;
    wire \current_shift_inst.control_input_1_cry_12 ;
    wire \current_shift_inst.control_input_1_axb_14 ;
    wire \current_shift_inst.control_inputZ0Z_14 ;
    wire \current_shift_inst.control_input_1_cry_13 ;
    wire \current_shift_inst.control_input_1_axb_15 ;
    wire \current_shift_inst.control_inputZ0Z_15 ;
    wire \current_shift_inst.control_input_1_cry_14 ;
    wire \current_shift_inst.control_input_1_cry_15 ;
    wire \current_shift_inst.control_input_1_axb_16 ;
    wire \current_shift_inst.control_inputZ0Z_16 ;
    wire bfn_11_22_0_;
    wire \current_shift_inst.control_input_1_axb_17 ;
    wire \current_shift_inst.control_inputZ0Z_17 ;
    wire \current_shift_inst.control_input_1_cry_16 ;
    wire \current_shift_inst.control_input_1_axb_18 ;
    wire \current_shift_inst.control_inputZ0Z_18 ;
    wire \current_shift_inst.control_input_1_cry_17 ;
    wire \current_shift_inst.control_input_1_axb_19 ;
    wire \current_shift_inst.control_inputZ0Z_19 ;
    wire \current_shift_inst.control_input_1_cry_18 ;
    wire \current_shift_inst.control_input_1_axb_20 ;
    wire \current_shift_inst.control_inputZ0Z_20 ;
    wire \current_shift_inst.control_input_1_cry_19 ;
    wire \current_shift_inst.control_input_1_axb_21 ;
    wire \current_shift_inst.control_inputZ0Z_21 ;
    wire \current_shift_inst.control_input_1_cry_20 ;
    wire \current_shift_inst.control_input_1_axb_22 ;
    wire \current_shift_inst.control_inputZ0Z_22 ;
    wire \current_shift_inst.control_input_1_cry_21 ;
    wire \current_shift_inst.control_input_1_axb_23 ;
    wire \current_shift_inst.control_inputZ0Z_23 ;
    wire \current_shift_inst.control_input_1_cry_22 ;
    wire \current_shift_inst.control_input_1_cry_23 ;
    wire \current_shift_inst.control_input_1_axb_24 ;
    wire \current_shift_inst.control_inputZ0Z_24 ;
    wire bfn_11_23_0_;
    wire \current_shift_inst.phase_valid_RNISLORZ0Z2 ;
    wire \current_shift_inst.control_input_1_cry_24 ;
    wire \current_shift_inst.control_input_1_cry_24_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ;
    wire \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_ ;
    wire \delay_measurement_inst.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.elapsed_time_hc_2 ;
    wire bfn_12_7_0_;
    wire \delay_measurement_inst.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_reg3lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_reg3lto9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_11 ;
    wire bfn_12_8_0_;
    wire \delay_measurement_inst.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_reg3lto15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.elapsed_time_hc_19 ;
    wire bfn_12_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_12_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.N_336_i_g ;
    wire \delay_measurement_inst.elapsed_time_hc_16 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire il_min_comp1_D2;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire s1_phy_c;
    wire \phase_controller_inst1.stoper_tr.N_21 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3 ;
    wire \current_shift_inst.z_i_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ;
    wire \current_shift_inst.timer_phase.N_188_i ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire bfn_12_24_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ;
    wire bfn_12_25_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_12_26_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_reg3lto14 ;
    wire \delay_measurement_inst.delay_hc_reg3 ;
    wire \delay_measurement_inst.elapsed_time_hc_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_13_7_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_13_8_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_13_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_13_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_337_i ;
    wire start_stop_c;
    wire red_c_i;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ;
    wire \current_shift_inst.un38_control_input_0_axb_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ;
    wire \current_shift_inst.start_timer_phaseZ0 ;
    wire \current_shift_inst.stop_timer_phaseZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ;
    wire \current_shift_inst.timer_phase.runningZ0 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_13_21_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_13_22_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_13_23_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire s2_phy_c;
    wire \delay_measurement_inst.un1_elapsed_time_hc ;
    wire \delay_measurement_inst.delay_hc_reg3lto31_0_0 ;
    wire measured_delay_hc_12;
    wire measured_delay_hc_14;
    wire measured_delay_hc_16;
    wire measured_delay_hc_17;
    wire measured_delay_hc_18;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ;
    wire \phase_controller_slave.stoper_tr.time_passed11_cascade_ ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire bfn_14_11_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_14_12_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_14_13_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.un4_control_input_axb_1 ;
    wire bfn_14_14_0_;
    wire \current_shift_inst.un4_control_input_axb_2 ;
    wire \current_shift_inst.un4_control_input_cry_1 ;
    wire \current_shift_inst.un4_control_input_axb_3 ;
    wire \current_shift_inst.un4_control_input_cry_2 ;
    wire \current_shift_inst.un4_control_input_cry_3 ;
    wire \current_shift_inst.un4_control_input_cry_4 ;
    wire \current_shift_inst.un4_control_input_cry_5 ;
    wire \current_shift_inst.un4_control_input_cry_6 ;
    wire \current_shift_inst.un4_control_input_cry_7 ;
    wire \current_shift_inst.un4_control_input_cry_8 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.un4_control_input_cry_9 ;
    wire \current_shift_inst.un4_control_input_cry_10 ;
    wire \current_shift_inst.un4_control_input_cry_11 ;
    wire \current_shift_inst.un4_control_input_cry_12 ;
    wire \current_shift_inst.un4_control_input_cry_13 ;
    wire \current_shift_inst.un4_control_input_cry_14 ;
    wire \current_shift_inst.un4_control_input_cry_15 ;
    wire \current_shift_inst.un4_control_input_cry_16 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.un4_control_input_cry_17 ;
    wire \current_shift_inst.un4_control_input_cry_18 ;
    wire \current_shift_inst.un4_control_input_cry_19 ;
    wire \current_shift_inst.un4_control_input_cry_20 ;
    wire \current_shift_inst.un4_control_input_cry_21 ;
    wire \current_shift_inst.un4_control_input_cry_22 ;
    wire \current_shift_inst.un4_control_input_cry_23 ;
    wire \current_shift_inst.un4_control_input_cry_24 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.un4_control_input_cry_25 ;
    wire \current_shift_inst.un4_control_input_cry_26 ;
    wire \current_shift_inst.un4_control_input_cry_27 ;
    wire \current_shift_inst.un4_control_input_cry_28 ;
    wire \current_shift_inst.un4_control_input_cry_29 ;
    wire \current_shift_inst.un4_control_input_cry_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ;
    wire \current_shift_inst.un38_control_input_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_fast_31 ;
    wire G_407;
    wire bfn_14_18_0_;
    wire \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ;
    wire G_406;
    wire \current_shift_inst.z_cry_0 ;
    wire \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ;
    wire \current_shift_inst.z_cry_1 ;
    wire \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ;
    wire \current_shift_inst.z_cry_2 ;
    wire \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ;
    wire \current_shift_inst.z_cry_3 ;
    wire \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ;
    wire \current_shift_inst.z_cry_4 ;
    wire \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ;
    wire \current_shift_inst.z_cry_5 ;
    wire \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ;
    wire \current_shift_inst.z_cry_6 ;
    wire \current_shift_inst.z_cry_7 ;
    wire \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ;
    wire bfn_14_19_0_;
    wire \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ;
    wire \current_shift_inst.z_cry_8 ;
    wire \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ;
    wire \current_shift_inst.z_cry_9 ;
    wire \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ;
    wire \current_shift_inst.z_cry_10 ;
    wire \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ;
    wire \current_shift_inst.z_cry_11 ;
    wire \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ;
    wire \current_shift_inst.z_cry_12 ;
    wire \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ;
    wire \current_shift_inst.z_cry_13 ;
    wire \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ;
    wire \current_shift_inst.z_cry_14 ;
    wire \current_shift_inst.z_cry_15 ;
    wire \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ;
    wire bfn_14_20_0_;
    wire \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ;
    wire \current_shift_inst.z_cry_16 ;
    wire \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ;
    wire \current_shift_inst.z_cry_17 ;
    wire \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ;
    wire \current_shift_inst.z_cry_18 ;
    wire \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ;
    wire \current_shift_inst.z_cry_19 ;
    wire \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ;
    wire \current_shift_inst.z_cry_20 ;
    wire \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ;
    wire \current_shift_inst.z_cry_21 ;
    wire \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ;
    wire \current_shift_inst.z_cry_22 ;
    wire \current_shift_inst.z_cry_23 ;
    wire \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ;
    wire bfn_14_21_0_;
    wire \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ;
    wire \current_shift_inst.z_cry_24 ;
    wire \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ;
    wire \current_shift_inst.z_cry_25 ;
    wire \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ;
    wire \current_shift_inst.z_cry_26 ;
    wire \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ;
    wire \current_shift_inst.z_cry_27 ;
    wire \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ;
    wire \current_shift_inst.z_cry_28 ;
    wire \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ;
    wire \current_shift_inst.z_cry_29 ;
    wire \current_shift_inst.z_cry_30 ;
    wire \current_shift_inst.z_31 ;
    wire bfn_14_22_0_;
    wire \current_shift_inst.timer_phase.counter_cry_0 ;
    wire \current_shift_inst.timer_phase.counter_cry_1 ;
    wire \current_shift_inst.timer_phase.counter_cry_2 ;
    wire \current_shift_inst.timer_phase.counter_cry_3 ;
    wire \current_shift_inst.timer_phase.counter_cry_4 ;
    wire \current_shift_inst.timer_phase.counter_cry_5 ;
    wire \current_shift_inst.timer_phase.counter_cry_6 ;
    wire \current_shift_inst.timer_phase.counter_cry_7 ;
    wire bfn_14_23_0_;
    wire \current_shift_inst.timer_phase.counter_cry_8 ;
    wire \current_shift_inst.timer_phase.counter_cry_9 ;
    wire \current_shift_inst.timer_phase.counter_cry_10 ;
    wire \current_shift_inst.timer_phase.counter_cry_11 ;
    wire \current_shift_inst.timer_phase.counter_cry_12 ;
    wire \current_shift_inst.timer_phase.counter_cry_13 ;
    wire \current_shift_inst.timer_phase.counter_cry_14 ;
    wire \current_shift_inst.timer_phase.counter_cry_15 ;
    wire bfn_14_24_0_;
    wire \current_shift_inst.timer_phase.counter_cry_16 ;
    wire \current_shift_inst.timer_phase.counter_cry_17 ;
    wire \current_shift_inst.timer_phase.counter_cry_18 ;
    wire \current_shift_inst.timer_phase.counter_cry_19 ;
    wire \current_shift_inst.timer_phase.counter_cry_20 ;
    wire \current_shift_inst.timer_phase.counter_cry_21 ;
    wire \current_shift_inst.timer_phase.counter_cry_22 ;
    wire \current_shift_inst.timer_phase.counter_cry_23 ;
    wire bfn_14_25_0_;
    wire \current_shift_inst.timer_phase.counter_cry_24 ;
    wire \current_shift_inst.timer_phase.counter_cry_25 ;
    wire \current_shift_inst.timer_phase.counter_cry_26 ;
    wire \current_shift_inst.timer_phase.counter_cry_27 ;
    wire \current_shift_inst.timer_phase.running_i ;
    wire \current_shift_inst.timer_phase.counter_cry_28 ;
    wire \current_shift_inst.timer_phase.N_192_i ;
    wire delay_tr_input_c;
    wire delay_tr_d1;
    wire measured_delay_hc_7;
    wire measured_delay_hc_2;
    wire measured_delay_hc_6;
    wire measured_delay_hc_4;
    wire measured_delay_hc_5;
    wire measured_delay_hc_3;
    wire measured_delay_hc_13;
    wire measured_delay_hc_9;
    wire measured_delay_hc_10;
    wire measured_delay_hc_11;
    wire measured_delay_hc_0;
    wire \phase_controller_inst1.stoper_hc.un2_startlt31 ;
    wire measured_delay_hc_1;
    wire measured_delay_hc_15;
    wire \phase_controller_inst1.stoper_hc.un1_startlt31_0 ;
    wire measured_delay_hc_8;
    wire measured_delay_hc_31;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_ ;
    wire measured_delay_tr_14;
    wire \current_shift_inst.un4_control_input_axb_4 ;
    wire \current_shift_inst.un4_control_input_axb_5 ;
    wire \current_shift_inst.un4_control_input_axb_6 ;
    wire \current_shift_inst.un4_control_input_axb_7 ;
    wire \current_shift_inst.un4_control_input_axb_8 ;
    wire \current_shift_inst.un4_control_input_axb_9 ;
    wire \current_shift_inst.un4_control_input_axb_10 ;
    wire \current_shift_inst.un4_control_input_axb_11 ;
    wire \current_shift_inst.un4_control_input_axb_22 ;
    wire \current_shift_inst.un4_control_input_axb_12 ;
    wire \current_shift_inst.un4_control_input_axb_19 ;
    wire \current_shift_inst.un4_control_input_axb_17 ;
    wire \current_shift_inst.un4_control_input_axb_15 ;
    wire \current_shift_inst.un4_control_input_axb_16 ;
    wire \current_shift_inst.un4_control_input_axb_18 ;
    wire \current_shift_inst.un4_control_input_axb_23 ;
    wire \current_shift_inst.un4_control_input_axb_27 ;
    wire \current_shift_inst.un4_control_input_axb_20 ;
    wire \current_shift_inst.un4_control_input_axb_30 ;
    wire \current_shift_inst.un4_control_input_axb_26 ;
    wire \current_shift_inst.un4_control_input_axb_29 ;
    wire \current_shift_inst.un4_control_input_axb_28 ;
    wire \current_shift_inst.un4_control_input_axb_25 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \current_shift_inst.un4_control_input_axb_21 ;
    wire \current_shift_inst.un4_control_input_axb_13 ;
    wire measured_delay_tr_12;
    wire measured_delay_tr_13;
    wire measured_delay_tr_11;
    wire measured_delay_tr_10;
    wire \current_shift_inst.N_1742_i ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ;
    wire \current_shift_inst.elapsed_time_ns_phase_1 ;
    wire bfn_15_21_0_;
    wire \current_shift_inst.elapsed_time_ns_phase_2 ;
    wire \current_shift_inst.z_5_2 ;
    wire \current_shift_inst.z_5_cry_1 ;
    wire \current_shift_inst.z_5_3 ;
    wire \current_shift_inst.z_5_cry_2 ;
    wire \current_shift_inst.z_5_4 ;
    wire \current_shift_inst.z_5_cry_3 ;
    wire \current_shift_inst.z_5_5 ;
    wire \current_shift_inst.z_5_cry_4 ;
    wire \current_shift_inst.z_5_6 ;
    wire \current_shift_inst.z_5_cry_5 ;
    wire \current_shift_inst.z_5_7 ;
    wire \current_shift_inst.z_5_cry_6 ;
    wire \current_shift_inst.z_5_8 ;
    wire \current_shift_inst.z_5_cry_7 ;
    wire \current_shift_inst.z_5_cry_8 ;
    wire \current_shift_inst.z_5_9 ;
    wire bfn_15_22_0_;
    wire \current_shift_inst.z_5_10 ;
    wire \current_shift_inst.z_5_cry_9 ;
    wire \current_shift_inst.z_5_11 ;
    wire \current_shift_inst.z_5_cry_10 ;
    wire \current_shift_inst.z_5_12 ;
    wire \current_shift_inst.z_5_cry_11 ;
    wire \current_shift_inst.z_5_13 ;
    wire \current_shift_inst.z_5_cry_12 ;
    wire \current_shift_inst.z_5_14 ;
    wire \current_shift_inst.z_5_cry_13 ;
    wire \current_shift_inst.z_5_15 ;
    wire \current_shift_inst.z_5_cry_14 ;
    wire \current_shift_inst.z_5_16 ;
    wire \current_shift_inst.z_5_cry_15 ;
    wire \current_shift_inst.z_5_cry_16 ;
    wire \current_shift_inst.z_5_17 ;
    wire bfn_15_23_0_;
    wire \current_shift_inst.z_5_18 ;
    wire \current_shift_inst.z_5_cry_17 ;
    wire \current_shift_inst.z_5_19 ;
    wire \current_shift_inst.z_5_cry_18 ;
    wire \current_shift_inst.z_5_20 ;
    wire \current_shift_inst.z_5_cry_19 ;
    wire \current_shift_inst.z_5_21 ;
    wire \current_shift_inst.z_5_cry_20 ;
    wire \current_shift_inst.z_5_22 ;
    wire \current_shift_inst.z_5_cry_21 ;
    wire \current_shift_inst.z_5_23 ;
    wire \current_shift_inst.z_5_cry_22 ;
    wire \current_shift_inst.z_5_24 ;
    wire \current_shift_inst.z_5_cry_23 ;
    wire \current_shift_inst.z_5_cry_24 ;
    wire \current_shift_inst.z_5_25 ;
    wire bfn_15_24_0_;
    wire \current_shift_inst.z_5_26 ;
    wire \current_shift_inst.z_5_cry_25 ;
    wire \current_shift_inst.z_5_27 ;
    wire \current_shift_inst.z_5_cry_26 ;
    wire \current_shift_inst.z_5_28 ;
    wire \current_shift_inst.z_5_cry_27 ;
    wire \current_shift_inst.z_5_29 ;
    wire \current_shift_inst.z_5_cry_28 ;
    wire \current_shift_inst.z_5_30 ;
    wire \current_shift_inst.z_5_cry_29 ;
    wire \current_shift_inst.z_5_cry_30 ;
    wire \current_shift_inst.z_5_cry_30_THRU_CO ;
    wire delay_hc_input_c;
    wire delay_hc_d1;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_16_8_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_8 ;
    wire bfn_16_9_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_16 ;
    wire bfn_16_10_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_1 ;
    wire bfn_16_11_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_9 ;
    wire bfn_16_12_0_;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_17 ;
    wire bfn_16_13_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ;
    wire measured_delay_tr_1;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_3 ;
    wire measured_delay_tr_9;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ;
    wire measured_delay_tr_3;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_20_li ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_2 ;
    wire measured_delay_tr_8;
    wire measured_delay_tr_7;
    wire measured_delay_tr_6;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6 ;
    wire measured_delay_tr_15;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ;
    wire measured_delay_tr_5;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_ ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_5 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ;
    wire bfn_16_15_0_;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ;
    wire bfn_16_16_0_;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ;
    wire bfn_16_17_0_;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ;
    wire bfn_16_18_0_;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.N_187_i_g ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire measured_delay_tr_18;
    wire measured_delay_tr_17;
    wire measured_delay_tr_19;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_3 ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.N_221_0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_424_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_3 ;
    wire bfn_16_22_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_1 ;
    wire \current_shift_inst.elapsed_time_ns_phase_4 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_2 ;
    wire \current_shift_inst.elapsed_time_ns_phase_5 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_3 ;
    wire \current_shift_inst.elapsed_time_ns_phase_6 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_4 ;
    wire \current_shift_inst.elapsed_time_ns_phase_7 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_5 ;
    wire \current_shift_inst.elapsed_time_ns_phase_8 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_6 ;
    wire \current_shift_inst.elapsed_time_ns_phase_9 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_7 ;
    wire \current_shift_inst.elapsed_time_ns_phase_10 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_8 ;
    wire \current_shift_inst.elapsed_time_ns_phase_11 ;
    wire bfn_16_23_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_9 ;
    wire \current_shift_inst.elapsed_time_ns_phase_12 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_10 ;
    wire \current_shift_inst.elapsed_time_ns_phase_13 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_11 ;
    wire \current_shift_inst.elapsed_time_ns_phase_14 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_12 ;
    wire \current_shift_inst.elapsed_time_ns_phase_15 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_13 ;
    wire \current_shift_inst.elapsed_time_ns_phase_16 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_14 ;
    wire \current_shift_inst.elapsed_time_ns_phase_17 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_15 ;
    wire \current_shift_inst.elapsed_time_ns_phase_18 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_16 ;
    wire \current_shift_inst.elapsed_time_ns_phase_19 ;
    wire bfn_16_24_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_17 ;
    wire \current_shift_inst.elapsed_time_ns_phase_20 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_18 ;
    wire \current_shift_inst.elapsed_time_ns_phase_21 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_19 ;
    wire \current_shift_inst.elapsed_time_ns_phase_22 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_20 ;
    wire \current_shift_inst.elapsed_time_ns_phase_23 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_21 ;
    wire \current_shift_inst.elapsed_time_ns_phase_24 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_22 ;
    wire \current_shift_inst.elapsed_time_ns_phase_25 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_23 ;
    wire \current_shift_inst.elapsed_time_ns_phase_26 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_24 ;
    wire \current_shift_inst.elapsed_time_ns_phase_27 ;
    wire bfn_16_25_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_25 ;
    wire \current_shift_inst.elapsed_time_ns_phase_28 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_28 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_26 ;
    wire \current_shift_inst.elapsed_time_ns_phase_29 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_27 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_29 ;
    wire \current_shift_inst.elapsed_time_ns_phase_30 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.elapsed_time_ns_phase_31 ;
    wire \current_shift_inst.timer_phase.N_188_i_g ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19 ;
    wire il_max_comp2_D1;
    wire il_min_comp2_D1;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_slave.N_214_cascade_ ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.start_timer_hcZ0 ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_slave.stoper_hc.time_passed11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_17_11_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_17_12_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_17_13_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_17_14_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_191_i ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un4_control_input_axb_14 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input_axb_24 ;
    wire CONSTANT_ONE_NET;
    wire \delay_measurement_inst.tr_stateZ0Z_0 ;
    wire delay_tr_d2;
    wire \delay_measurement_inst.prev_tr_sigZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_ ;
    wire \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_390_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_379 ;
    wire \delay_measurement_inst.N_280_i ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_ ;
    wire \delay_measurement_inst.N_409_1 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire bfn_17_23_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_17_24_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_17_25_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_17_26_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_339_i ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_18_8_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ;
    wire bfn_18_9_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ;
    wire bfn_18_10_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ;
    wire \phase_controller_slave.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_slave.hc_time_passed ;
    wire \phase_controller_slave.stateZ0Z_2 ;
    wire s4_phy_c;
    wire \phase_controller_slave.stateZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.time_passed11 ;
    wire \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_ ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire il_max_comp2_D2;
    wire \phase_controller_slave.N_213 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stateZ0Z_3 ;
    wire shift_flag_start;
    wire s3_phy_c;
    wire \phase_controller_slave.start_timer_trZ0 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ;
    wire measured_delay_tr_16;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ;
    wire measured_delay_tr_4;
    wire \delay_measurement_inst.N_425 ;
    wire \delay_measurement_inst.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ;
    wire measured_delay_tr_2;
    wire \delay_measurement_inst.N_280_i_0 ;
    wire \delay_measurement_inst.N_286_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_415 ;
    wire \delay_measurement_inst.N_373 ;
    wire \delay_measurement_inst.elapsed_time_tr_3 ;
    wire bfn_18_23_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.elapsed_time_tr_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.elapsed_time_tr_11 ;
    wire bfn_18_24_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.elapsed_time_tr_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.elapsed_time_tr_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire \delay_measurement_inst.elapsed_time_tr_19 ;
    wire bfn_18_25_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_18_26_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \phase_controller_slave.stateZ0Z_1 ;
    wire il_min_comp2_D2;
    wire \phase_controller_slave.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_slave.tr_time_passed ;
    wire \phase_controller_slave.stateZ0Z_0 ;
    wire \phase_controller_slave.N_211 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_tr_1 ;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire \delay_measurement_inst.delay_tr_timer.N_338_i ;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__20536),
            .RESETB(N__31431),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__43473),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__43335),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__18516,N__18544,N__18517,N__18545,N__18518,N__18174,N__18582,N__18423,N__19705,N__18152,N__18239,N__18319,N__18330,N__18277,N__18288}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__43341,N__43338,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__43336,N__43340,N__43337,N__43339}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__43501),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__43494),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64}),
            .ADDSUBBOT(),
            .A({dangling_wire_65,N__18552,N__18486,N__18550,N__18485,N__18551,N__18484,N__18553,N__18481,N__18546,N__18480,N__18547,N__18482,N__18548,N__18483,N__18549}),
            .C({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .B({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,N__43500,N__43497,dangling_wire_89,dangling_wire_90,dangling_wire_91,N__43495,N__43499,N__43496,N__43498}),
            .OHOLDTOP(),
            .O({dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__49352),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__49354),
            .DIN(N__49353),
            .DOUT(N__49352),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__49354),
            .PADOUT(N__49353),
            .PADIN(N__49352),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__49343),
            .DIN(N__49342),
            .DOUT(N__49341),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__49343),
            .PADOUT(N__49342),
            .PADIN(N__49341),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__49334),
            .DIN(N__49333),
            .DOUT(N__49332),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__49334),
            .PADOUT(N__49333),
            .PADIN(N__49332),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__49325),
            .DIN(N__49324),
            .DOUT(N__49323),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__49325),
            .PADOUT(N__49324),
            .PADIN(N__49323),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24697),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__49316),
            .DIN(N__49315),
            .DOUT(N__49314),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__49316),
            .PADOUT(N__49315),
            .PADIN(N__49314),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__49307),
            .DIN(N__49306),
            .DOUT(N__49305),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__49307),
            .PADOUT(N__49306),
            .PADIN(N__49305),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33664),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_iopad (
            .OE(N__49298),
            .DIN(N__49297),
            .DOUT(N__49296),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_preio (
            .PADOEN(N__49298),
            .PADOUT(N__49297),
            .PADIN(N__49296),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_iopad (
            .OE(N__49289),
            .DIN(N__49288),
            .DOUT(N__49287),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_preio (
            .PADOEN(N__49289),
            .PADOUT(N__49288),
            .PADIN(N__49287),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__49280),
            .DIN(N__49279),
            .DOUT(N__49278),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__49280),
            .PADOUT(N__49279),
            .PADIN(N__49278),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__49271),
            .DIN(N__49270),
            .DOUT(N__49269),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__49271),
            .PADOUT(N__49270),
            .PADIN(N__49269),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__30046),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__49262),
            .DIN(N__49261),
            .DOUT(N__49260),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__49262),
            .PADOUT(N__49261),
            .PADIN(N__49260),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44785),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__49253),
            .DIN(N__49252),
            .DOUT(N__49251),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__49253),
            .PADOUT(N__49252),
            .PADIN(N__49251),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__49244),
            .DIN(N__49243),
            .DOUT(N__49242),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__49244),
            .PADOUT(N__49243),
            .PADIN(N__49242),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__45691),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11881 (
            .O(N__49225),
            .I(N__49221));
    InMux I__11880 (
            .O(N__49224),
            .I(N__49218));
    LocalMux I__11879 (
            .O(N__49221),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__11878 (
            .O(N__49218),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__11877 (
            .O(N__49213),
            .I(N__49208));
    CascadeMux I__11876 (
            .O(N__49212),
            .I(N__49205));
    InMux I__11875 (
            .O(N__49211),
            .I(N__49202));
    InMux I__11874 (
            .O(N__49208),
            .I(N__49197));
    InMux I__11873 (
            .O(N__49205),
            .I(N__49197));
    LocalMux I__11872 (
            .O(N__49202),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__11871 (
            .O(N__49197),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__11870 (
            .O(N__49192),
            .I(N__49189));
    LocalMux I__11869 (
            .O(N__49189),
            .I(N__49186));
    Span4Mux_v I__11868 (
            .O(N__49186),
            .I(N__49183));
    Odrv4 I__11867 (
            .O(N__49183),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__11866 (
            .O(N__49180),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__11865 (
            .O(N__49177),
            .I(N__49173));
    InMux I__11864 (
            .O(N__49176),
            .I(N__49170));
    LocalMux I__11863 (
            .O(N__49173),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__11862 (
            .O(N__49170),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__11861 (
            .O(N__49165),
            .I(N__49160));
    CascadeMux I__11860 (
            .O(N__49164),
            .I(N__49157));
    InMux I__11859 (
            .O(N__49163),
            .I(N__49154));
    InMux I__11858 (
            .O(N__49160),
            .I(N__49149));
    InMux I__11857 (
            .O(N__49157),
            .I(N__49149));
    LocalMux I__11856 (
            .O(N__49154),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__11855 (
            .O(N__49149),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__11854 (
            .O(N__49144),
            .I(N__49141));
    LocalMux I__11853 (
            .O(N__49141),
            .I(N__49138));
    Span4Mux_v I__11852 (
            .O(N__49138),
            .I(N__49135));
    Odrv4 I__11851 (
            .O(N__49135),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ));
    InMux I__11850 (
            .O(N__49132),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__11849 (
            .O(N__49129),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__11848 (
            .O(N__49126),
            .I(N__49121));
    InMux I__11847 (
            .O(N__49125),
            .I(N__49116));
    InMux I__11846 (
            .O(N__49124),
            .I(N__49116));
    LocalMux I__11845 (
            .O(N__49121),
            .I(N__49111));
    LocalMux I__11844 (
            .O(N__49116),
            .I(N__49108));
    InMux I__11843 (
            .O(N__49115),
            .I(N__49105));
    CascadeMux I__11842 (
            .O(N__49114),
            .I(N__49096));
    Span4Mux_h I__11841 (
            .O(N__49111),
            .I(N__49088));
    Span4Mux_h I__11840 (
            .O(N__49108),
            .I(N__49088));
    LocalMux I__11839 (
            .O(N__49105),
            .I(N__49088));
    InMux I__11838 (
            .O(N__49104),
            .I(N__49077));
    InMux I__11837 (
            .O(N__49103),
            .I(N__49077));
    InMux I__11836 (
            .O(N__49102),
            .I(N__49077));
    InMux I__11835 (
            .O(N__49101),
            .I(N__49077));
    InMux I__11834 (
            .O(N__49100),
            .I(N__49077));
    InMux I__11833 (
            .O(N__49099),
            .I(N__49072));
    InMux I__11832 (
            .O(N__49096),
            .I(N__49072));
    InMux I__11831 (
            .O(N__49095),
            .I(N__49069));
    Span4Mux_v I__11830 (
            .O(N__49088),
            .I(N__49066));
    LocalMux I__11829 (
            .O(N__49077),
            .I(N__49063));
    LocalMux I__11828 (
            .O(N__49072),
            .I(N__49058));
    LocalMux I__11827 (
            .O(N__49069),
            .I(N__49058));
    Span4Mux_h I__11826 (
            .O(N__49066),
            .I(N__49053));
    Span4Mux_v I__11825 (
            .O(N__49063),
            .I(N__49053));
    Span4Mux_v I__11824 (
            .O(N__49058),
            .I(N__49050));
    Span4Mux_v I__11823 (
            .O(N__49053),
            .I(N__49047));
    Span4Mux_h I__11822 (
            .O(N__49050),
            .I(N__49044));
    Odrv4 I__11821 (
            .O(N__49047),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__11820 (
            .O(N__49044),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    CascadeMux I__11819 (
            .O(N__49039),
            .I(N__49036));
    InMux I__11818 (
            .O(N__49036),
            .I(N__49026));
    InMux I__11817 (
            .O(N__49035),
            .I(N__49026));
    InMux I__11816 (
            .O(N__49034),
            .I(N__49026));
    InMux I__11815 (
            .O(N__49033),
            .I(N__49023));
    LocalMux I__11814 (
            .O(N__49026),
            .I(N__49018));
    LocalMux I__11813 (
            .O(N__49023),
            .I(N__49018));
    Odrv4 I__11812 (
            .O(N__49018),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    InMux I__11811 (
            .O(N__49015),
            .I(N__49010));
    InMux I__11810 (
            .O(N__49014),
            .I(N__49005));
    InMux I__11809 (
            .O(N__49013),
            .I(N__49005));
    LocalMux I__11808 (
            .O(N__49010),
            .I(N__49002));
    LocalMux I__11807 (
            .O(N__49005),
            .I(N__48999));
    Span4Mux_v I__11806 (
            .O(N__49002),
            .I(N__48996));
    Span4Mux_v I__11805 (
            .O(N__48999),
            .I(N__48993));
    Span4Mux_h I__11804 (
            .O(N__48996),
            .I(N__48990));
    Odrv4 I__11803 (
            .O(N__48993),
            .I(il_min_comp2_D2));
    Odrv4 I__11802 (
            .O(N__48990),
            .I(il_min_comp2_D2));
    InMux I__11801 (
            .O(N__48985),
            .I(N__48982));
    LocalMux I__11800 (
            .O(N__48982),
            .I(N__48979));
    Span4Mux_h I__11799 (
            .O(N__48979),
            .I(N__48976));
    Odrv4 I__11798 (
            .O(N__48976),
            .I(\phase_controller_slave.start_timer_tr_0_sqmuxa ));
    InMux I__11797 (
            .O(N__48973),
            .I(N__48968));
    InMux I__11796 (
            .O(N__48972),
            .I(N__48965));
    InMux I__11795 (
            .O(N__48971),
            .I(N__48962));
    LocalMux I__11794 (
            .O(N__48968),
            .I(N__48959));
    LocalMux I__11793 (
            .O(N__48965),
            .I(\phase_controller_slave.tr_time_passed ));
    LocalMux I__11792 (
            .O(N__48962),
            .I(\phase_controller_slave.tr_time_passed ));
    Odrv4 I__11791 (
            .O(N__48959),
            .I(\phase_controller_slave.tr_time_passed ));
    InMux I__11790 (
            .O(N__48952),
            .I(N__48949));
    LocalMux I__11789 (
            .O(N__48949),
            .I(N__48945));
    InMux I__11788 (
            .O(N__48948),
            .I(N__48942));
    Span4Mux_h I__11787 (
            .O(N__48945),
            .I(N__48939));
    LocalMux I__11786 (
            .O(N__48942),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    Odrv4 I__11785 (
            .O(N__48939),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    InMux I__11784 (
            .O(N__48934),
            .I(N__48928));
    InMux I__11783 (
            .O(N__48933),
            .I(N__48928));
    LocalMux I__11782 (
            .O(N__48928),
            .I(N__48925));
    Odrv4 I__11781 (
            .O(N__48925),
            .I(\phase_controller_slave.N_211 ));
    InMux I__11780 (
            .O(N__48922),
            .I(N__48919));
    LocalMux I__11779 (
            .O(N__48919),
            .I(N__48916));
    Span4Mux_v I__11778 (
            .O(N__48916),
            .I(N__48913));
    Span4Mux_h I__11777 (
            .O(N__48913),
            .I(N__48908));
    InMux I__11776 (
            .O(N__48912),
            .I(N__48905));
    InMux I__11775 (
            .O(N__48911),
            .I(N__48902));
    Odrv4 I__11774 (
            .O(N__48908),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__11773 (
            .O(N__48905),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__11772 (
            .O(N__48902),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__11771 (
            .O(N__48895),
            .I(N__48891));
    InMux I__11770 (
            .O(N__48894),
            .I(N__48888));
    LocalMux I__11769 (
            .O(N__48891),
            .I(N__48885));
    LocalMux I__11768 (
            .O(N__48888),
            .I(N__48882));
    Span4Mux_h I__11767 (
            .O(N__48885),
            .I(N__48879));
    Odrv12 I__11766 (
            .O(N__48882),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    Odrv4 I__11765 (
            .O(N__48879),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    ClkMux I__11764 (
            .O(N__48874),
            .I(N__48349));
    ClkMux I__11763 (
            .O(N__48873),
            .I(N__48349));
    ClkMux I__11762 (
            .O(N__48872),
            .I(N__48349));
    ClkMux I__11761 (
            .O(N__48871),
            .I(N__48349));
    ClkMux I__11760 (
            .O(N__48870),
            .I(N__48349));
    ClkMux I__11759 (
            .O(N__48869),
            .I(N__48349));
    ClkMux I__11758 (
            .O(N__48868),
            .I(N__48349));
    ClkMux I__11757 (
            .O(N__48867),
            .I(N__48349));
    ClkMux I__11756 (
            .O(N__48866),
            .I(N__48349));
    ClkMux I__11755 (
            .O(N__48865),
            .I(N__48349));
    ClkMux I__11754 (
            .O(N__48864),
            .I(N__48349));
    ClkMux I__11753 (
            .O(N__48863),
            .I(N__48349));
    ClkMux I__11752 (
            .O(N__48862),
            .I(N__48349));
    ClkMux I__11751 (
            .O(N__48861),
            .I(N__48349));
    ClkMux I__11750 (
            .O(N__48860),
            .I(N__48349));
    ClkMux I__11749 (
            .O(N__48859),
            .I(N__48349));
    ClkMux I__11748 (
            .O(N__48858),
            .I(N__48349));
    ClkMux I__11747 (
            .O(N__48857),
            .I(N__48349));
    ClkMux I__11746 (
            .O(N__48856),
            .I(N__48349));
    ClkMux I__11745 (
            .O(N__48855),
            .I(N__48349));
    ClkMux I__11744 (
            .O(N__48854),
            .I(N__48349));
    ClkMux I__11743 (
            .O(N__48853),
            .I(N__48349));
    ClkMux I__11742 (
            .O(N__48852),
            .I(N__48349));
    ClkMux I__11741 (
            .O(N__48851),
            .I(N__48349));
    ClkMux I__11740 (
            .O(N__48850),
            .I(N__48349));
    ClkMux I__11739 (
            .O(N__48849),
            .I(N__48349));
    ClkMux I__11738 (
            .O(N__48848),
            .I(N__48349));
    ClkMux I__11737 (
            .O(N__48847),
            .I(N__48349));
    ClkMux I__11736 (
            .O(N__48846),
            .I(N__48349));
    ClkMux I__11735 (
            .O(N__48845),
            .I(N__48349));
    ClkMux I__11734 (
            .O(N__48844),
            .I(N__48349));
    ClkMux I__11733 (
            .O(N__48843),
            .I(N__48349));
    ClkMux I__11732 (
            .O(N__48842),
            .I(N__48349));
    ClkMux I__11731 (
            .O(N__48841),
            .I(N__48349));
    ClkMux I__11730 (
            .O(N__48840),
            .I(N__48349));
    ClkMux I__11729 (
            .O(N__48839),
            .I(N__48349));
    ClkMux I__11728 (
            .O(N__48838),
            .I(N__48349));
    ClkMux I__11727 (
            .O(N__48837),
            .I(N__48349));
    ClkMux I__11726 (
            .O(N__48836),
            .I(N__48349));
    ClkMux I__11725 (
            .O(N__48835),
            .I(N__48349));
    ClkMux I__11724 (
            .O(N__48834),
            .I(N__48349));
    ClkMux I__11723 (
            .O(N__48833),
            .I(N__48349));
    ClkMux I__11722 (
            .O(N__48832),
            .I(N__48349));
    ClkMux I__11721 (
            .O(N__48831),
            .I(N__48349));
    ClkMux I__11720 (
            .O(N__48830),
            .I(N__48349));
    ClkMux I__11719 (
            .O(N__48829),
            .I(N__48349));
    ClkMux I__11718 (
            .O(N__48828),
            .I(N__48349));
    ClkMux I__11717 (
            .O(N__48827),
            .I(N__48349));
    ClkMux I__11716 (
            .O(N__48826),
            .I(N__48349));
    ClkMux I__11715 (
            .O(N__48825),
            .I(N__48349));
    ClkMux I__11714 (
            .O(N__48824),
            .I(N__48349));
    ClkMux I__11713 (
            .O(N__48823),
            .I(N__48349));
    ClkMux I__11712 (
            .O(N__48822),
            .I(N__48349));
    ClkMux I__11711 (
            .O(N__48821),
            .I(N__48349));
    ClkMux I__11710 (
            .O(N__48820),
            .I(N__48349));
    ClkMux I__11709 (
            .O(N__48819),
            .I(N__48349));
    ClkMux I__11708 (
            .O(N__48818),
            .I(N__48349));
    ClkMux I__11707 (
            .O(N__48817),
            .I(N__48349));
    ClkMux I__11706 (
            .O(N__48816),
            .I(N__48349));
    ClkMux I__11705 (
            .O(N__48815),
            .I(N__48349));
    ClkMux I__11704 (
            .O(N__48814),
            .I(N__48349));
    ClkMux I__11703 (
            .O(N__48813),
            .I(N__48349));
    ClkMux I__11702 (
            .O(N__48812),
            .I(N__48349));
    ClkMux I__11701 (
            .O(N__48811),
            .I(N__48349));
    ClkMux I__11700 (
            .O(N__48810),
            .I(N__48349));
    ClkMux I__11699 (
            .O(N__48809),
            .I(N__48349));
    ClkMux I__11698 (
            .O(N__48808),
            .I(N__48349));
    ClkMux I__11697 (
            .O(N__48807),
            .I(N__48349));
    ClkMux I__11696 (
            .O(N__48806),
            .I(N__48349));
    ClkMux I__11695 (
            .O(N__48805),
            .I(N__48349));
    ClkMux I__11694 (
            .O(N__48804),
            .I(N__48349));
    ClkMux I__11693 (
            .O(N__48803),
            .I(N__48349));
    ClkMux I__11692 (
            .O(N__48802),
            .I(N__48349));
    ClkMux I__11691 (
            .O(N__48801),
            .I(N__48349));
    ClkMux I__11690 (
            .O(N__48800),
            .I(N__48349));
    ClkMux I__11689 (
            .O(N__48799),
            .I(N__48349));
    ClkMux I__11688 (
            .O(N__48798),
            .I(N__48349));
    ClkMux I__11687 (
            .O(N__48797),
            .I(N__48349));
    ClkMux I__11686 (
            .O(N__48796),
            .I(N__48349));
    ClkMux I__11685 (
            .O(N__48795),
            .I(N__48349));
    ClkMux I__11684 (
            .O(N__48794),
            .I(N__48349));
    ClkMux I__11683 (
            .O(N__48793),
            .I(N__48349));
    ClkMux I__11682 (
            .O(N__48792),
            .I(N__48349));
    ClkMux I__11681 (
            .O(N__48791),
            .I(N__48349));
    ClkMux I__11680 (
            .O(N__48790),
            .I(N__48349));
    ClkMux I__11679 (
            .O(N__48789),
            .I(N__48349));
    ClkMux I__11678 (
            .O(N__48788),
            .I(N__48349));
    ClkMux I__11677 (
            .O(N__48787),
            .I(N__48349));
    ClkMux I__11676 (
            .O(N__48786),
            .I(N__48349));
    ClkMux I__11675 (
            .O(N__48785),
            .I(N__48349));
    ClkMux I__11674 (
            .O(N__48784),
            .I(N__48349));
    ClkMux I__11673 (
            .O(N__48783),
            .I(N__48349));
    ClkMux I__11672 (
            .O(N__48782),
            .I(N__48349));
    ClkMux I__11671 (
            .O(N__48781),
            .I(N__48349));
    ClkMux I__11670 (
            .O(N__48780),
            .I(N__48349));
    ClkMux I__11669 (
            .O(N__48779),
            .I(N__48349));
    ClkMux I__11668 (
            .O(N__48778),
            .I(N__48349));
    ClkMux I__11667 (
            .O(N__48777),
            .I(N__48349));
    ClkMux I__11666 (
            .O(N__48776),
            .I(N__48349));
    ClkMux I__11665 (
            .O(N__48775),
            .I(N__48349));
    ClkMux I__11664 (
            .O(N__48774),
            .I(N__48349));
    ClkMux I__11663 (
            .O(N__48773),
            .I(N__48349));
    ClkMux I__11662 (
            .O(N__48772),
            .I(N__48349));
    ClkMux I__11661 (
            .O(N__48771),
            .I(N__48349));
    ClkMux I__11660 (
            .O(N__48770),
            .I(N__48349));
    ClkMux I__11659 (
            .O(N__48769),
            .I(N__48349));
    ClkMux I__11658 (
            .O(N__48768),
            .I(N__48349));
    ClkMux I__11657 (
            .O(N__48767),
            .I(N__48349));
    ClkMux I__11656 (
            .O(N__48766),
            .I(N__48349));
    ClkMux I__11655 (
            .O(N__48765),
            .I(N__48349));
    ClkMux I__11654 (
            .O(N__48764),
            .I(N__48349));
    ClkMux I__11653 (
            .O(N__48763),
            .I(N__48349));
    ClkMux I__11652 (
            .O(N__48762),
            .I(N__48349));
    ClkMux I__11651 (
            .O(N__48761),
            .I(N__48349));
    ClkMux I__11650 (
            .O(N__48760),
            .I(N__48349));
    ClkMux I__11649 (
            .O(N__48759),
            .I(N__48349));
    ClkMux I__11648 (
            .O(N__48758),
            .I(N__48349));
    ClkMux I__11647 (
            .O(N__48757),
            .I(N__48349));
    ClkMux I__11646 (
            .O(N__48756),
            .I(N__48349));
    ClkMux I__11645 (
            .O(N__48755),
            .I(N__48349));
    ClkMux I__11644 (
            .O(N__48754),
            .I(N__48349));
    ClkMux I__11643 (
            .O(N__48753),
            .I(N__48349));
    ClkMux I__11642 (
            .O(N__48752),
            .I(N__48349));
    ClkMux I__11641 (
            .O(N__48751),
            .I(N__48349));
    ClkMux I__11640 (
            .O(N__48750),
            .I(N__48349));
    ClkMux I__11639 (
            .O(N__48749),
            .I(N__48349));
    ClkMux I__11638 (
            .O(N__48748),
            .I(N__48349));
    ClkMux I__11637 (
            .O(N__48747),
            .I(N__48349));
    ClkMux I__11636 (
            .O(N__48746),
            .I(N__48349));
    ClkMux I__11635 (
            .O(N__48745),
            .I(N__48349));
    ClkMux I__11634 (
            .O(N__48744),
            .I(N__48349));
    ClkMux I__11633 (
            .O(N__48743),
            .I(N__48349));
    ClkMux I__11632 (
            .O(N__48742),
            .I(N__48349));
    ClkMux I__11631 (
            .O(N__48741),
            .I(N__48349));
    ClkMux I__11630 (
            .O(N__48740),
            .I(N__48349));
    ClkMux I__11629 (
            .O(N__48739),
            .I(N__48349));
    ClkMux I__11628 (
            .O(N__48738),
            .I(N__48349));
    ClkMux I__11627 (
            .O(N__48737),
            .I(N__48349));
    ClkMux I__11626 (
            .O(N__48736),
            .I(N__48349));
    ClkMux I__11625 (
            .O(N__48735),
            .I(N__48349));
    ClkMux I__11624 (
            .O(N__48734),
            .I(N__48349));
    ClkMux I__11623 (
            .O(N__48733),
            .I(N__48349));
    ClkMux I__11622 (
            .O(N__48732),
            .I(N__48349));
    ClkMux I__11621 (
            .O(N__48731),
            .I(N__48349));
    ClkMux I__11620 (
            .O(N__48730),
            .I(N__48349));
    ClkMux I__11619 (
            .O(N__48729),
            .I(N__48349));
    ClkMux I__11618 (
            .O(N__48728),
            .I(N__48349));
    ClkMux I__11617 (
            .O(N__48727),
            .I(N__48349));
    ClkMux I__11616 (
            .O(N__48726),
            .I(N__48349));
    ClkMux I__11615 (
            .O(N__48725),
            .I(N__48349));
    ClkMux I__11614 (
            .O(N__48724),
            .I(N__48349));
    ClkMux I__11613 (
            .O(N__48723),
            .I(N__48349));
    ClkMux I__11612 (
            .O(N__48722),
            .I(N__48349));
    ClkMux I__11611 (
            .O(N__48721),
            .I(N__48349));
    ClkMux I__11610 (
            .O(N__48720),
            .I(N__48349));
    ClkMux I__11609 (
            .O(N__48719),
            .I(N__48349));
    ClkMux I__11608 (
            .O(N__48718),
            .I(N__48349));
    ClkMux I__11607 (
            .O(N__48717),
            .I(N__48349));
    ClkMux I__11606 (
            .O(N__48716),
            .I(N__48349));
    ClkMux I__11605 (
            .O(N__48715),
            .I(N__48349));
    ClkMux I__11604 (
            .O(N__48714),
            .I(N__48349));
    ClkMux I__11603 (
            .O(N__48713),
            .I(N__48349));
    ClkMux I__11602 (
            .O(N__48712),
            .I(N__48349));
    ClkMux I__11601 (
            .O(N__48711),
            .I(N__48349));
    ClkMux I__11600 (
            .O(N__48710),
            .I(N__48349));
    ClkMux I__11599 (
            .O(N__48709),
            .I(N__48349));
    ClkMux I__11598 (
            .O(N__48708),
            .I(N__48349));
    ClkMux I__11597 (
            .O(N__48707),
            .I(N__48349));
    ClkMux I__11596 (
            .O(N__48706),
            .I(N__48349));
    ClkMux I__11595 (
            .O(N__48705),
            .I(N__48349));
    ClkMux I__11594 (
            .O(N__48704),
            .I(N__48349));
    ClkMux I__11593 (
            .O(N__48703),
            .I(N__48349));
    ClkMux I__11592 (
            .O(N__48702),
            .I(N__48349));
    ClkMux I__11591 (
            .O(N__48701),
            .I(N__48349));
    ClkMux I__11590 (
            .O(N__48700),
            .I(N__48349));
    GlobalMux I__11589 (
            .O(N__48349),
            .I(clk_100mhz_0));
    CEMux I__11588 (
            .O(N__48346),
            .I(N__48340));
    CEMux I__11587 (
            .O(N__48345),
            .I(N__48335));
    CEMux I__11586 (
            .O(N__48344),
            .I(N__48332));
    CEMux I__11585 (
            .O(N__48343),
            .I(N__48329));
    LocalMux I__11584 (
            .O(N__48340),
            .I(N__48326));
    CEMux I__11583 (
            .O(N__48339),
            .I(N__48323));
    CEMux I__11582 (
            .O(N__48338),
            .I(N__48320));
    LocalMux I__11581 (
            .O(N__48335),
            .I(N__48317));
    LocalMux I__11580 (
            .O(N__48332),
            .I(N__48312));
    LocalMux I__11579 (
            .O(N__48329),
            .I(N__48312));
    Span4Mux_h I__11578 (
            .O(N__48326),
            .I(N__48309));
    LocalMux I__11577 (
            .O(N__48323),
            .I(N__48306));
    LocalMux I__11576 (
            .O(N__48320),
            .I(N__48303));
    Span12Mux_s8_h I__11575 (
            .O(N__48317),
            .I(N__48300));
    Span4Mux_v I__11574 (
            .O(N__48312),
            .I(N__48297));
    Span4Mux_v I__11573 (
            .O(N__48309),
            .I(N__48292));
    Span4Mux_v I__11572 (
            .O(N__48306),
            .I(N__48292));
    Span4Mux_h I__11571 (
            .O(N__48303),
            .I(N__48289));
    Odrv12 I__11570 (
            .O(N__48300),
            .I(\delay_measurement_inst.delay_tr_timer.N_338_i ));
    Odrv4 I__11569 (
            .O(N__48297),
            .I(\delay_measurement_inst.delay_tr_timer.N_338_i ));
    Odrv4 I__11568 (
            .O(N__48292),
            .I(\delay_measurement_inst.delay_tr_timer.N_338_i ));
    Odrv4 I__11567 (
            .O(N__48289),
            .I(\delay_measurement_inst.delay_tr_timer.N_338_i ));
    CascadeMux I__11566 (
            .O(N__48280),
            .I(N__48272));
    InMux I__11565 (
            .O(N__48279),
            .I(N__48269));
    InMux I__11564 (
            .O(N__48278),
            .I(N__48266));
    InMux I__11563 (
            .O(N__48277),
            .I(N__48263));
    InMux I__11562 (
            .O(N__48276),
            .I(N__48260));
    InMux I__11561 (
            .O(N__48275),
            .I(N__48257));
    InMux I__11560 (
            .O(N__48272),
            .I(N__48254));
    LocalMux I__11559 (
            .O(N__48269),
            .I(N__48251));
    LocalMux I__11558 (
            .O(N__48266),
            .I(N__48248));
    LocalMux I__11557 (
            .O(N__48263),
            .I(N__48245));
    LocalMux I__11556 (
            .O(N__48260),
            .I(N__48242));
    LocalMux I__11555 (
            .O(N__48257),
            .I(N__48167));
    LocalMux I__11554 (
            .O(N__48254),
            .I(N__48114));
    Glb2LocalMux I__11553 (
            .O(N__48251),
            .I(N__47779));
    Glb2LocalMux I__11552 (
            .O(N__48248),
            .I(N__47779));
    Glb2LocalMux I__11551 (
            .O(N__48245),
            .I(N__47779));
    Glb2LocalMux I__11550 (
            .O(N__48242),
            .I(N__47779));
    SRMux I__11549 (
            .O(N__48241),
            .I(N__47779));
    SRMux I__11548 (
            .O(N__48240),
            .I(N__47779));
    SRMux I__11547 (
            .O(N__48239),
            .I(N__47779));
    SRMux I__11546 (
            .O(N__48238),
            .I(N__47779));
    SRMux I__11545 (
            .O(N__48237),
            .I(N__47779));
    SRMux I__11544 (
            .O(N__48236),
            .I(N__47779));
    SRMux I__11543 (
            .O(N__48235),
            .I(N__47779));
    SRMux I__11542 (
            .O(N__48234),
            .I(N__47779));
    SRMux I__11541 (
            .O(N__48233),
            .I(N__47779));
    SRMux I__11540 (
            .O(N__48232),
            .I(N__47779));
    SRMux I__11539 (
            .O(N__48231),
            .I(N__47779));
    SRMux I__11538 (
            .O(N__48230),
            .I(N__47779));
    SRMux I__11537 (
            .O(N__48229),
            .I(N__47779));
    SRMux I__11536 (
            .O(N__48228),
            .I(N__47779));
    SRMux I__11535 (
            .O(N__48227),
            .I(N__47779));
    SRMux I__11534 (
            .O(N__48226),
            .I(N__47779));
    SRMux I__11533 (
            .O(N__48225),
            .I(N__47779));
    SRMux I__11532 (
            .O(N__48224),
            .I(N__47779));
    SRMux I__11531 (
            .O(N__48223),
            .I(N__47779));
    SRMux I__11530 (
            .O(N__48222),
            .I(N__47779));
    SRMux I__11529 (
            .O(N__48221),
            .I(N__47779));
    SRMux I__11528 (
            .O(N__48220),
            .I(N__47779));
    SRMux I__11527 (
            .O(N__48219),
            .I(N__47779));
    SRMux I__11526 (
            .O(N__48218),
            .I(N__47779));
    SRMux I__11525 (
            .O(N__48217),
            .I(N__47779));
    SRMux I__11524 (
            .O(N__48216),
            .I(N__47779));
    SRMux I__11523 (
            .O(N__48215),
            .I(N__47779));
    SRMux I__11522 (
            .O(N__48214),
            .I(N__47779));
    SRMux I__11521 (
            .O(N__48213),
            .I(N__47779));
    SRMux I__11520 (
            .O(N__48212),
            .I(N__47779));
    SRMux I__11519 (
            .O(N__48211),
            .I(N__47779));
    SRMux I__11518 (
            .O(N__48210),
            .I(N__47779));
    SRMux I__11517 (
            .O(N__48209),
            .I(N__47779));
    SRMux I__11516 (
            .O(N__48208),
            .I(N__47779));
    SRMux I__11515 (
            .O(N__48207),
            .I(N__47779));
    SRMux I__11514 (
            .O(N__48206),
            .I(N__47779));
    SRMux I__11513 (
            .O(N__48205),
            .I(N__47779));
    SRMux I__11512 (
            .O(N__48204),
            .I(N__47779));
    SRMux I__11511 (
            .O(N__48203),
            .I(N__47779));
    SRMux I__11510 (
            .O(N__48202),
            .I(N__47779));
    SRMux I__11509 (
            .O(N__48201),
            .I(N__47779));
    SRMux I__11508 (
            .O(N__48200),
            .I(N__47779));
    SRMux I__11507 (
            .O(N__48199),
            .I(N__47779));
    SRMux I__11506 (
            .O(N__48198),
            .I(N__47779));
    SRMux I__11505 (
            .O(N__48197),
            .I(N__47779));
    SRMux I__11504 (
            .O(N__48196),
            .I(N__47779));
    SRMux I__11503 (
            .O(N__48195),
            .I(N__47779));
    SRMux I__11502 (
            .O(N__48194),
            .I(N__47779));
    SRMux I__11501 (
            .O(N__48193),
            .I(N__47779));
    SRMux I__11500 (
            .O(N__48192),
            .I(N__47779));
    SRMux I__11499 (
            .O(N__48191),
            .I(N__47779));
    SRMux I__11498 (
            .O(N__48190),
            .I(N__47779));
    SRMux I__11497 (
            .O(N__48189),
            .I(N__47779));
    SRMux I__11496 (
            .O(N__48188),
            .I(N__47779));
    SRMux I__11495 (
            .O(N__48187),
            .I(N__47779));
    SRMux I__11494 (
            .O(N__48186),
            .I(N__47779));
    SRMux I__11493 (
            .O(N__48185),
            .I(N__47779));
    SRMux I__11492 (
            .O(N__48184),
            .I(N__47779));
    SRMux I__11491 (
            .O(N__48183),
            .I(N__47779));
    SRMux I__11490 (
            .O(N__48182),
            .I(N__47779));
    SRMux I__11489 (
            .O(N__48181),
            .I(N__47779));
    SRMux I__11488 (
            .O(N__48180),
            .I(N__47779));
    SRMux I__11487 (
            .O(N__48179),
            .I(N__47779));
    SRMux I__11486 (
            .O(N__48178),
            .I(N__47779));
    SRMux I__11485 (
            .O(N__48177),
            .I(N__47779));
    SRMux I__11484 (
            .O(N__48176),
            .I(N__47779));
    SRMux I__11483 (
            .O(N__48175),
            .I(N__47779));
    SRMux I__11482 (
            .O(N__48174),
            .I(N__47779));
    SRMux I__11481 (
            .O(N__48173),
            .I(N__47779));
    SRMux I__11480 (
            .O(N__48172),
            .I(N__47779));
    SRMux I__11479 (
            .O(N__48171),
            .I(N__47779));
    SRMux I__11478 (
            .O(N__48170),
            .I(N__47779));
    Glb2LocalMux I__11477 (
            .O(N__48167),
            .I(N__47779));
    SRMux I__11476 (
            .O(N__48166),
            .I(N__47779));
    SRMux I__11475 (
            .O(N__48165),
            .I(N__47779));
    SRMux I__11474 (
            .O(N__48164),
            .I(N__47779));
    SRMux I__11473 (
            .O(N__48163),
            .I(N__47779));
    SRMux I__11472 (
            .O(N__48162),
            .I(N__47779));
    SRMux I__11471 (
            .O(N__48161),
            .I(N__47779));
    SRMux I__11470 (
            .O(N__48160),
            .I(N__47779));
    SRMux I__11469 (
            .O(N__48159),
            .I(N__47779));
    SRMux I__11468 (
            .O(N__48158),
            .I(N__47779));
    SRMux I__11467 (
            .O(N__48157),
            .I(N__47779));
    SRMux I__11466 (
            .O(N__48156),
            .I(N__47779));
    SRMux I__11465 (
            .O(N__48155),
            .I(N__47779));
    SRMux I__11464 (
            .O(N__48154),
            .I(N__47779));
    SRMux I__11463 (
            .O(N__48153),
            .I(N__47779));
    SRMux I__11462 (
            .O(N__48152),
            .I(N__47779));
    SRMux I__11461 (
            .O(N__48151),
            .I(N__47779));
    SRMux I__11460 (
            .O(N__48150),
            .I(N__47779));
    SRMux I__11459 (
            .O(N__48149),
            .I(N__47779));
    SRMux I__11458 (
            .O(N__48148),
            .I(N__47779));
    SRMux I__11457 (
            .O(N__48147),
            .I(N__47779));
    SRMux I__11456 (
            .O(N__48146),
            .I(N__47779));
    SRMux I__11455 (
            .O(N__48145),
            .I(N__47779));
    SRMux I__11454 (
            .O(N__48144),
            .I(N__47779));
    SRMux I__11453 (
            .O(N__48143),
            .I(N__47779));
    SRMux I__11452 (
            .O(N__48142),
            .I(N__47779));
    SRMux I__11451 (
            .O(N__48141),
            .I(N__47779));
    SRMux I__11450 (
            .O(N__48140),
            .I(N__47779));
    SRMux I__11449 (
            .O(N__48139),
            .I(N__47779));
    SRMux I__11448 (
            .O(N__48138),
            .I(N__47779));
    SRMux I__11447 (
            .O(N__48137),
            .I(N__47779));
    SRMux I__11446 (
            .O(N__48136),
            .I(N__47779));
    SRMux I__11445 (
            .O(N__48135),
            .I(N__47779));
    SRMux I__11444 (
            .O(N__48134),
            .I(N__47779));
    SRMux I__11443 (
            .O(N__48133),
            .I(N__47779));
    SRMux I__11442 (
            .O(N__48132),
            .I(N__47779));
    SRMux I__11441 (
            .O(N__48131),
            .I(N__47779));
    SRMux I__11440 (
            .O(N__48130),
            .I(N__47779));
    SRMux I__11439 (
            .O(N__48129),
            .I(N__47779));
    SRMux I__11438 (
            .O(N__48128),
            .I(N__47779));
    SRMux I__11437 (
            .O(N__48127),
            .I(N__47779));
    SRMux I__11436 (
            .O(N__48126),
            .I(N__47779));
    SRMux I__11435 (
            .O(N__48125),
            .I(N__47779));
    SRMux I__11434 (
            .O(N__48124),
            .I(N__47779));
    SRMux I__11433 (
            .O(N__48123),
            .I(N__47779));
    SRMux I__11432 (
            .O(N__48122),
            .I(N__47779));
    SRMux I__11431 (
            .O(N__48121),
            .I(N__47779));
    SRMux I__11430 (
            .O(N__48120),
            .I(N__47779));
    SRMux I__11429 (
            .O(N__48119),
            .I(N__47779));
    SRMux I__11428 (
            .O(N__48118),
            .I(N__47779));
    SRMux I__11427 (
            .O(N__48117),
            .I(N__47779));
    Glb2LocalMux I__11426 (
            .O(N__48114),
            .I(N__47779));
    SRMux I__11425 (
            .O(N__48113),
            .I(N__47779));
    SRMux I__11424 (
            .O(N__48112),
            .I(N__47779));
    SRMux I__11423 (
            .O(N__48111),
            .I(N__47779));
    SRMux I__11422 (
            .O(N__48110),
            .I(N__47779));
    SRMux I__11421 (
            .O(N__48109),
            .I(N__47779));
    SRMux I__11420 (
            .O(N__48108),
            .I(N__47779));
    SRMux I__11419 (
            .O(N__48107),
            .I(N__47779));
    SRMux I__11418 (
            .O(N__48106),
            .I(N__47779));
    SRMux I__11417 (
            .O(N__48105),
            .I(N__47779));
    SRMux I__11416 (
            .O(N__48104),
            .I(N__47779));
    SRMux I__11415 (
            .O(N__48103),
            .I(N__47779));
    SRMux I__11414 (
            .O(N__48102),
            .I(N__47779));
    SRMux I__11413 (
            .O(N__48101),
            .I(N__47779));
    SRMux I__11412 (
            .O(N__48100),
            .I(N__47779));
    SRMux I__11411 (
            .O(N__48099),
            .I(N__47779));
    SRMux I__11410 (
            .O(N__48098),
            .I(N__47779));
    SRMux I__11409 (
            .O(N__48097),
            .I(N__47779));
    SRMux I__11408 (
            .O(N__48096),
            .I(N__47779));
    SRMux I__11407 (
            .O(N__48095),
            .I(N__47779));
    SRMux I__11406 (
            .O(N__48094),
            .I(N__47779));
    SRMux I__11405 (
            .O(N__48093),
            .I(N__47779));
    SRMux I__11404 (
            .O(N__48092),
            .I(N__47779));
    SRMux I__11403 (
            .O(N__48091),
            .I(N__47779));
    SRMux I__11402 (
            .O(N__48090),
            .I(N__47779));
    SRMux I__11401 (
            .O(N__48089),
            .I(N__47779));
    SRMux I__11400 (
            .O(N__48088),
            .I(N__47779));
    GlobalMux I__11399 (
            .O(N__47779),
            .I(N__47776));
    gio2CtrlBuf I__11398 (
            .O(N__47776),
            .I(red_c_g));
    CascadeMux I__11397 (
            .O(N__47773),
            .I(N__47768));
    CascadeMux I__11396 (
            .O(N__47772),
            .I(N__47765));
    InMux I__11395 (
            .O(N__47771),
            .I(N__47762));
    InMux I__11394 (
            .O(N__47768),
            .I(N__47757));
    InMux I__11393 (
            .O(N__47765),
            .I(N__47757));
    LocalMux I__11392 (
            .O(N__47762),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__11391 (
            .O(N__47757),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__11390 (
            .O(N__47752),
            .I(N__47749));
    LocalMux I__11389 (
            .O(N__47749),
            .I(N__47746));
    Span4Mux_v I__11388 (
            .O(N__47746),
            .I(N__47743));
    Odrv4 I__11387 (
            .O(N__47743),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__11386 (
            .O(N__47740),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__11385 (
            .O(N__47737),
            .I(N__47732));
    CascadeMux I__11384 (
            .O(N__47736),
            .I(N__47729));
    InMux I__11383 (
            .O(N__47735),
            .I(N__47726));
    InMux I__11382 (
            .O(N__47732),
            .I(N__47721));
    InMux I__11381 (
            .O(N__47729),
            .I(N__47721));
    LocalMux I__11380 (
            .O(N__47726),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__11379 (
            .O(N__47721),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__11378 (
            .O(N__47716),
            .I(N__47713));
    LocalMux I__11377 (
            .O(N__47713),
            .I(N__47710));
    Span4Mux_v I__11376 (
            .O(N__47710),
            .I(N__47707));
    Odrv4 I__11375 (
            .O(N__47707),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__11374 (
            .O(N__47704),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__11373 (
            .O(N__47701),
            .I(N__47696));
    InMux I__11372 (
            .O(N__47700),
            .I(N__47691));
    InMux I__11371 (
            .O(N__47699),
            .I(N__47691));
    LocalMux I__11370 (
            .O(N__47696),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__11369 (
            .O(N__47691),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__11368 (
            .O(N__47686),
            .I(N__47683));
    LocalMux I__11367 (
            .O(N__47683),
            .I(N__47680));
    Span4Mux_h I__11366 (
            .O(N__47680),
            .I(N__47677));
    Odrv4 I__11365 (
            .O(N__47677),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__11364 (
            .O(N__47674),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__11363 (
            .O(N__47671),
            .I(N__47666));
    InMux I__11362 (
            .O(N__47670),
            .I(N__47661));
    InMux I__11361 (
            .O(N__47669),
            .I(N__47661));
    LocalMux I__11360 (
            .O(N__47666),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__11359 (
            .O(N__47661),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    CascadeMux I__11358 (
            .O(N__47656),
            .I(N__47653));
    InMux I__11357 (
            .O(N__47653),
            .I(N__47650));
    LocalMux I__11356 (
            .O(N__47650),
            .I(N__47647));
    Span4Mux_h I__11355 (
            .O(N__47647),
            .I(N__47644));
    Odrv4 I__11354 (
            .O(N__47644),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__11353 (
            .O(N__47641),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__11352 (
            .O(N__47638),
            .I(N__47633));
    CascadeMux I__11351 (
            .O(N__47637),
            .I(N__47630));
    InMux I__11350 (
            .O(N__47636),
            .I(N__47627));
    InMux I__11349 (
            .O(N__47633),
            .I(N__47622));
    InMux I__11348 (
            .O(N__47630),
            .I(N__47622));
    LocalMux I__11347 (
            .O(N__47627),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__11346 (
            .O(N__47622),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__11345 (
            .O(N__47617),
            .I(N__47614));
    LocalMux I__11344 (
            .O(N__47614),
            .I(N__47611));
    Span4Mux_h I__11343 (
            .O(N__47611),
            .I(N__47608));
    Odrv4 I__11342 (
            .O(N__47608),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__11341 (
            .O(N__47605),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__11340 (
            .O(N__47602),
            .I(N__47597));
    CascadeMux I__11339 (
            .O(N__47601),
            .I(N__47594));
    InMux I__11338 (
            .O(N__47600),
            .I(N__47591));
    InMux I__11337 (
            .O(N__47597),
            .I(N__47586));
    InMux I__11336 (
            .O(N__47594),
            .I(N__47586));
    LocalMux I__11335 (
            .O(N__47591),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__11334 (
            .O(N__47586),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__11333 (
            .O(N__47581),
            .I(N__47578));
    LocalMux I__11332 (
            .O(N__47578),
            .I(N__47575));
    Span4Mux_h I__11331 (
            .O(N__47575),
            .I(N__47572));
    Odrv4 I__11330 (
            .O(N__47572),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__11329 (
            .O(N__47569),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__11328 (
            .O(N__47566),
            .I(N__47561));
    InMux I__11327 (
            .O(N__47565),
            .I(N__47558));
    InMux I__11326 (
            .O(N__47564),
            .I(N__47555));
    LocalMux I__11325 (
            .O(N__47561),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__11324 (
            .O(N__47558),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__11323 (
            .O(N__47555),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__11322 (
            .O(N__47548),
            .I(N__47545));
    LocalMux I__11321 (
            .O(N__47545),
            .I(N__47542));
    Odrv4 I__11320 (
            .O(N__47542),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__11319 (
            .O(N__47539),
            .I(bfn_18_26_0_));
    InMux I__11318 (
            .O(N__47536),
            .I(N__47531));
    InMux I__11317 (
            .O(N__47535),
            .I(N__47528));
    InMux I__11316 (
            .O(N__47534),
            .I(N__47525));
    LocalMux I__11315 (
            .O(N__47531),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__11314 (
            .O(N__47528),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__11313 (
            .O(N__47525),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    CascadeMux I__11312 (
            .O(N__47518),
            .I(N__47515));
    InMux I__11311 (
            .O(N__47515),
            .I(N__47512));
    LocalMux I__11310 (
            .O(N__47512),
            .I(N__47509));
    Odrv4 I__11309 (
            .O(N__47509),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__11308 (
            .O(N__47506),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    CascadeMux I__11307 (
            .O(N__47503),
            .I(N__47498));
    CascadeMux I__11306 (
            .O(N__47502),
            .I(N__47495));
    InMux I__11305 (
            .O(N__47501),
            .I(N__47492));
    InMux I__11304 (
            .O(N__47498),
            .I(N__47487));
    InMux I__11303 (
            .O(N__47495),
            .I(N__47487));
    LocalMux I__11302 (
            .O(N__47492),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__11301 (
            .O(N__47487),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__11300 (
            .O(N__47482),
            .I(N__47478));
    CascadeMux I__11299 (
            .O(N__47481),
            .I(N__47475));
    LocalMux I__11298 (
            .O(N__47478),
            .I(N__47472));
    InMux I__11297 (
            .O(N__47475),
            .I(N__47469));
    Span4Mux_h I__11296 (
            .O(N__47472),
            .I(N__47466));
    LocalMux I__11295 (
            .O(N__47469),
            .I(N__47463));
    Span4Mux_v I__11294 (
            .O(N__47466),
            .I(N__47460));
    Span4Mux_h I__11293 (
            .O(N__47463),
            .I(N__47457));
    Odrv4 I__11292 (
            .O(N__47460),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    Odrv4 I__11291 (
            .O(N__47457),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    InMux I__11290 (
            .O(N__47452),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__11289 (
            .O(N__47449),
            .I(N__47444));
    CascadeMux I__11288 (
            .O(N__47448),
            .I(N__47441));
    InMux I__11287 (
            .O(N__47447),
            .I(N__47438));
    InMux I__11286 (
            .O(N__47444),
            .I(N__47433));
    InMux I__11285 (
            .O(N__47441),
            .I(N__47433));
    LocalMux I__11284 (
            .O(N__47438),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__11283 (
            .O(N__47433),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__11282 (
            .O(N__47428),
            .I(N__47422));
    InMux I__11281 (
            .O(N__47427),
            .I(N__47419));
    InMux I__11280 (
            .O(N__47426),
            .I(N__47413));
    InMux I__11279 (
            .O(N__47425),
            .I(N__47413));
    LocalMux I__11278 (
            .O(N__47422),
            .I(N__47410));
    LocalMux I__11277 (
            .O(N__47419),
            .I(N__47407));
    InMux I__11276 (
            .O(N__47418),
            .I(N__47404));
    LocalMux I__11275 (
            .O(N__47413),
            .I(N__47399));
    Span4Mux_h I__11274 (
            .O(N__47410),
            .I(N__47399));
    Span4Mux_h I__11273 (
            .O(N__47407),
            .I(N__47394));
    LocalMux I__11272 (
            .O(N__47404),
            .I(N__47394));
    Span4Mux_v I__11271 (
            .O(N__47399),
            .I(N__47391));
    Span4Mux_h I__11270 (
            .O(N__47394),
            .I(N__47388));
    Odrv4 I__11269 (
            .O(N__47391),
            .I(\delay_measurement_inst.elapsed_time_tr_14 ));
    Odrv4 I__11268 (
            .O(N__47388),
            .I(\delay_measurement_inst.elapsed_time_tr_14 ));
    InMux I__11267 (
            .O(N__47383),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__11266 (
            .O(N__47380),
            .I(N__47375));
    InMux I__11265 (
            .O(N__47379),
            .I(N__47370));
    InMux I__11264 (
            .O(N__47378),
            .I(N__47370));
    LocalMux I__11263 (
            .O(N__47375),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__11262 (
            .O(N__47370),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__11261 (
            .O(N__47365),
            .I(N__47358));
    CascadeMux I__11260 (
            .O(N__47364),
            .I(N__47355));
    CascadeMux I__11259 (
            .O(N__47363),
            .I(N__47351));
    InMux I__11258 (
            .O(N__47362),
            .I(N__47348));
    InMux I__11257 (
            .O(N__47361),
            .I(N__47345));
    LocalMux I__11256 (
            .O(N__47358),
            .I(N__47342));
    InMux I__11255 (
            .O(N__47355),
            .I(N__47339));
    InMux I__11254 (
            .O(N__47354),
            .I(N__47336));
    InMux I__11253 (
            .O(N__47351),
            .I(N__47333));
    LocalMux I__11252 (
            .O(N__47348),
            .I(N__47328));
    LocalMux I__11251 (
            .O(N__47345),
            .I(N__47328));
    Span4Mux_h I__11250 (
            .O(N__47342),
            .I(N__47319));
    LocalMux I__11249 (
            .O(N__47339),
            .I(N__47319));
    LocalMux I__11248 (
            .O(N__47336),
            .I(N__47319));
    LocalMux I__11247 (
            .O(N__47333),
            .I(N__47319));
    Span4Mux_v I__11246 (
            .O(N__47328),
            .I(N__47314));
    Span4Mux_h I__11245 (
            .O(N__47319),
            .I(N__47314));
    Odrv4 I__11244 (
            .O(N__47314),
            .I(\delay_measurement_inst.elapsed_time_tr_15 ));
    InMux I__11243 (
            .O(N__47311),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__11242 (
            .O(N__47308),
            .I(N__47303));
    InMux I__11241 (
            .O(N__47307),
            .I(N__47298));
    InMux I__11240 (
            .O(N__47306),
            .I(N__47298));
    LocalMux I__11239 (
            .O(N__47303),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__11238 (
            .O(N__47298),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__11237 (
            .O(N__47293),
            .I(N__47290));
    LocalMux I__11236 (
            .O(N__47290),
            .I(N__47286));
    InMux I__11235 (
            .O(N__47289),
            .I(N__47283));
    Span4Mux_v I__11234 (
            .O(N__47286),
            .I(N__47279));
    LocalMux I__11233 (
            .O(N__47283),
            .I(N__47276));
    InMux I__11232 (
            .O(N__47282),
            .I(N__47273));
    Span4Mux_v I__11231 (
            .O(N__47279),
            .I(N__47268));
    Span4Mux_v I__11230 (
            .O(N__47276),
            .I(N__47268));
    LocalMux I__11229 (
            .O(N__47273),
            .I(N__47265));
    Span4Mux_h I__11228 (
            .O(N__47268),
            .I(N__47262));
    Odrv12 I__11227 (
            .O(N__47265),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    Odrv4 I__11226 (
            .O(N__47262),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    InMux I__11225 (
            .O(N__47257),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__11224 (
            .O(N__47254),
            .I(N__47249));
    CascadeMux I__11223 (
            .O(N__47253),
            .I(N__47246));
    InMux I__11222 (
            .O(N__47252),
            .I(N__47243));
    InMux I__11221 (
            .O(N__47249),
            .I(N__47238));
    InMux I__11220 (
            .O(N__47246),
            .I(N__47238));
    LocalMux I__11219 (
            .O(N__47243),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__11218 (
            .O(N__47238),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__11217 (
            .O(N__47233),
            .I(N__47229));
    InMux I__11216 (
            .O(N__47232),
            .I(N__47225));
    LocalMux I__11215 (
            .O(N__47229),
            .I(N__47222));
    InMux I__11214 (
            .O(N__47228),
            .I(N__47219));
    LocalMux I__11213 (
            .O(N__47225),
            .I(N__47216));
    Span12Mux_h I__11212 (
            .O(N__47222),
            .I(N__47211));
    LocalMux I__11211 (
            .O(N__47219),
            .I(N__47211));
    Span4Mux_h I__11210 (
            .O(N__47216),
            .I(N__47208));
    Odrv12 I__11209 (
            .O(N__47211),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    Odrv4 I__11208 (
            .O(N__47208),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    InMux I__11207 (
            .O(N__47203),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__11206 (
            .O(N__47200),
            .I(N__47195));
    CascadeMux I__11205 (
            .O(N__47199),
            .I(N__47192));
    InMux I__11204 (
            .O(N__47198),
            .I(N__47189));
    InMux I__11203 (
            .O(N__47195),
            .I(N__47184));
    InMux I__11202 (
            .O(N__47192),
            .I(N__47184));
    LocalMux I__11201 (
            .O(N__47189),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__11200 (
            .O(N__47184),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__11199 (
            .O(N__47179),
            .I(N__47176));
    LocalMux I__11198 (
            .O(N__47176),
            .I(N__47173));
    Span4Mux_h I__11197 (
            .O(N__47173),
            .I(N__47169));
    InMux I__11196 (
            .O(N__47172),
            .I(N__47165));
    Span4Mux_h I__11195 (
            .O(N__47169),
            .I(N__47162));
    InMux I__11194 (
            .O(N__47168),
            .I(N__47159));
    LocalMux I__11193 (
            .O(N__47165),
            .I(N__47156));
    Sp12to4 I__11192 (
            .O(N__47162),
            .I(N__47151));
    LocalMux I__11191 (
            .O(N__47159),
            .I(N__47151));
    Span4Mux_h I__11190 (
            .O(N__47156),
            .I(N__47148));
    Odrv12 I__11189 (
            .O(N__47151),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    Odrv4 I__11188 (
            .O(N__47148),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    InMux I__11187 (
            .O(N__47143),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__11186 (
            .O(N__47140),
            .I(N__47135));
    InMux I__11185 (
            .O(N__47139),
            .I(N__47132));
    InMux I__11184 (
            .O(N__47138),
            .I(N__47129));
    LocalMux I__11183 (
            .O(N__47135),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__11182 (
            .O(N__47132),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__11181 (
            .O(N__47129),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__11180 (
            .O(N__47122),
            .I(N__47119));
    LocalMux I__11179 (
            .O(N__47119),
            .I(N__47114));
    CascadeMux I__11178 (
            .O(N__47118),
            .I(N__47111));
    CascadeMux I__11177 (
            .O(N__47117),
            .I(N__47108));
    Span4Mux_h I__11176 (
            .O(N__47114),
            .I(N__47105));
    InMux I__11175 (
            .O(N__47111),
            .I(N__47102));
    InMux I__11174 (
            .O(N__47108),
            .I(N__47099));
    Span4Mux_v I__11173 (
            .O(N__47105),
            .I(N__47096));
    LocalMux I__11172 (
            .O(N__47102),
            .I(N__47093));
    LocalMux I__11171 (
            .O(N__47099),
            .I(N__47090));
    Span4Mux_h I__11170 (
            .O(N__47096),
            .I(N__47087));
    Span4Mux_v I__11169 (
            .O(N__47093),
            .I(N__47082));
    Span4Mux_h I__11168 (
            .O(N__47090),
            .I(N__47082));
    Odrv4 I__11167 (
            .O(N__47087),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    Odrv4 I__11166 (
            .O(N__47082),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    InMux I__11165 (
            .O(N__47077),
            .I(bfn_18_25_0_));
    InMux I__11164 (
            .O(N__47074),
            .I(N__47069));
    InMux I__11163 (
            .O(N__47073),
            .I(N__47066));
    InMux I__11162 (
            .O(N__47072),
            .I(N__47063));
    LocalMux I__11161 (
            .O(N__47069),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__11160 (
            .O(N__47066),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__11159 (
            .O(N__47063),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__11158 (
            .O(N__47056),
            .I(N__47053));
    LocalMux I__11157 (
            .O(N__47053),
            .I(N__47050));
    Span4Mux_h I__11156 (
            .O(N__47050),
            .I(N__47047));
    Odrv4 I__11155 (
            .O(N__47047),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__11154 (
            .O(N__47044),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__11153 (
            .O(N__47041),
            .I(N__47036));
    CascadeMux I__11152 (
            .O(N__47040),
            .I(N__47033));
    InMux I__11151 (
            .O(N__47039),
            .I(N__47030));
    InMux I__11150 (
            .O(N__47036),
            .I(N__47025));
    InMux I__11149 (
            .O(N__47033),
            .I(N__47025));
    LocalMux I__11148 (
            .O(N__47030),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__11147 (
            .O(N__47025),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__11146 (
            .O(N__47020),
            .I(N__47015));
    InMux I__11145 (
            .O(N__47019),
            .I(N__47012));
    InMux I__11144 (
            .O(N__47018),
            .I(N__47009));
    LocalMux I__11143 (
            .O(N__47015),
            .I(N__47002));
    LocalMux I__11142 (
            .O(N__47012),
            .I(N__47002));
    LocalMux I__11141 (
            .O(N__47009),
            .I(N__47002));
    Span4Mux_h I__11140 (
            .O(N__47002),
            .I(N__46999));
    Odrv4 I__11139 (
            .O(N__46999),
            .I(\delay_measurement_inst.elapsed_time_tr_6 ));
    InMux I__11138 (
            .O(N__46996),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__11137 (
            .O(N__46993),
            .I(N__46988));
    InMux I__11136 (
            .O(N__46992),
            .I(N__46983));
    InMux I__11135 (
            .O(N__46991),
            .I(N__46983));
    LocalMux I__11134 (
            .O(N__46988),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__11133 (
            .O(N__46983),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__11132 (
            .O(N__46978),
            .I(N__46975));
    LocalMux I__11131 (
            .O(N__46975),
            .I(N__46972));
    Span4Mux_v I__11130 (
            .O(N__46972),
            .I(N__46967));
    InMux I__11129 (
            .O(N__46971),
            .I(N__46964));
    InMux I__11128 (
            .O(N__46970),
            .I(N__46961));
    Span4Mux_v I__11127 (
            .O(N__46967),
            .I(N__46958));
    LocalMux I__11126 (
            .O(N__46964),
            .I(N__46953));
    LocalMux I__11125 (
            .O(N__46961),
            .I(N__46953));
    Span4Mux_h I__11124 (
            .O(N__46958),
            .I(N__46950));
    Span4Mux_h I__11123 (
            .O(N__46953),
            .I(N__46947));
    Odrv4 I__11122 (
            .O(N__46950),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    Odrv4 I__11121 (
            .O(N__46947),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    InMux I__11120 (
            .O(N__46942),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__11119 (
            .O(N__46939),
            .I(N__46934));
    InMux I__11118 (
            .O(N__46938),
            .I(N__46929));
    InMux I__11117 (
            .O(N__46937),
            .I(N__46929));
    LocalMux I__11116 (
            .O(N__46934),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__11115 (
            .O(N__46929),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__11114 (
            .O(N__46924),
            .I(N__46921));
    LocalMux I__11113 (
            .O(N__46921),
            .I(N__46918));
    Span4Mux_h I__11112 (
            .O(N__46918),
            .I(N__46913));
    InMux I__11111 (
            .O(N__46917),
            .I(N__46910));
    InMux I__11110 (
            .O(N__46916),
            .I(N__46907));
    Span4Mux_h I__11109 (
            .O(N__46913),
            .I(N__46904));
    LocalMux I__11108 (
            .O(N__46910),
            .I(N__46899));
    LocalMux I__11107 (
            .O(N__46907),
            .I(N__46899));
    Span4Mux_v I__11106 (
            .O(N__46904),
            .I(N__46896));
    Span4Mux_h I__11105 (
            .O(N__46899),
            .I(N__46893));
    Odrv4 I__11104 (
            .O(N__46896),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    Odrv4 I__11103 (
            .O(N__46893),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    InMux I__11102 (
            .O(N__46888),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__11101 (
            .O(N__46885),
            .I(N__46880));
    CascadeMux I__11100 (
            .O(N__46884),
            .I(N__46877));
    InMux I__11099 (
            .O(N__46883),
            .I(N__46874));
    InMux I__11098 (
            .O(N__46880),
            .I(N__46869));
    InMux I__11097 (
            .O(N__46877),
            .I(N__46869));
    LocalMux I__11096 (
            .O(N__46874),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__11095 (
            .O(N__46869),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    CascadeMux I__11094 (
            .O(N__46864),
            .I(N__46861));
    InMux I__11093 (
            .O(N__46861),
            .I(N__46857));
    CascadeMux I__11092 (
            .O(N__46860),
            .I(N__46853));
    LocalMux I__11091 (
            .O(N__46857),
            .I(N__46849));
    InMux I__11090 (
            .O(N__46856),
            .I(N__46846));
    InMux I__11089 (
            .O(N__46853),
            .I(N__46843));
    InMux I__11088 (
            .O(N__46852),
            .I(N__46840));
    Span4Mux_h I__11087 (
            .O(N__46849),
            .I(N__46837));
    LocalMux I__11086 (
            .O(N__46846),
            .I(N__46834));
    LocalMux I__11085 (
            .O(N__46843),
            .I(N__46831));
    LocalMux I__11084 (
            .O(N__46840),
            .I(N__46828));
    Span4Mux_v I__11083 (
            .O(N__46837),
            .I(N__46825));
    Span4Mux_v I__11082 (
            .O(N__46834),
            .I(N__46818));
    Span4Mux_v I__11081 (
            .O(N__46831),
            .I(N__46818));
    Span4Mux_h I__11080 (
            .O(N__46828),
            .I(N__46818));
    Odrv4 I__11079 (
            .O(N__46825),
            .I(\delay_measurement_inst.elapsed_time_tr_9 ));
    Odrv4 I__11078 (
            .O(N__46818),
            .I(\delay_measurement_inst.elapsed_time_tr_9 ));
    InMux I__11077 (
            .O(N__46813),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__11076 (
            .O(N__46810),
            .I(N__46805));
    CascadeMux I__11075 (
            .O(N__46809),
            .I(N__46802));
    InMux I__11074 (
            .O(N__46808),
            .I(N__46799));
    InMux I__11073 (
            .O(N__46805),
            .I(N__46794));
    InMux I__11072 (
            .O(N__46802),
            .I(N__46794));
    LocalMux I__11071 (
            .O(N__46799),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__11070 (
            .O(N__46794),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__11069 (
            .O(N__46789),
            .I(N__46785));
    InMux I__11068 (
            .O(N__46788),
            .I(N__46782));
    LocalMux I__11067 (
            .O(N__46785),
            .I(N__46779));
    LocalMux I__11066 (
            .O(N__46782),
            .I(N__46776));
    Span12Mux_v I__11065 (
            .O(N__46779),
            .I(N__46773));
    Span4Mux_h I__11064 (
            .O(N__46776),
            .I(N__46770));
    Odrv12 I__11063 (
            .O(N__46773),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    Odrv4 I__11062 (
            .O(N__46770),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    InMux I__11061 (
            .O(N__46765),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__11060 (
            .O(N__46762),
            .I(N__46757));
    InMux I__11059 (
            .O(N__46761),
            .I(N__46754));
    InMux I__11058 (
            .O(N__46760),
            .I(N__46751));
    LocalMux I__11057 (
            .O(N__46757),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__11056 (
            .O(N__46754),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__11055 (
            .O(N__46751),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__11054 (
            .O(N__46744),
            .I(N__46741));
    LocalMux I__11053 (
            .O(N__46741),
            .I(N__46737));
    InMux I__11052 (
            .O(N__46740),
            .I(N__46734));
    Span4Mux_v I__11051 (
            .O(N__46737),
            .I(N__46731));
    LocalMux I__11050 (
            .O(N__46734),
            .I(N__46728));
    Span4Mux_h I__11049 (
            .O(N__46731),
            .I(N__46725));
    Span4Mux_h I__11048 (
            .O(N__46728),
            .I(N__46722));
    Odrv4 I__11047 (
            .O(N__46725),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    Odrv4 I__11046 (
            .O(N__46722),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    InMux I__11045 (
            .O(N__46717),
            .I(bfn_18_24_0_));
    InMux I__11044 (
            .O(N__46714),
            .I(N__46709));
    InMux I__11043 (
            .O(N__46713),
            .I(N__46706));
    InMux I__11042 (
            .O(N__46712),
            .I(N__46703));
    LocalMux I__11041 (
            .O(N__46709),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__11040 (
            .O(N__46706),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__11039 (
            .O(N__46703),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__11038 (
            .O(N__46696),
            .I(N__46693));
    LocalMux I__11037 (
            .O(N__46693),
            .I(N__46689));
    InMux I__11036 (
            .O(N__46692),
            .I(N__46686));
    Span4Mux_v I__11035 (
            .O(N__46689),
            .I(N__46683));
    LocalMux I__11034 (
            .O(N__46686),
            .I(N__46680));
    Span4Mux_h I__11033 (
            .O(N__46683),
            .I(N__46677));
    Span4Mux_h I__11032 (
            .O(N__46680),
            .I(N__46674));
    Odrv4 I__11031 (
            .O(N__46677),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    Odrv4 I__11030 (
            .O(N__46674),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    InMux I__11029 (
            .O(N__46669),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__11028 (
            .O(N__46666),
            .I(N__46663));
    InMux I__11027 (
            .O(N__46663),
            .I(N__46660));
    LocalMux I__11026 (
            .O(N__46660),
            .I(N__46657));
    Span4Mux_h I__11025 (
            .O(N__46657),
            .I(N__46654));
    Span4Mux_v I__11024 (
            .O(N__46654),
            .I(N__46651));
    Odrv4 I__11023 (
            .O(N__46651),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    CEMux I__11022 (
            .O(N__46648),
            .I(N__46645));
    LocalMux I__11021 (
            .O(N__46645),
            .I(N__46638));
    CEMux I__11020 (
            .O(N__46644),
            .I(N__46635));
    CEMux I__11019 (
            .O(N__46643),
            .I(N__46632));
    CEMux I__11018 (
            .O(N__46642),
            .I(N__46629));
    CEMux I__11017 (
            .O(N__46641),
            .I(N__46625));
    Span4Mux_v I__11016 (
            .O(N__46638),
            .I(N__46622));
    LocalMux I__11015 (
            .O(N__46635),
            .I(N__46619));
    LocalMux I__11014 (
            .O(N__46632),
            .I(N__46616));
    LocalMux I__11013 (
            .O(N__46629),
            .I(N__46613));
    CEMux I__11012 (
            .O(N__46628),
            .I(N__46610));
    LocalMux I__11011 (
            .O(N__46625),
            .I(N__46607));
    Span4Mux_v I__11010 (
            .O(N__46622),
            .I(N__46604));
    Span4Mux_v I__11009 (
            .O(N__46619),
            .I(N__46601));
    Span4Mux_v I__11008 (
            .O(N__46616),
            .I(N__46598));
    Span4Mux_v I__11007 (
            .O(N__46613),
            .I(N__46593));
    LocalMux I__11006 (
            .O(N__46610),
            .I(N__46593));
    Span4Mux_h I__11005 (
            .O(N__46607),
            .I(N__46590));
    Sp12to4 I__11004 (
            .O(N__46604),
            .I(N__46583));
    Sp12to4 I__11003 (
            .O(N__46601),
            .I(N__46583));
    Sp12to4 I__11002 (
            .O(N__46598),
            .I(N__46583));
    Span4Mux_v I__11001 (
            .O(N__46593),
            .I(N__46580));
    Span4Mux_h I__11000 (
            .O(N__46590),
            .I(N__46577));
    Odrv12 I__10999 (
            .O(N__46583),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__10998 (
            .O(N__46580),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__10997 (
            .O(N__46577),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    CascadeMux I__10996 (
            .O(N__46570),
            .I(N__46566));
    InMux I__10995 (
            .O(N__46569),
            .I(N__46563));
    InMux I__10994 (
            .O(N__46566),
            .I(N__46560));
    LocalMux I__10993 (
            .O(N__46563),
            .I(N__46556));
    LocalMux I__10992 (
            .O(N__46560),
            .I(N__46553));
    CascadeMux I__10991 (
            .O(N__46559),
            .I(N__46550));
    Span4Mux_h I__10990 (
            .O(N__46556),
            .I(N__46547));
    Span12Mux_v I__10989 (
            .O(N__46553),
            .I(N__46544));
    InMux I__10988 (
            .O(N__46550),
            .I(N__46541));
    Span4Mux_h I__10987 (
            .O(N__46547),
            .I(N__46538));
    Odrv12 I__10986 (
            .O(N__46544),
            .I(measured_delay_tr_4));
    LocalMux I__10985 (
            .O(N__46541),
            .I(measured_delay_tr_4));
    Odrv4 I__10984 (
            .O(N__46538),
            .I(measured_delay_tr_4));
    InMux I__10983 (
            .O(N__46531),
            .I(N__46528));
    LocalMux I__10982 (
            .O(N__46528),
            .I(N__46523));
    InMux I__10981 (
            .O(N__46527),
            .I(N__46520));
    InMux I__10980 (
            .O(N__46526),
            .I(N__46517));
    Span4Mux_h I__10979 (
            .O(N__46523),
            .I(N__46513));
    LocalMux I__10978 (
            .O(N__46520),
            .I(N__46510));
    LocalMux I__10977 (
            .O(N__46517),
            .I(N__46507));
    InMux I__10976 (
            .O(N__46516),
            .I(N__46504));
    Span4Mux_h I__10975 (
            .O(N__46513),
            .I(N__46498));
    Span4Mux_h I__10974 (
            .O(N__46510),
            .I(N__46491));
    Span4Mux_v I__10973 (
            .O(N__46507),
            .I(N__46491));
    LocalMux I__10972 (
            .O(N__46504),
            .I(N__46491));
    InMux I__10971 (
            .O(N__46503),
            .I(N__46486));
    InMux I__10970 (
            .O(N__46502),
            .I(N__46486));
    InMux I__10969 (
            .O(N__46501),
            .I(N__46483));
    Odrv4 I__10968 (
            .O(N__46498),
            .I(\delay_measurement_inst.N_425 ));
    Odrv4 I__10967 (
            .O(N__46491),
            .I(\delay_measurement_inst.N_425 ));
    LocalMux I__10966 (
            .O(N__46486),
            .I(\delay_measurement_inst.N_425 ));
    LocalMux I__10965 (
            .O(N__46483),
            .I(\delay_measurement_inst.N_425 ));
    InMux I__10964 (
            .O(N__46474),
            .I(N__46470));
    InMux I__10963 (
            .O(N__46473),
            .I(N__46467));
    LocalMux I__10962 (
            .O(N__46470),
            .I(N__46464));
    LocalMux I__10961 (
            .O(N__46467),
            .I(N__46460));
    Span4Mux_h I__10960 (
            .O(N__46464),
            .I(N__46457));
    InMux I__10959 (
            .O(N__46463),
            .I(N__46454));
    Odrv4 I__10958 (
            .O(N__46460),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    Odrv4 I__10957 (
            .O(N__46457),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    LocalMux I__10956 (
            .O(N__46454),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    InMux I__10955 (
            .O(N__46447),
            .I(N__46443));
    InMux I__10954 (
            .O(N__46446),
            .I(N__46440));
    LocalMux I__10953 (
            .O(N__46443),
            .I(N__46433));
    LocalMux I__10952 (
            .O(N__46440),
            .I(N__46433));
    InMux I__10951 (
            .O(N__46439),
            .I(N__46430));
    InMux I__10950 (
            .O(N__46438),
            .I(N__46427));
    Span4Mux_v I__10949 (
            .O(N__46433),
            .I(N__46424));
    LocalMux I__10948 (
            .O(N__46430),
            .I(N__46419));
    LocalMux I__10947 (
            .O(N__46427),
            .I(N__46419));
    Span4Mux_h I__10946 (
            .O(N__46424),
            .I(N__46412));
    Span4Mux_v I__10945 (
            .O(N__46419),
            .I(N__46409));
    InMux I__10944 (
            .O(N__46418),
            .I(N__46402));
    InMux I__10943 (
            .O(N__46417),
            .I(N__46402));
    InMux I__10942 (
            .O(N__46416),
            .I(N__46402));
    InMux I__10941 (
            .O(N__46415),
            .I(N__46399));
    Odrv4 I__10940 (
            .O(N__46412),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    Odrv4 I__10939 (
            .O(N__46409),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    LocalMux I__10938 (
            .O(N__46402),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    LocalMux I__10937 (
            .O(N__46399),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    InMux I__10936 (
            .O(N__46390),
            .I(N__46387));
    LocalMux I__10935 (
            .O(N__46387),
            .I(N__46383));
    InMux I__10934 (
            .O(N__46386),
            .I(N__46379));
    Span4Mux_h I__10933 (
            .O(N__46383),
            .I(N__46376));
    InMux I__10932 (
            .O(N__46382),
            .I(N__46373));
    LocalMux I__10931 (
            .O(N__46379),
            .I(N__46370));
    Span4Mux_v I__10930 (
            .O(N__46376),
            .I(N__46367));
    LocalMux I__10929 (
            .O(N__46373),
            .I(N__46364));
    Span4Mux_h I__10928 (
            .O(N__46370),
            .I(N__46361));
    Odrv4 I__10927 (
            .O(N__46367),
            .I(measured_delay_tr_2));
    Odrv12 I__10926 (
            .O(N__46364),
            .I(measured_delay_tr_2));
    Odrv4 I__10925 (
            .O(N__46361),
            .I(measured_delay_tr_2));
    CEMux I__10924 (
            .O(N__46354),
            .I(N__46351));
    LocalMux I__10923 (
            .O(N__46351),
            .I(N__46346));
    CEMux I__10922 (
            .O(N__46350),
            .I(N__46340));
    CEMux I__10921 (
            .O(N__46349),
            .I(N__46337));
    Span4Mux_v I__10920 (
            .O(N__46346),
            .I(N__46334));
    CEMux I__10919 (
            .O(N__46345),
            .I(N__46331));
    CEMux I__10918 (
            .O(N__46344),
            .I(N__46328));
    CEMux I__10917 (
            .O(N__46343),
            .I(N__46325));
    LocalMux I__10916 (
            .O(N__46340),
            .I(N__46322));
    LocalMux I__10915 (
            .O(N__46337),
            .I(N__46319));
    Span4Mux_h I__10914 (
            .O(N__46334),
            .I(N__46314));
    LocalMux I__10913 (
            .O(N__46331),
            .I(N__46314));
    LocalMux I__10912 (
            .O(N__46328),
            .I(N__46311));
    LocalMux I__10911 (
            .O(N__46325),
            .I(N__46308));
    Span4Mux_v I__10910 (
            .O(N__46322),
            .I(N__46305));
    Span4Mux_v I__10909 (
            .O(N__46319),
            .I(N__46302));
    Span4Mux_h I__10908 (
            .O(N__46314),
            .I(N__46297));
    Span4Mux_h I__10907 (
            .O(N__46311),
            .I(N__46297));
    Span4Mux_h I__10906 (
            .O(N__46308),
            .I(N__46294));
    Odrv4 I__10905 (
            .O(N__46305),
            .I(\delay_measurement_inst.N_280_i_0 ));
    Odrv4 I__10904 (
            .O(N__46302),
            .I(\delay_measurement_inst.N_280_i_0 ));
    Odrv4 I__10903 (
            .O(N__46297),
            .I(\delay_measurement_inst.N_280_i_0 ));
    Odrv4 I__10902 (
            .O(N__46294),
            .I(\delay_measurement_inst.N_280_i_0 ));
    InMux I__10901 (
            .O(N__46285),
            .I(N__46279));
    InMux I__10900 (
            .O(N__46284),
            .I(N__46279));
    LocalMux I__10899 (
            .O(N__46279),
            .I(N__46276));
    Span4Mux_h I__10898 (
            .O(N__46276),
            .I(N__46273));
    Odrv4 I__10897 (
            .O(N__46273),
            .I(\delay_measurement_inst.N_286_1 ));
    InMux I__10896 (
            .O(N__46270),
            .I(N__46265));
    InMux I__10895 (
            .O(N__46269),
            .I(N__46262));
    InMux I__10894 (
            .O(N__46268),
            .I(N__46259));
    LocalMux I__10893 (
            .O(N__46265),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ));
    LocalMux I__10892 (
            .O(N__46262),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ));
    LocalMux I__10891 (
            .O(N__46259),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ));
    InMux I__10890 (
            .O(N__46252),
            .I(N__46245));
    InMux I__10889 (
            .O(N__46251),
            .I(N__46245));
    InMux I__10888 (
            .O(N__46250),
            .I(N__46242));
    LocalMux I__10887 (
            .O(N__46245),
            .I(N__46235));
    LocalMux I__10886 (
            .O(N__46242),
            .I(N__46232));
    InMux I__10885 (
            .O(N__46241),
            .I(N__46229));
    InMux I__10884 (
            .O(N__46240),
            .I(N__46226));
    InMux I__10883 (
            .O(N__46239),
            .I(N__46221));
    InMux I__10882 (
            .O(N__46238),
            .I(N__46221));
    Span4Mux_h I__10881 (
            .O(N__46235),
            .I(N__46216));
    Span4Mux_v I__10880 (
            .O(N__46232),
            .I(N__46213));
    LocalMux I__10879 (
            .O(N__46229),
            .I(N__46210));
    LocalMux I__10878 (
            .O(N__46226),
            .I(N__46205));
    LocalMux I__10877 (
            .O(N__46221),
            .I(N__46205));
    InMux I__10876 (
            .O(N__46220),
            .I(N__46202));
    InMux I__10875 (
            .O(N__46219),
            .I(N__46199));
    Span4Mux_v I__10874 (
            .O(N__46216),
            .I(N__46196));
    Span4Mux_h I__10873 (
            .O(N__46213),
            .I(N__46191));
    Span4Mux_v I__10872 (
            .O(N__46210),
            .I(N__46191));
    Span12Mux_h I__10871 (
            .O(N__46205),
            .I(N__46184));
    LocalMux I__10870 (
            .O(N__46202),
            .I(N__46184));
    LocalMux I__10869 (
            .O(N__46199),
            .I(N__46184));
    Odrv4 I__10868 (
            .O(N__46196),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    Odrv4 I__10867 (
            .O(N__46191),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    Odrv12 I__10866 (
            .O(N__46184),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    CascadeMux I__10865 (
            .O(N__46177),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16_cascade_ ));
    InMux I__10864 (
            .O(N__46174),
            .I(N__46171));
    LocalMux I__10863 (
            .O(N__46171),
            .I(\delay_measurement_inst.delay_tr_timer.N_415 ));
    CascadeMux I__10862 (
            .O(N__46168),
            .I(N__46162));
    CascadeMux I__10861 (
            .O(N__46167),
            .I(N__46159));
    CascadeMux I__10860 (
            .O(N__46166),
            .I(N__46156));
    InMux I__10859 (
            .O(N__46165),
            .I(N__46148));
    InMux I__10858 (
            .O(N__46162),
            .I(N__46148));
    InMux I__10857 (
            .O(N__46159),
            .I(N__46145));
    InMux I__10856 (
            .O(N__46156),
            .I(N__46142));
    InMux I__10855 (
            .O(N__46155),
            .I(N__46139));
    InMux I__10854 (
            .O(N__46154),
            .I(N__46136));
    CascadeMux I__10853 (
            .O(N__46153),
            .I(N__46132));
    LocalMux I__10852 (
            .O(N__46148),
            .I(N__46129));
    LocalMux I__10851 (
            .O(N__46145),
            .I(N__46122));
    LocalMux I__10850 (
            .O(N__46142),
            .I(N__46122));
    LocalMux I__10849 (
            .O(N__46139),
            .I(N__46122));
    LocalMux I__10848 (
            .O(N__46136),
            .I(N__46119));
    CascadeMux I__10847 (
            .O(N__46135),
            .I(N__46116));
    InMux I__10846 (
            .O(N__46132),
            .I(N__46113));
    Span4Mux_v I__10845 (
            .O(N__46129),
            .I(N__46108));
    Span4Mux_v I__10844 (
            .O(N__46122),
            .I(N__46108));
    Span4Mux_h I__10843 (
            .O(N__46119),
            .I(N__46105));
    InMux I__10842 (
            .O(N__46116),
            .I(N__46102));
    LocalMux I__10841 (
            .O(N__46113),
            .I(N__46099));
    Span4Mux_h I__10840 (
            .O(N__46108),
            .I(N__46094));
    Span4Mux_v I__10839 (
            .O(N__46105),
            .I(N__46094));
    LocalMux I__10838 (
            .O(N__46102),
            .I(\delay_measurement_inst.N_373 ));
    Odrv4 I__10837 (
            .O(N__46099),
            .I(\delay_measurement_inst.N_373 ));
    Odrv4 I__10836 (
            .O(N__46094),
            .I(\delay_measurement_inst.N_373 ));
    InMux I__10835 (
            .O(N__46087),
            .I(N__46083));
    CascadeMux I__10834 (
            .O(N__46086),
            .I(N__46080));
    LocalMux I__10833 (
            .O(N__46083),
            .I(N__46076));
    InMux I__10832 (
            .O(N__46080),
            .I(N__46073));
    InMux I__10831 (
            .O(N__46079),
            .I(N__46070));
    Span4Mux_h I__10830 (
            .O(N__46076),
            .I(N__46065));
    LocalMux I__10829 (
            .O(N__46073),
            .I(N__46065));
    LocalMux I__10828 (
            .O(N__46070),
            .I(N__46062));
    Span4Mux_h I__10827 (
            .O(N__46065),
            .I(N__46059));
    Span4Mux_h I__10826 (
            .O(N__46062),
            .I(N__46056));
    Odrv4 I__10825 (
            .O(N__46059),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    Odrv4 I__10824 (
            .O(N__46056),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    InMux I__10823 (
            .O(N__46051),
            .I(N__46048));
    LocalMux I__10822 (
            .O(N__46048),
            .I(N__46043));
    InMux I__10821 (
            .O(N__46047),
            .I(N__46040));
    InMux I__10820 (
            .O(N__46046),
            .I(N__46037));
    Odrv4 I__10819 (
            .O(N__46043),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__10818 (
            .O(N__46040),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__10817 (
            .O(N__46037),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__10816 (
            .O(N__46030),
            .I(N__46025));
    InMux I__10815 (
            .O(N__46029),
            .I(N__46022));
    InMux I__10814 (
            .O(N__46028),
            .I(N__46019));
    LocalMux I__10813 (
            .O(N__46025),
            .I(N__46016));
    LocalMux I__10812 (
            .O(N__46022),
            .I(N__46013));
    LocalMux I__10811 (
            .O(N__46019),
            .I(N__46010));
    Span4Mux_h I__10810 (
            .O(N__46016),
            .I(N__46007));
    Span4Mux_h I__10809 (
            .O(N__46013),
            .I(N__46004));
    Odrv12 I__10808 (
            .O(N__46010),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    Odrv4 I__10807 (
            .O(N__46007),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    Odrv4 I__10806 (
            .O(N__46004),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    InMux I__10805 (
            .O(N__45997),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__10804 (
            .O(N__45994),
            .I(N__45989));
    CascadeMux I__10803 (
            .O(N__45993),
            .I(N__45986));
    InMux I__10802 (
            .O(N__45992),
            .I(N__45983));
    InMux I__10801 (
            .O(N__45989),
            .I(N__45978));
    InMux I__10800 (
            .O(N__45986),
            .I(N__45978));
    LocalMux I__10799 (
            .O(N__45983),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__10798 (
            .O(N__45978),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    CascadeMux I__10797 (
            .O(N__45973),
            .I(N__45970));
    InMux I__10796 (
            .O(N__45970),
            .I(N__45965));
    InMux I__10795 (
            .O(N__45969),
            .I(N__45962));
    InMux I__10794 (
            .O(N__45968),
            .I(N__45959));
    LocalMux I__10793 (
            .O(N__45965),
            .I(N__45954));
    LocalMux I__10792 (
            .O(N__45962),
            .I(N__45954));
    LocalMux I__10791 (
            .O(N__45959),
            .I(N__45951));
    Span4Mux_h I__10790 (
            .O(N__45954),
            .I(N__45948));
    Span4Mux_h I__10789 (
            .O(N__45951),
            .I(N__45945));
    Odrv4 I__10788 (
            .O(N__45948),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    Odrv4 I__10787 (
            .O(N__45945),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    InMux I__10786 (
            .O(N__45940),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__10785 (
            .O(N__45937),
            .I(N__45934));
    LocalMux I__10784 (
            .O(N__45934),
            .I(N__45931));
    Span4Mux_v I__10783 (
            .O(N__45931),
            .I(N__45927));
    InMux I__10782 (
            .O(N__45930),
            .I(N__45924));
    Sp12to4 I__10781 (
            .O(N__45927),
            .I(N__45917));
    LocalMux I__10780 (
            .O(N__45924),
            .I(N__45917));
    InMux I__10779 (
            .O(N__45923),
            .I(N__45914));
    InMux I__10778 (
            .O(N__45922),
            .I(N__45911));
    Odrv12 I__10777 (
            .O(N__45917),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    LocalMux I__10776 (
            .O(N__45914),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    LocalMux I__10775 (
            .O(N__45911),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    InMux I__10774 (
            .O(N__45904),
            .I(N__45901));
    LocalMux I__10773 (
            .O(N__45901),
            .I(N__45897));
    InMux I__10772 (
            .O(N__45900),
            .I(N__45893));
    Span4Mux_h I__10771 (
            .O(N__45897),
            .I(N__45890));
    InMux I__10770 (
            .O(N__45896),
            .I(N__45887));
    LocalMux I__10769 (
            .O(N__45893),
            .I(N__45884));
    Odrv4 I__10768 (
            .O(N__45890),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    LocalMux I__10767 (
            .O(N__45887),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    Odrv4 I__10766 (
            .O(N__45884),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    CascadeMux I__10765 (
            .O(N__45877),
            .I(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_ ));
    InMux I__10764 (
            .O(N__45874),
            .I(N__45867));
    InMux I__10763 (
            .O(N__45873),
            .I(N__45862));
    InMux I__10762 (
            .O(N__45872),
            .I(N__45862));
    InMux I__10761 (
            .O(N__45871),
            .I(N__45858));
    InMux I__10760 (
            .O(N__45870),
            .I(N__45855));
    LocalMux I__10759 (
            .O(N__45867),
            .I(N__45852));
    LocalMux I__10758 (
            .O(N__45862),
            .I(N__45849));
    InMux I__10757 (
            .O(N__45861),
            .I(N__45846));
    LocalMux I__10756 (
            .O(N__45858),
            .I(N__45841));
    LocalMux I__10755 (
            .O(N__45855),
            .I(N__45841));
    Span4Mux_h I__10754 (
            .O(N__45852),
            .I(N__45838));
    Span4Mux_v I__10753 (
            .O(N__45849),
            .I(N__45833));
    LocalMux I__10752 (
            .O(N__45846),
            .I(N__45833));
    Span4Mux_h I__10751 (
            .O(N__45841),
            .I(N__45830));
    Odrv4 I__10750 (
            .O(N__45838),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__10749 (
            .O(N__45833),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__10748 (
            .O(N__45830),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__10747 (
            .O(N__45823),
            .I(N__45819));
    InMux I__10746 (
            .O(N__45822),
            .I(N__45815));
    InMux I__10745 (
            .O(N__45819),
            .I(N__45812));
    InMux I__10744 (
            .O(N__45818),
            .I(N__45809));
    LocalMux I__10743 (
            .O(N__45815),
            .I(N__45802));
    LocalMux I__10742 (
            .O(N__45812),
            .I(N__45802));
    LocalMux I__10741 (
            .O(N__45809),
            .I(N__45802));
    Span4Mux_v I__10740 (
            .O(N__45802),
            .I(N__45799));
    Odrv4 I__10739 (
            .O(N__45799),
            .I(il_max_comp2_D2));
    InMux I__10738 (
            .O(N__45796),
            .I(N__45793));
    LocalMux I__10737 (
            .O(N__45793),
            .I(N__45790));
    Odrv12 I__10736 (
            .O(N__45790),
            .I(\phase_controller_slave.N_213 ));
    InMux I__10735 (
            .O(N__45787),
            .I(N__45784));
    LocalMux I__10734 (
            .O(N__45784),
            .I(N__45781));
    Odrv12 I__10733 (
            .O(N__45781),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ));
    InMux I__10732 (
            .O(N__45778),
            .I(N__45775));
    LocalMux I__10731 (
            .O(N__45775),
            .I(N__45771));
    InMux I__10730 (
            .O(N__45774),
            .I(N__45768));
    Span4Mux_h I__10729 (
            .O(N__45771),
            .I(N__45763));
    LocalMux I__10728 (
            .O(N__45768),
            .I(N__45763));
    Odrv4 I__10727 (
            .O(N__45763),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__10726 (
            .O(N__45760),
            .I(N__45753));
    InMux I__10725 (
            .O(N__45759),
            .I(N__45750));
    InMux I__10724 (
            .O(N__45758),
            .I(N__45747));
    InMux I__10723 (
            .O(N__45757),
            .I(N__45744));
    InMux I__10722 (
            .O(N__45756),
            .I(N__45741));
    LocalMux I__10721 (
            .O(N__45753),
            .I(N__45736));
    LocalMux I__10720 (
            .O(N__45750),
            .I(N__45736));
    LocalMux I__10719 (
            .O(N__45747),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__10718 (
            .O(N__45744),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__10717 (
            .O(N__45741),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    Odrv4 I__10716 (
            .O(N__45736),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    InMux I__10715 (
            .O(N__45727),
            .I(N__45723));
    InMux I__10714 (
            .O(N__45726),
            .I(N__45720));
    LocalMux I__10713 (
            .O(N__45723),
            .I(N__45715));
    LocalMux I__10712 (
            .O(N__45720),
            .I(N__45715));
    Span4Mux_v I__10711 (
            .O(N__45715),
            .I(N__45710));
    InMux I__10710 (
            .O(N__45714),
            .I(N__45707));
    InMux I__10709 (
            .O(N__45713),
            .I(N__45704));
    Span4Mux_h I__10708 (
            .O(N__45710),
            .I(N__45701));
    LocalMux I__10707 (
            .O(N__45707),
            .I(N__45696));
    LocalMux I__10706 (
            .O(N__45704),
            .I(N__45696));
    Odrv4 I__10705 (
            .O(N__45701),
            .I(shift_flag_start));
    Odrv4 I__10704 (
            .O(N__45696),
            .I(shift_flag_start));
    IoInMux I__10703 (
            .O(N__45691),
            .I(N__45688));
    LocalMux I__10702 (
            .O(N__45688),
            .I(N__45685));
    Span4Mux_s1_v I__10701 (
            .O(N__45685),
            .I(N__45681));
    InMux I__10700 (
            .O(N__45684),
            .I(N__45678));
    Span4Mux_v I__10699 (
            .O(N__45681),
            .I(N__45673));
    LocalMux I__10698 (
            .O(N__45678),
            .I(N__45673));
    Span4Mux_v I__10697 (
            .O(N__45673),
            .I(N__45670));
    Sp12to4 I__10696 (
            .O(N__45670),
            .I(N__45667));
    Span12Mux_h I__10695 (
            .O(N__45667),
            .I(N__45663));
    InMux I__10694 (
            .O(N__45666),
            .I(N__45660));
    Odrv12 I__10693 (
            .O(N__45663),
            .I(s3_phy_c));
    LocalMux I__10692 (
            .O(N__45660),
            .I(s3_phy_c));
    CascadeMux I__10691 (
            .O(N__45655),
            .I(N__45644));
    CascadeMux I__10690 (
            .O(N__45654),
            .I(N__45640));
    CascadeMux I__10689 (
            .O(N__45653),
            .I(N__45637));
    CascadeMux I__10688 (
            .O(N__45652),
            .I(N__45634));
    CascadeMux I__10687 (
            .O(N__45651),
            .I(N__45631));
    CascadeMux I__10686 (
            .O(N__45650),
            .I(N__45622));
    CascadeMux I__10685 (
            .O(N__45649),
            .I(N__45615));
    CascadeMux I__10684 (
            .O(N__45648),
            .I(N__45612));
    CascadeMux I__10683 (
            .O(N__45647),
            .I(N__45609));
    InMux I__10682 (
            .O(N__45644),
            .I(N__45604));
    InMux I__10681 (
            .O(N__45643),
            .I(N__45604));
    InMux I__10680 (
            .O(N__45640),
            .I(N__45586));
    InMux I__10679 (
            .O(N__45637),
            .I(N__45586));
    InMux I__10678 (
            .O(N__45634),
            .I(N__45586));
    InMux I__10677 (
            .O(N__45631),
            .I(N__45586));
    InMux I__10676 (
            .O(N__45630),
            .I(N__45586));
    InMux I__10675 (
            .O(N__45629),
            .I(N__45586));
    InMux I__10674 (
            .O(N__45628),
            .I(N__45586));
    InMux I__10673 (
            .O(N__45627),
            .I(N__45586));
    InMux I__10672 (
            .O(N__45626),
            .I(N__45581));
    InMux I__10671 (
            .O(N__45625),
            .I(N__45581));
    InMux I__10670 (
            .O(N__45622),
            .I(N__45564));
    InMux I__10669 (
            .O(N__45621),
            .I(N__45564));
    InMux I__10668 (
            .O(N__45620),
            .I(N__45564));
    InMux I__10667 (
            .O(N__45619),
            .I(N__45564));
    InMux I__10666 (
            .O(N__45618),
            .I(N__45564));
    InMux I__10665 (
            .O(N__45615),
            .I(N__45564));
    InMux I__10664 (
            .O(N__45612),
            .I(N__45564));
    InMux I__10663 (
            .O(N__45609),
            .I(N__45564));
    LocalMux I__10662 (
            .O(N__45604),
            .I(N__45561));
    CascadeMux I__10661 (
            .O(N__45603),
            .I(N__45557));
    LocalMux I__10660 (
            .O(N__45586),
            .I(N__45552));
    LocalMux I__10659 (
            .O(N__45581),
            .I(N__45547));
    LocalMux I__10658 (
            .O(N__45564),
            .I(N__45547));
    Span4Mux_h I__10657 (
            .O(N__45561),
            .I(N__45544));
    InMux I__10656 (
            .O(N__45560),
            .I(N__45541));
    InMux I__10655 (
            .O(N__45557),
            .I(N__45538));
    InMux I__10654 (
            .O(N__45556),
            .I(N__45533));
    InMux I__10653 (
            .O(N__45555),
            .I(N__45533));
    Span4Mux_h I__10652 (
            .O(N__45552),
            .I(N__45528));
    Span4Mux_v I__10651 (
            .O(N__45547),
            .I(N__45528));
    Span4Mux_h I__10650 (
            .O(N__45544),
            .I(N__45523));
    LocalMux I__10649 (
            .O(N__45541),
            .I(N__45523));
    LocalMux I__10648 (
            .O(N__45538),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    LocalMux I__10647 (
            .O(N__45533),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__10646 (
            .O(N__45528),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__10645 (
            .O(N__45523),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    InMux I__10644 (
            .O(N__45514),
            .I(N__45481));
    InMux I__10643 (
            .O(N__45513),
            .I(N__45481));
    InMux I__10642 (
            .O(N__45512),
            .I(N__45481));
    InMux I__10641 (
            .O(N__45511),
            .I(N__45481));
    InMux I__10640 (
            .O(N__45510),
            .I(N__45481));
    InMux I__10639 (
            .O(N__45509),
            .I(N__45481));
    InMux I__10638 (
            .O(N__45508),
            .I(N__45481));
    InMux I__10637 (
            .O(N__45507),
            .I(N__45481));
    InMux I__10636 (
            .O(N__45506),
            .I(N__45464));
    InMux I__10635 (
            .O(N__45505),
            .I(N__45464));
    InMux I__10634 (
            .O(N__45504),
            .I(N__45464));
    InMux I__10633 (
            .O(N__45503),
            .I(N__45464));
    InMux I__10632 (
            .O(N__45502),
            .I(N__45464));
    InMux I__10631 (
            .O(N__45501),
            .I(N__45464));
    InMux I__10630 (
            .O(N__45500),
            .I(N__45464));
    InMux I__10629 (
            .O(N__45499),
            .I(N__45464));
    CascadeMux I__10628 (
            .O(N__45498),
            .I(N__45461));
    LocalMux I__10627 (
            .O(N__45481),
            .I(N__45451));
    LocalMux I__10626 (
            .O(N__45464),
            .I(N__45451));
    InMux I__10625 (
            .O(N__45461),
            .I(N__45446));
    InMux I__10624 (
            .O(N__45460),
            .I(N__45446));
    InMux I__10623 (
            .O(N__45459),
            .I(N__45443));
    InMux I__10622 (
            .O(N__45458),
            .I(N__45438));
    InMux I__10621 (
            .O(N__45457),
            .I(N__45438));
    InMux I__10620 (
            .O(N__45456),
            .I(N__45435));
    Span4Mux_v I__10619 (
            .O(N__45451),
            .I(N__45430));
    LocalMux I__10618 (
            .O(N__45446),
            .I(N__45427));
    LocalMux I__10617 (
            .O(N__45443),
            .I(N__45424));
    LocalMux I__10616 (
            .O(N__45438),
            .I(N__45419));
    LocalMux I__10615 (
            .O(N__45435),
            .I(N__45419));
    InMux I__10614 (
            .O(N__45434),
            .I(N__45414));
    InMux I__10613 (
            .O(N__45433),
            .I(N__45414));
    Sp12to4 I__10612 (
            .O(N__45430),
            .I(N__45409));
    Span12Mux_v I__10611 (
            .O(N__45427),
            .I(N__45409));
    Span4Mux_h I__10610 (
            .O(N__45424),
            .I(N__45406));
    Span4Mux_h I__10609 (
            .O(N__45419),
            .I(N__45403));
    LocalMux I__10608 (
            .O(N__45414),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv12 I__10607 (
            .O(N__45409),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__10606 (
            .O(N__45406),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__10605 (
            .O(N__45403),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    CascadeMux I__10604 (
            .O(N__45394),
            .I(N__45371));
    InMux I__10603 (
            .O(N__45393),
            .I(N__45366));
    InMux I__10602 (
            .O(N__45392),
            .I(N__45366));
    CascadeMux I__10601 (
            .O(N__45391),
            .I(N__45362));
    InMux I__10600 (
            .O(N__45390),
            .I(N__45344));
    InMux I__10599 (
            .O(N__45389),
            .I(N__45344));
    InMux I__10598 (
            .O(N__45388),
            .I(N__45344));
    InMux I__10597 (
            .O(N__45387),
            .I(N__45344));
    InMux I__10596 (
            .O(N__45386),
            .I(N__45344));
    InMux I__10595 (
            .O(N__45385),
            .I(N__45344));
    InMux I__10594 (
            .O(N__45384),
            .I(N__45344));
    InMux I__10593 (
            .O(N__45383),
            .I(N__45344));
    InMux I__10592 (
            .O(N__45382),
            .I(N__45327));
    InMux I__10591 (
            .O(N__45381),
            .I(N__45327));
    InMux I__10590 (
            .O(N__45380),
            .I(N__45327));
    InMux I__10589 (
            .O(N__45379),
            .I(N__45327));
    InMux I__10588 (
            .O(N__45378),
            .I(N__45327));
    InMux I__10587 (
            .O(N__45377),
            .I(N__45327));
    InMux I__10586 (
            .O(N__45376),
            .I(N__45327));
    InMux I__10585 (
            .O(N__45375),
            .I(N__45327));
    InMux I__10584 (
            .O(N__45374),
            .I(N__45323));
    InMux I__10583 (
            .O(N__45371),
            .I(N__45320));
    LocalMux I__10582 (
            .O(N__45366),
            .I(N__45317));
    InMux I__10581 (
            .O(N__45365),
            .I(N__45314));
    InMux I__10580 (
            .O(N__45362),
            .I(N__45309));
    InMux I__10579 (
            .O(N__45361),
            .I(N__45309));
    LocalMux I__10578 (
            .O(N__45344),
            .I(N__45304));
    LocalMux I__10577 (
            .O(N__45327),
            .I(N__45304));
    InMux I__10576 (
            .O(N__45326),
            .I(N__45301));
    LocalMux I__10575 (
            .O(N__45323),
            .I(N__45292));
    LocalMux I__10574 (
            .O(N__45320),
            .I(N__45292));
    Span4Mux_v I__10573 (
            .O(N__45317),
            .I(N__45292));
    LocalMux I__10572 (
            .O(N__45314),
            .I(N__45292));
    LocalMux I__10571 (
            .O(N__45309),
            .I(N__45287));
    Span4Mux_v I__10570 (
            .O(N__45304),
            .I(N__45287));
    LocalMux I__10569 (
            .O(N__45301),
            .I(N__45284));
    Span4Mux_h I__10568 (
            .O(N__45292),
            .I(N__45281));
    Odrv4 I__10567 (
            .O(N__45287),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv12 I__10566 (
            .O(N__45284),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__10565 (
            .O(N__45281),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    InMux I__10564 (
            .O(N__45274),
            .I(N__45271));
    LocalMux I__10563 (
            .O(N__45271),
            .I(N__45267));
    InMux I__10562 (
            .O(N__45270),
            .I(N__45264));
    Span4Mux_h I__10561 (
            .O(N__45267),
            .I(N__45260));
    LocalMux I__10560 (
            .O(N__45264),
            .I(N__45257));
    InMux I__10559 (
            .O(N__45263),
            .I(N__45254));
    Span4Mux_v I__10558 (
            .O(N__45260),
            .I(N__45250));
    Span12Mux_s11_v I__10557 (
            .O(N__45257),
            .I(N__45245));
    LocalMux I__10556 (
            .O(N__45254),
            .I(N__45245));
    InMux I__10555 (
            .O(N__45253),
            .I(N__45242));
    Odrv4 I__10554 (
            .O(N__45250),
            .I(measured_delay_tr_16));
    Odrv12 I__10553 (
            .O(N__45245),
            .I(measured_delay_tr_16));
    LocalMux I__10552 (
            .O(N__45242),
            .I(measured_delay_tr_16));
    InMux I__10551 (
            .O(N__45235),
            .I(N__45232));
    LocalMux I__10550 (
            .O(N__45232),
            .I(N__45229));
    Span4Mux_h I__10549 (
            .O(N__45229),
            .I(N__45226));
    Odrv4 I__10548 (
            .O(N__45226),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ));
    CEMux I__10547 (
            .O(N__45223),
            .I(N__45220));
    LocalMux I__10546 (
            .O(N__45220),
            .I(N__45216));
    CEMux I__10545 (
            .O(N__45219),
            .I(N__45213));
    Span4Mux_v I__10544 (
            .O(N__45216),
            .I(N__45206));
    LocalMux I__10543 (
            .O(N__45213),
            .I(N__45206));
    CEMux I__10542 (
            .O(N__45212),
            .I(N__45203));
    CEMux I__10541 (
            .O(N__45211),
            .I(N__45200));
    Span4Mux_h I__10540 (
            .O(N__45206),
            .I(N__45197));
    LocalMux I__10539 (
            .O(N__45203),
            .I(N__45193));
    LocalMux I__10538 (
            .O(N__45200),
            .I(N__45190));
    Span4Mux_h I__10537 (
            .O(N__45197),
            .I(N__45187));
    CEMux I__10536 (
            .O(N__45196),
            .I(N__45184));
    Span4Mux_h I__10535 (
            .O(N__45193),
            .I(N__45181));
    Span4Mux_h I__10534 (
            .O(N__45190),
            .I(N__45176));
    Span4Mux_v I__10533 (
            .O(N__45187),
            .I(N__45176));
    LocalMux I__10532 (
            .O(N__45184),
            .I(N__45173));
    Odrv4 I__10531 (
            .O(N__45181),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__10530 (
            .O(N__45176),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv12 I__10529 (
            .O(N__45173),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    CascadeMux I__10528 (
            .O(N__45166),
            .I(N__45161));
    CascadeMux I__10527 (
            .O(N__45165),
            .I(N__45158));
    InMux I__10526 (
            .O(N__45164),
            .I(N__45142));
    InMux I__10525 (
            .O(N__45161),
            .I(N__45142));
    InMux I__10524 (
            .O(N__45158),
            .I(N__45142));
    InMux I__10523 (
            .O(N__45157),
            .I(N__45142));
    InMux I__10522 (
            .O(N__45156),
            .I(N__45142));
    InMux I__10521 (
            .O(N__45155),
            .I(N__45138));
    InMux I__10520 (
            .O(N__45154),
            .I(N__45128));
    InMux I__10519 (
            .O(N__45153),
            .I(N__45125));
    LocalMux I__10518 (
            .O(N__45142),
            .I(N__45122));
    InMux I__10517 (
            .O(N__45141),
            .I(N__45119));
    LocalMux I__10516 (
            .O(N__45138),
            .I(N__45116));
    InMux I__10515 (
            .O(N__45137),
            .I(N__45113));
    InMux I__10514 (
            .O(N__45136),
            .I(N__45106));
    InMux I__10513 (
            .O(N__45135),
            .I(N__45106));
    InMux I__10512 (
            .O(N__45134),
            .I(N__45106));
    InMux I__10511 (
            .O(N__45133),
            .I(N__45099));
    InMux I__10510 (
            .O(N__45132),
            .I(N__45099));
    InMux I__10509 (
            .O(N__45131),
            .I(N__45099));
    LocalMux I__10508 (
            .O(N__45128),
            .I(N__45094));
    LocalMux I__10507 (
            .O(N__45125),
            .I(N__45094));
    Span4Mux_h I__10506 (
            .O(N__45122),
            .I(N__45089));
    LocalMux I__10505 (
            .O(N__45119),
            .I(N__45089));
    Span4Mux_v I__10504 (
            .O(N__45116),
            .I(N__45084));
    LocalMux I__10503 (
            .O(N__45113),
            .I(N__45084));
    LocalMux I__10502 (
            .O(N__45106),
            .I(N__45079));
    LocalMux I__10501 (
            .O(N__45099),
            .I(N__45079));
    Span4Mux_h I__10500 (
            .O(N__45094),
            .I(N__45076));
    Span4Mux_v I__10499 (
            .O(N__45089),
            .I(N__45071));
    Span4Mux_h I__10498 (
            .O(N__45084),
            .I(N__45071));
    Span4Mux_h I__10497 (
            .O(N__45079),
            .I(N__45068));
    Span4Mux_h I__10496 (
            .O(N__45076),
            .I(N__45065));
    Odrv4 I__10495 (
            .O(N__45071),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    Odrv4 I__10494 (
            .O(N__45068),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    Odrv4 I__10493 (
            .O(N__45065),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    CascadeMux I__10492 (
            .O(N__45058),
            .I(N__45054));
    InMux I__10491 (
            .O(N__45057),
            .I(N__45049));
    InMux I__10490 (
            .O(N__45054),
            .I(N__45044));
    InMux I__10489 (
            .O(N__45053),
            .I(N__45044));
    InMux I__10488 (
            .O(N__45052),
            .I(N__45041));
    LocalMux I__10487 (
            .O(N__45049),
            .I(N__45038));
    LocalMux I__10486 (
            .O(N__45044),
            .I(N__45035));
    LocalMux I__10485 (
            .O(N__45041),
            .I(N__45030));
    Span4Mux_v I__10484 (
            .O(N__45038),
            .I(N__45027));
    Span12Mux_h I__10483 (
            .O(N__45035),
            .I(N__45024));
    InMux I__10482 (
            .O(N__45034),
            .I(N__45019));
    InMux I__10481 (
            .O(N__45033),
            .I(N__45019));
    Span4Mux_h I__10480 (
            .O(N__45030),
            .I(N__45014));
    Span4Mux_h I__10479 (
            .O(N__45027),
            .I(N__45014));
    Odrv12 I__10478 (
            .O(N__45024),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ));
    LocalMux I__10477 (
            .O(N__45019),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ));
    Odrv4 I__10476 (
            .O(N__45014),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ));
    InMux I__10475 (
            .O(N__45007),
            .I(N__44995));
    InMux I__10474 (
            .O(N__45006),
            .I(N__44995));
    InMux I__10473 (
            .O(N__45005),
            .I(N__44995));
    InMux I__10472 (
            .O(N__45004),
            .I(N__44995));
    LocalMux I__10471 (
            .O(N__44995),
            .I(N__44990));
    InMux I__10470 (
            .O(N__44994),
            .I(N__44987));
    InMux I__10469 (
            .O(N__44993),
            .I(N__44984));
    Span4Mux_h I__10468 (
            .O(N__44990),
            .I(N__44979));
    LocalMux I__10467 (
            .O(N__44987),
            .I(N__44979));
    LocalMux I__10466 (
            .O(N__44984),
            .I(N__44976));
    Span4Mux_v I__10465 (
            .O(N__44979),
            .I(N__44969));
    Span4Mux_v I__10464 (
            .O(N__44976),
            .I(N__44966));
    InMux I__10463 (
            .O(N__44975),
            .I(N__44963));
    InMux I__10462 (
            .O(N__44974),
            .I(N__44956));
    InMux I__10461 (
            .O(N__44973),
            .I(N__44956));
    InMux I__10460 (
            .O(N__44972),
            .I(N__44956));
    Span4Mux_h I__10459 (
            .O(N__44969),
            .I(N__44953));
    Odrv4 I__10458 (
            .O(N__44966),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    LocalMux I__10457 (
            .O(N__44963),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    LocalMux I__10456 (
            .O(N__44956),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    Odrv4 I__10455 (
            .O(N__44953),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    InMux I__10454 (
            .O(N__44944),
            .I(N__44940));
    InMux I__10453 (
            .O(N__44943),
            .I(N__44937));
    LocalMux I__10452 (
            .O(N__44940),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__10451 (
            .O(N__44937),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__10450 (
            .O(N__44932),
            .I(N__44929));
    LocalMux I__10449 (
            .O(N__44929),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ));
    InMux I__10448 (
            .O(N__44926),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__10447 (
            .O(N__44923),
            .I(N__44919));
    InMux I__10446 (
            .O(N__44922),
            .I(N__44916));
    LocalMux I__10445 (
            .O(N__44919),
            .I(N__44913));
    LocalMux I__10444 (
            .O(N__44916),
            .I(N__44910));
    Odrv4 I__10443 (
            .O(N__44913),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__10442 (
            .O(N__44910),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__10441 (
            .O(N__44905),
            .I(N__44902));
    InMux I__10440 (
            .O(N__44902),
            .I(N__44899));
    LocalMux I__10439 (
            .O(N__44899),
            .I(N__44896));
    Odrv4 I__10438 (
            .O(N__44896),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ));
    InMux I__10437 (
            .O(N__44893),
            .I(bfn_18_10_0_));
    InMux I__10436 (
            .O(N__44890),
            .I(N__44886));
    InMux I__10435 (
            .O(N__44889),
            .I(N__44883));
    LocalMux I__10434 (
            .O(N__44886),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__10433 (
            .O(N__44883),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__10432 (
            .O(N__44878),
            .I(N__44875));
    LocalMux I__10431 (
            .O(N__44875),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ));
    InMux I__10430 (
            .O(N__44872),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__10429 (
            .O(N__44869),
            .I(N__44866));
    LocalMux I__10428 (
            .O(N__44866),
            .I(N__44862));
    InMux I__10427 (
            .O(N__44865),
            .I(N__44859));
    Span4Mux_h I__10426 (
            .O(N__44862),
            .I(N__44854));
    LocalMux I__10425 (
            .O(N__44859),
            .I(N__44854));
    Span4Mux_h I__10424 (
            .O(N__44854),
            .I(N__44851));
    Odrv4 I__10423 (
            .O(N__44851),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__10422 (
            .O(N__44848),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__10421 (
            .O(N__44845),
            .I(N__44842));
    LocalMux I__10420 (
            .O(N__44842),
            .I(N__44839));
    Span4Mux_v I__10419 (
            .O(N__44839),
            .I(N__44836));
    Odrv4 I__10418 (
            .O(N__44836),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ));
    InMux I__10417 (
            .O(N__44833),
            .I(N__44830));
    LocalMux I__10416 (
            .O(N__44830),
            .I(N__44827));
    Odrv4 I__10415 (
            .O(N__44827),
            .I(\phase_controller_slave.start_timer_hc_0_sqmuxa ));
    InMux I__10414 (
            .O(N__44824),
            .I(N__44818));
    InMux I__10413 (
            .O(N__44823),
            .I(N__44811));
    InMux I__10412 (
            .O(N__44822),
            .I(N__44811));
    InMux I__10411 (
            .O(N__44821),
            .I(N__44811));
    LocalMux I__10410 (
            .O(N__44818),
            .I(\phase_controller_slave.hc_time_passed ));
    LocalMux I__10409 (
            .O(N__44811),
            .I(\phase_controller_slave.hc_time_passed ));
    CascadeMux I__10408 (
            .O(N__44806),
            .I(N__44802));
    CascadeMux I__10407 (
            .O(N__44805),
            .I(N__44799));
    InMux I__10406 (
            .O(N__44802),
            .I(N__44795));
    InMux I__10405 (
            .O(N__44799),
            .I(N__44790));
    InMux I__10404 (
            .O(N__44798),
            .I(N__44790));
    LocalMux I__10403 (
            .O(N__44795),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    LocalMux I__10402 (
            .O(N__44790),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    IoInMux I__10401 (
            .O(N__44785),
            .I(N__44782));
    LocalMux I__10400 (
            .O(N__44782),
            .I(N__44779));
    IoSpan4Mux I__10399 (
            .O(N__44779),
            .I(N__44776));
    Span4Mux_s3_v I__10398 (
            .O(N__44776),
            .I(N__44773));
    Span4Mux_v I__10397 (
            .O(N__44773),
            .I(N__44770));
    Sp12to4 I__10396 (
            .O(N__44770),
            .I(N__44767));
    Span12Mux_h I__10395 (
            .O(N__44767),
            .I(N__44763));
    CascadeMux I__10394 (
            .O(N__44766),
            .I(N__44760));
    Span12Mux_v I__10393 (
            .O(N__44763),
            .I(N__44757));
    InMux I__10392 (
            .O(N__44760),
            .I(N__44754));
    Odrv12 I__10391 (
            .O(N__44757),
            .I(s4_phy_c));
    LocalMux I__10390 (
            .O(N__44754),
            .I(s4_phy_c));
    InMux I__10389 (
            .O(N__44749),
            .I(N__44745));
    InMux I__10388 (
            .O(N__44748),
            .I(N__44742));
    LocalMux I__10387 (
            .O(N__44745),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__10386 (
            .O(N__44742),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__10385 (
            .O(N__44737),
            .I(N__44734));
    LocalMux I__10384 (
            .O(N__44734),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ));
    InMux I__10383 (
            .O(N__44731),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__10382 (
            .O(N__44728),
            .I(N__44725));
    LocalMux I__10381 (
            .O(N__44725),
            .I(N__44722));
    Span4Mux_h I__10380 (
            .O(N__44722),
            .I(N__44718));
    InMux I__10379 (
            .O(N__44721),
            .I(N__44715));
    Odrv4 I__10378 (
            .O(N__44718),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__10377 (
            .O(N__44715),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__10376 (
            .O(N__44710),
            .I(N__44707));
    LocalMux I__10375 (
            .O(N__44707),
            .I(N__44704));
    Span4Mux_h I__10374 (
            .O(N__44704),
            .I(N__44701));
    Odrv4 I__10373 (
            .O(N__44701),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ));
    InMux I__10372 (
            .O(N__44698),
            .I(bfn_18_9_0_));
    InMux I__10371 (
            .O(N__44695),
            .I(N__44691));
    InMux I__10370 (
            .O(N__44694),
            .I(N__44688));
    LocalMux I__10369 (
            .O(N__44691),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__10368 (
            .O(N__44688),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__10367 (
            .O(N__44683),
            .I(N__44680));
    LocalMux I__10366 (
            .O(N__44680),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ));
    InMux I__10365 (
            .O(N__44677),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__10364 (
            .O(N__44674),
            .I(N__44670));
    InMux I__10363 (
            .O(N__44673),
            .I(N__44667));
    LocalMux I__10362 (
            .O(N__44670),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__10361 (
            .O(N__44667),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__10360 (
            .O(N__44662),
            .I(N__44659));
    LocalMux I__10359 (
            .O(N__44659),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ));
    InMux I__10358 (
            .O(N__44656),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__10357 (
            .O(N__44653),
            .I(N__44649));
    InMux I__10356 (
            .O(N__44652),
            .I(N__44646));
    LocalMux I__10355 (
            .O(N__44649),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__10354 (
            .O(N__44646),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__10353 (
            .O(N__44641),
            .I(N__44638));
    LocalMux I__10352 (
            .O(N__44638),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ));
    InMux I__10351 (
            .O(N__44635),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__10350 (
            .O(N__44632),
            .I(N__44628));
    InMux I__10349 (
            .O(N__44631),
            .I(N__44625));
    LocalMux I__10348 (
            .O(N__44628),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__10347 (
            .O(N__44625),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__10346 (
            .O(N__44620),
            .I(N__44617));
    LocalMux I__10345 (
            .O(N__44617),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ));
    InMux I__10344 (
            .O(N__44614),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__10343 (
            .O(N__44611),
            .I(N__44607));
    InMux I__10342 (
            .O(N__44610),
            .I(N__44604));
    LocalMux I__10341 (
            .O(N__44607),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__10340 (
            .O(N__44604),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__10339 (
            .O(N__44599),
            .I(N__44596));
    LocalMux I__10338 (
            .O(N__44596),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ));
    InMux I__10337 (
            .O(N__44593),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__10336 (
            .O(N__44590),
            .I(N__44586));
    InMux I__10335 (
            .O(N__44589),
            .I(N__44583));
    LocalMux I__10334 (
            .O(N__44586),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__10333 (
            .O(N__44583),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__10332 (
            .O(N__44578),
            .I(N__44575));
    LocalMux I__10331 (
            .O(N__44575),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ));
    InMux I__10330 (
            .O(N__44572),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__10329 (
            .O(N__44569),
            .I(N__44531));
    InMux I__10328 (
            .O(N__44568),
            .I(N__44531));
    InMux I__10327 (
            .O(N__44567),
            .I(N__44531));
    InMux I__10326 (
            .O(N__44566),
            .I(N__44531));
    InMux I__10325 (
            .O(N__44565),
            .I(N__44526));
    InMux I__10324 (
            .O(N__44564),
            .I(N__44526));
    InMux I__10323 (
            .O(N__44563),
            .I(N__44517));
    InMux I__10322 (
            .O(N__44562),
            .I(N__44517));
    InMux I__10321 (
            .O(N__44561),
            .I(N__44517));
    InMux I__10320 (
            .O(N__44560),
            .I(N__44517));
    InMux I__10319 (
            .O(N__44559),
            .I(N__44508));
    InMux I__10318 (
            .O(N__44558),
            .I(N__44508));
    InMux I__10317 (
            .O(N__44557),
            .I(N__44508));
    InMux I__10316 (
            .O(N__44556),
            .I(N__44508));
    InMux I__10315 (
            .O(N__44555),
            .I(N__44499));
    InMux I__10314 (
            .O(N__44554),
            .I(N__44499));
    InMux I__10313 (
            .O(N__44553),
            .I(N__44499));
    InMux I__10312 (
            .O(N__44552),
            .I(N__44499));
    InMux I__10311 (
            .O(N__44551),
            .I(N__44490));
    InMux I__10310 (
            .O(N__44550),
            .I(N__44490));
    InMux I__10309 (
            .O(N__44549),
            .I(N__44490));
    InMux I__10308 (
            .O(N__44548),
            .I(N__44490));
    InMux I__10307 (
            .O(N__44547),
            .I(N__44481));
    InMux I__10306 (
            .O(N__44546),
            .I(N__44481));
    InMux I__10305 (
            .O(N__44545),
            .I(N__44481));
    InMux I__10304 (
            .O(N__44544),
            .I(N__44481));
    InMux I__10303 (
            .O(N__44543),
            .I(N__44472));
    InMux I__10302 (
            .O(N__44542),
            .I(N__44472));
    InMux I__10301 (
            .O(N__44541),
            .I(N__44472));
    InMux I__10300 (
            .O(N__44540),
            .I(N__44472));
    LocalMux I__10299 (
            .O(N__44531),
            .I(N__44461));
    LocalMux I__10298 (
            .O(N__44526),
            .I(N__44461));
    LocalMux I__10297 (
            .O(N__44517),
            .I(N__44461));
    LocalMux I__10296 (
            .O(N__44508),
            .I(N__44461));
    LocalMux I__10295 (
            .O(N__44499),
            .I(N__44461));
    LocalMux I__10294 (
            .O(N__44490),
            .I(N__44458));
    LocalMux I__10293 (
            .O(N__44481),
            .I(N__44451));
    LocalMux I__10292 (
            .O(N__44472),
            .I(N__44451));
    Span4Mux_v I__10291 (
            .O(N__44461),
            .I(N__44451));
    Odrv12 I__10290 (
            .O(N__44458),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__10289 (
            .O(N__44451),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__10288 (
            .O(N__44446),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__10287 (
            .O(N__44443),
            .I(N__44437));
    CEMux I__10286 (
            .O(N__44442),
            .I(N__44434));
    CEMux I__10285 (
            .O(N__44441),
            .I(N__44431));
    CEMux I__10284 (
            .O(N__44440),
            .I(N__44428));
    LocalMux I__10283 (
            .O(N__44437),
            .I(N__44425));
    LocalMux I__10282 (
            .O(N__44434),
            .I(N__44422));
    LocalMux I__10281 (
            .O(N__44431),
            .I(N__44417));
    LocalMux I__10280 (
            .O(N__44428),
            .I(N__44417));
    Span4Mux_v I__10279 (
            .O(N__44425),
            .I(N__44410));
    Span4Mux_v I__10278 (
            .O(N__44422),
            .I(N__44410));
    Span4Mux_v I__10277 (
            .O(N__44417),
            .I(N__44410));
    Odrv4 I__10276 (
            .O(N__44410),
            .I(\delay_measurement_inst.delay_tr_timer.N_339_i ));
    InMux I__10275 (
            .O(N__44407),
            .I(N__44404));
    LocalMux I__10274 (
            .O(N__44404),
            .I(N__44401));
    Odrv4 I__10273 (
            .O(N__44401),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    CascadeMux I__10272 (
            .O(N__44398),
            .I(N__44394));
    InMux I__10271 (
            .O(N__44397),
            .I(N__44390));
    InMux I__10270 (
            .O(N__44394),
            .I(N__44387));
    InMux I__10269 (
            .O(N__44393),
            .I(N__44384));
    LocalMux I__10268 (
            .O(N__44390),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__10267 (
            .O(N__44387),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__10266 (
            .O(N__44384),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__10265 (
            .O(N__44377),
            .I(N__44373));
    InMux I__10264 (
            .O(N__44376),
            .I(N__44370));
    LocalMux I__10263 (
            .O(N__44373),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__10262 (
            .O(N__44370),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__10261 (
            .O(N__44365),
            .I(N__44362));
    LocalMux I__10260 (
            .O(N__44362),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ));
    InMux I__10259 (
            .O(N__44359),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__10258 (
            .O(N__44356),
            .I(N__44353));
    LocalMux I__10257 (
            .O(N__44353),
            .I(N__44350));
    Span4Mux_h I__10256 (
            .O(N__44350),
            .I(N__44347));
    Odrv4 I__10255 (
            .O(N__44347),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ));
    CascadeMux I__10254 (
            .O(N__44344),
            .I(N__44341));
    InMux I__10253 (
            .O(N__44341),
            .I(N__44337));
    InMux I__10252 (
            .O(N__44340),
            .I(N__44334));
    LocalMux I__10251 (
            .O(N__44337),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__10250 (
            .O(N__44334),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__10249 (
            .O(N__44329),
            .I(N__44326));
    LocalMux I__10248 (
            .O(N__44326),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ));
    InMux I__10247 (
            .O(N__44323),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__10246 (
            .O(N__44320),
            .I(N__44316));
    InMux I__10245 (
            .O(N__44319),
            .I(N__44313));
    LocalMux I__10244 (
            .O(N__44316),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__10243 (
            .O(N__44313),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__10242 (
            .O(N__44308),
            .I(N__44305));
    InMux I__10241 (
            .O(N__44305),
            .I(N__44302));
    LocalMux I__10240 (
            .O(N__44302),
            .I(N__44299));
    Odrv4 I__10239 (
            .O(N__44299),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ));
    InMux I__10238 (
            .O(N__44296),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__10237 (
            .O(N__44293),
            .I(N__44289));
    InMux I__10236 (
            .O(N__44292),
            .I(N__44286));
    LocalMux I__10235 (
            .O(N__44289),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__10234 (
            .O(N__44286),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__10233 (
            .O(N__44281),
            .I(N__44278));
    InMux I__10232 (
            .O(N__44278),
            .I(N__44275));
    LocalMux I__10231 (
            .O(N__44275),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ));
    InMux I__10230 (
            .O(N__44272),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__10229 (
            .O(N__44269),
            .I(N__44265));
    InMux I__10228 (
            .O(N__44268),
            .I(N__44262));
    LocalMux I__10227 (
            .O(N__44265),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__10226 (
            .O(N__44262),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__10225 (
            .O(N__44257),
            .I(N__44254));
    LocalMux I__10224 (
            .O(N__44254),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ));
    InMux I__10223 (
            .O(N__44251),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__10222 (
            .O(N__44248),
            .I(N__44245));
    LocalMux I__10221 (
            .O(N__44245),
            .I(N__44241));
    InMux I__10220 (
            .O(N__44244),
            .I(N__44238));
    Span4Mux_h I__10219 (
            .O(N__44241),
            .I(N__44235));
    LocalMux I__10218 (
            .O(N__44238),
            .I(N__44232));
    Odrv4 I__10217 (
            .O(N__44235),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__10216 (
            .O(N__44232),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__10215 (
            .O(N__44227),
            .I(N__44224));
    LocalMux I__10214 (
            .O(N__44224),
            .I(N__44221));
    Span4Mux_h I__10213 (
            .O(N__44221),
            .I(N__44218));
    Odrv4 I__10212 (
            .O(N__44218),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ));
    InMux I__10211 (
            .O(N__44215),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__10210 (
            .O(N__44212),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__10209 (
            .O(N__44209),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__10208 (
            .O(N__44206),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__10207 (
            .O(N__44203),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__10206 (
            .O(N__44200),
            .I(bfn_17_26_0_));
    InMux I__10205 (
            .O(N__44197),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__10204 (
            .O(N__44194),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__10203 (
            .O(N__44191),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__10202 (
            .O(N__44188),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__10201 (
            .O(N__44185),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__10200 (
            .O(N__44182),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__10199 (
            .O(N__44179),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__10198 (
            .O(N__44176),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__10197 (
            .O(N__44173),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__10196 (
            .O(N__44170),
            .I(bfn_17_25_0_));
    InMux I__10195 (
            .O(N__44167),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__10194 (
            .O(N__44164),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__10193 (
            .O(N__44161),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__10192 (
            .O(N__44158),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__10191 (
            .O(N__44155),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__10190 (
            .O(N__44152),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__10189 (
            .O(N__44149),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__10188 (
            .O(N__44146),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__10187 (
            .O(N__44143),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__10186 (
            .O(N__44140),
            .I(bfn_17_24_0_));
    InMux I__10185 (
            .O(N__44137),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__10184 (
            .O(N__44134),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__10183 (
            .O(N__44131),
            .I(N__44128));
    LocalMux I__10182 (
            .O(N__44128),
            .I(N__44124));
    InMux I__10181 (
            .O(N__44127),
            .I(N__44121));
    Odrv4 I__10180 (
            .O(N__44124),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__10179 (
            .O(N__44121),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__10178 (
            .O(N__44116),
            .I(N__44111));
    InMux I__10177 (
            .O(N__44115),
            .I(N__44108));
    InMux I__10176 (
            .O(N__44114),
            .I(N__44105));
    LocalMux I__10175 (
            .O(N__44111),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__10174 (
            .O(N__44108),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__10173 (
            .O(N__44105),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__10172 (
            .O(N__44098),
            .I(N__44094));
    InMux I__10171 (
            .O(N__44097),
            .I(N__44091));
    LocalMux I__10170 (
            .O(N__44094),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ));
    LocalMux I__10169 (
            .O(N__44091),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ));
    CascadeMux I__10168 (
            .O(N__44086),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_ ));
    InMux I__10167 (
            .O(N__44083),
            .I(N__44068));
    InMux I__10166 (
            .O(N__44082),
            .I(N__44068));
    InMux I__10165 (
            .O(N__44081),
            .I(N__44068));
    InMux I__10164 (
            .O(N__44080),
            .I(N__44068));
    InMux I__10163 (
            .O(N__44079),
            .I(N__44068));
    LocalMux I__10162 (
            .O(N__44068),
            .I(N__44065));
    Span4Mux_h I__10161 (
            .O(N__44065),
            .I(N__44062));
    Odrv4 I__10160 (
            .O(N__44062),
            .I(\delay_measurement_inst.N_409_1 ));
    InMux I__10159 (
            .O(N__44059),
            .I(N__44053));
    InMux I__10158 (
            .O(N__44058),
            .I(N__44050));
    InMux I__10157 (
            .O(N__44057),
            .I(N__44045));
    InMux I__10156 (
            .O(N__44056),
            .I(N__44045));
    LocalMux I__10155 (
            .O(N__44053),
            .I(N__44042));
    LocalMux I__10154 (
            .O(N__44050),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__10153 (
            .O(N__44045),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__10152 (
            .O(N__44042),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    CascadeMux I__10151 (
            .O(N__44035),
            .I(N__44032));
    InMux I__10150 (
            .O(N__44032),
            .I(N__44029));
    LocalMux I__10149 (
            .O(N__44029),
            .I(N__44026));
    Span4Mux_h I__10148 (
            .O(N__44026),
            .I(N__44023));
    Odrv4 I__10147 (
            .O(N__44023),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__10146 (
            .O(N__44020),
            .I(bfn_17_23_0_));
    InMux I__10145 (
            .O(N__44017),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__10144 (
            .O(N__44014),
            .I(N__44011));
    LocalMux I__10143 (
            .O(N__44011),
            .I(N__44007));
    InMux I__10142 (
            .O(N__44010),
            .I(N__44003));
    Span4Mux_v I__10141 (
            .O(N__44007),
            .I(N__44000));
    InMux I__10140 (
            .O(N__44006),
            .I(N__43997));
    LocalMux I__10139 (
            .O(N__44003),
            .I(N__43994));
    Odrv4 I__10138 (
            .O(N__44000),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__10137 (
            .O(N__43997),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    Odrv12 I__10136 (
            .O(N__43994),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    InMux I__10135 (
            .O(N__43987),
            .I(N__43982));
    InMux I__10134 (
            .O(N__43986),
            .I(N__43976));
    InMux I__10133 (
            .O(N__43985),
            .I(N__43976));
    LocalMux I__10132 (
            .O(N__43982),
            .I(N__43973));
    InMux I__10131 (
            .O(N__43981),
            .I(N__43970));
    LocalMux I__10130 (
            .O(N__43976),
            .I(N__43967));
    Sp12to4 I__10129 (
            .O(N__43973),
            .I(N__43962));
    LocalMux I__10128 (
            .O(N__43970),
            .I(N__43962));
    Span12Mux_v I__10127 (
            .O(N__43967),
            .I(N__43959));
    Span12Mux_v I__10126 (
            .O(N__43962),
            .I(N__43956));
    Odrv12 I__10125 (
            .O(N__43959),
            .I(delay_tr_d2));
    Odrv12 I__10124 (
            .O(N__43956),
            .I(delay_tr_d2));
    InMux I__10123 (
            .O(N__43951),
            .I(N__43948));
    LocalMux I__10122 (
            .O(N__43948),
            .I(N__43944));
    InMux I__10121 (
            .O(N__43947),
            .I(N__43940));
    Span4Mux_h I__10120 (
            .O(N__43944),
            .I(N__43937));
    InMux I__10119 (
            .O(N__43943),
            .I(N__43934));
    LocalMux I__10118 (
            .O(N__43940),
            .I(N__43931));
    Odrv4 I__10117 (
            .O(N__43937),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__10116 (
            .O(N__43934),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    Odrv12 I__10115 (
            .O(N__43931),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    CascadeMux I__10114 (
            .O(N__43924),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4_cascade_ ));
    InMux I__10113 (
            .O(N__43921),
            .I(N__43918));
    LocalMux I__10112 (
            .O(N__43918),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5 ));
    CascadeMux I__10111 (
            .O(N__43915),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_ ));
    InMux I__10110 (
            .O(N__43912),
            .I(N__43909));
    LocalMux I__10109 (
            .O(N__43909),
            .I(N__43905));
    InMux I__10108 (
            .O(N__43908),
            .I(N__43902));
    Span4Mux_h I__10107 (
            .O(N__43905),
            .I(N__43899));
    LocalMux I__10106 (
            .O(N__43902),
            .I(N__43896));
    Span4Mux_h I__10105 (
            .O(N__43899),
            .I(N__43893));
    Odrv12 I__10104 (
            .O(N__43896),
            .I(\delay_measurement_inst.tr_state_RNIMR6LZ0Z_0 ));
    Odrv4 I__10103 (
            .O(N__43893),
            .I(\delay_measurement_inst.tr_state_RNIMR6LZ0Z_0 ));
    CascadeMux I__10102 (
            .O(N__43888),
            .I(\delay_measurement_inst.delay_tr_timer.N_390_cascade_ ));
    InMux I__10101 (
            .O(N__43885),
            .I(N__43882));
    LocalMux I__10100 (
            .O(N__43882),
            .I(\delay_measurement_inst.delay_tr_timer.N_379 ));
    InMux I__10099 (
            .O(N__43879),
            .I(N__43873));
    InMux I__10098 (
            .O(N__43878),
            .I(N__43870));
    InMux I__10097 (
            .O(N__43877),
            .I(N__43865));
    InMux I__10096 (
            .O(N__43876),
            .I(N__43865));
    LocalMux I__10095 (
            .O(N__43873),
            .I(N__43860));
    LocalMux I__10094 (
            .O(N__43870),
            .I(N__43860));
    LocalMux I__10093 (
            .O(N__43865),
            .I(N__43857));
    Span4Mux_v I__10092 (
            .O(N__43860),
            .I(N__43852));
    Span4Mux_v I__10091 (
            .O(N__43857),
            .I(N__43852));
    Span4Mux_h I__10090 (
            .O(N__43852),
            .I(N__43848));
    InMux I__10089 (
            .O(N__43851),
            .I(N__43845));
    Odrv4 I__10088 (
            .O(N__43848),
            .I(\delay_measurement_inst.N_280_i ));
    LocalMux I__10087 (
            .O(N__43845),
            .I(\delay_measurement_inst.N_280_i ));
    InMux I__10086 (
            .O(N__43840),
            .I(bfn_17_14_0_));
    CascadeMux I__10085 (
            .O(N__43837),
            .I(N__43833));
    InMux I__10084 (
            .O(N__43836),
            .I(N__43830));
    InMux I__10083 (
            .O(N__43833),
            .I(N__43827));
    LocalMux I__10082 (
            .O(N__43830),
            .I(N__43821));
    LocalMux I__10081 (
            .O(N__43827),
            .I(N__43821));
    InMux I__10080 (
            .O(N__43826),
            .I(N__43818));
    Span4Mux_v I__10079 (
            .O(N__43821),
            .I(N__43815));
    LocalMux I__10078 (
            .O(N__43818),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__10077 (
            .O(N__43815),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__10076 (
            .O(N__43810),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__10075 (
            .O(N__43807),
            .I(N__43803));
    CascadeMux I__10074 (
            .O(N__43806),
            .I(N__43800));
    InMux I__10073 (
            .O(N__43803),
            .I(N__43794));
    InMux I__10072 (
            .O(N__43800),
            .I(N__43794));
    InMux I__10071 (
            .O(N__43799),
            .I(N__43791));
    LocalMux I__10070 (
            .O(N__43794),
            .I(N__43788));
    LocalMux I__10069 (
            .O(N__43791),
            .I(N__43783));
    Span4Mux_v I__10068 (
            .O(N__43788),
            .I(N__43783));
    Odrv4 I__10067 (
            .O(N__43783),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__10066 (
            .O(N__43780),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    CascadeMux I__10065 (
            .O(N__43777),
            .I(N__43773));
    InMux I__10064 (
            .O(N__43776),
            .I(N__43769));
    InMux I__10063 (
            .O(N__43773),
            .I(N__43766));
    InMux I__10062 (
            .O(N__43772),
            .I(N__43763));
    LocalMux I__10061 (
            .O(N__43769),
            .I(N__43758));
    LocalMux I__10060 (
            .O(N__43766),
            .I(N__43758));
    LocalMux I__10059 (
            .O(N__43763),
            .I(N__43753));
    Span4Mux_v I__10058 (
            .O(N__43758),
            .I(N__43753));
    Odrv4 I__10057 (
            .O(N__43753),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__10056 (
            .O(N__43750),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__10055 (
            .O(N__43747),
            .I(N__43744));
    LocalMux I__10054 (
            .O(N__43744),
            .I(N__43740));
    InMux I__10053 (
            .O(N__43743),
            .I(N__43737));
    Span4Mux_v I__10052 (
            .O(N__43740),
            .I(N__43734));
    LocalMux I__10051 (
            .O(N__43737),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__10050 (
            .O(N__43734),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__10049 (
            .O(N__43729),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__10048 (
            .O(N__43726),
            .I(N__43694));
    InMux I__10047 (
            .O(N__43725),
            .I(N__43694));
    InMux I__10046 (
            .O(N__43724),
            .I(N__43694));
    InMux I__10045 (
            .O(N__43723),
            .I(N__43694));
    InMux I__10044 (
            .O(N__43722),
            .I(N__43685));
    InMux I__10043 (
            .O(N__43721),
            .I(N__43685));
    InMux I__10042 (
            .O(N__43720),
            .I(N__43685));
    InMux I__10041 (
            .O(N__43719),
            .I(N__43685));
    InMux I__10040 (
            .O(N__43718),
            .I(N__43676));
    InMux I__10039 (
            .O(N__43717),
            .I(N__43676));
    InMux I__10038 (
            .O(N__43716),
            .I(N__43676));
    InMux I__10037 (
            .O(N__43715),
            .I(N__43676));
    InMux I__10036 (
            .O(N__43714),
            .I(N__43667));
    InMux I__10035 (
            .O(N__43713),
            .I(N__43667));
    InMux I__10034 (
            .O(N__43712),
            .I(N__43667));
    InMux I__10033 (
            .O(N__43711),
            .I(N__43667));
    InMux I__10032 (
            .O(N__43710),
            .I(N__43658));
    InMux I__10031 (
            .O(N__43709),
            .I(N__43658));
    InMux I__10030 (
            .O(N__43708),
            .I(N__43658));
    InMux I__10029 (
            .O(N__43707),
            .I(N__43658));
    InMux I__10028 (
            .O(N__43706),
            .I(N__43649));
    InMux I__10027 (
            .O(N__43705),
            .I(N__43649));
    InMux I__10026 (
            .O(N__43704),
            .I(N__43649));
    InMux I__10025 (
            .O(N__43703),
            .I(N__43649));
    LocalMux I__10024 (
            .O(N__43694),
            .I(N__43634));
    LocalMux I__10023 (
            .O(N__43685),
            .I(N__43634));
    LocalMux I__10022 (
            .O(N__43676),
            .I(N__43634));
    LocalMux I__10021 (
            .O(N__43667),
            .I(N__43634));
    LocalMux I__10020 (
            .O(N__43658),
            .I(N__43629));
    LocalMux I__10019 (
            .O(N__43649),
            .I(N__43629));
    InMux I__10018 (
            .O(N__43648),
            .I(N__43624));
    InMux I__10017 (
            .O(N__43647),
            .I(N__43624));
    InMux I__10016 (
            .O(N__43646),
            .I(N__43615));
    InMux I__10015 (
            .O(N__43645),
            .I(N__43615));
    InMux I__10014 (
            .O(N__43644),
            .I(N__43615));
    InMux I__10013 (
            .O(N__43643),
            .I(N__43615));
    Span4Mux_v I__10012 (
            .O(N__43634),
            .I(N__43606));
    Span4Mux_v I__10011 (
            .O(N__43629),
            .I(N__43606));
    LocalMux I__10010 (
            .O(N__43624),
            .I(N__43606));
    LocalMux I__10009 (
            .O(N__43615),
            .I(N__43606));
    Span4Mux_h I__10008 (
            .O(N__43606),
            .I(N__43603));
    Odrv4 I__10007 (
            .O(N__43603),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__10006 (
            .O(N__43600),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CascadeMux I__10005 (
            .O(N__43597),
            .I(N__43594));
    InMux I__10004 (
            .O(N__43594),
            .I(N__43591));
    LocalMux I__10003 (
            .O(N__43591),
            .I(N__43587));
    InMux I__10002 (
            .O(N__43590),
            .I(N__43584));
    Span4Mux_v I__10001 (
            .O(N__43587),
            .I(N__43581));
    LocalMux I__10000 (
            .O(N__43584),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__9999 (
            .O(N__43581),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__9998 (
            .O(N__43576),
            .I(N__43573));
    LocalMux I__9997 (
            .O(N__43573),
            .I(N__43568));
    CEMux I__9996 (
            .O(N__43572),
            .I(N__43565));
    CEMux I__9995 (
            .O(N__43571),
            .I(N__43562));
    Span4Mux_v I__9994 (
            .O(N__43568),
            .I(N__43556));
    LocalMux I__9993 (
            .O(N__43565),
            .I(N__43556));
    LocalMux I__9992 (
            .O(N__43562),
            .I(N__43553));
    CEMux I__9991 (
            .O(N__43561),
            .I(N__43550));
    Span4Mux_v I__9990 (
            .O(N__43556),
            .I(N__43545));
    Span4Mux_v I__9989 (
            .O(N__43553),
            .I(N__43545));
    LocalMux I__9988 (
            .O(N__43550),
            .I(N__43542));
    Span4Mux_h I__9987 (
            .O(N__43545),
            .I(N__43539));
    Span4Mux_h I__9986 (
            .O(N__43542),
            .I(N__43536));
    Odrv4 I__9985 (
            .O(N__43539),
            .I(\current_shift_inst.timer_s1.N_191_i ));
    Odrv4 I__9984 (
            .O(N__43536),
            .I(\current_shift_inst.timer_s1.N_191_i ));
    InMux I__9983 (
            .O(N__43531),
            .I(N__43528));
    LocalMux I__9982 (
            .O(N__43528),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ));
    InMux I__9981 (
            .O(N__43525),
            .I(N__43522));
    LocalMux I__9980 (
            .O(N__43522),
            .I(N__43519));
    Odrv12 I__9979 (
            .O(N__43519),
            .I(\current_shift_inst.un4_control_input_axb_14 ));
    InMux I__9978 (
            .O(N__43516),
            .I(N__43513));
    LocalMux I__9977 (
            .O(N__43513),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ));
    InMux I__9976 (
            .O(N__43510),
            .I(N__43507));
    LocalMux I__9975 (
            .O(N__43507),
            .I(N__43504));
    Odrv12 I__9974 (
            .O(N__43504),
            .I(\current_shift_inst.un4_control_input_axb_24 ));
    InMux I__9973 (
            .O(N__43501),
            .I(N__43490));
    InMux I__9972 (
            .O(N__43500),
            .I(N__43483));
    InMux I__9971 (
            .O(N__43499),
            .I(N__43483));
    InMux I__9970 (
            .O(N__43498),
            .I(N__43483));
    InMux I__9969 (
            .O(N__43497),
            .I(N__43474));
    InMux I__9968 (
            .O(N__43496),
            .I(N__43474));
    InMux I__9967 (
            .O(N__43495),
            .I(N__43474));
    InMux I__9966 (
            .O(N__43494),
            .I(N__43474));
    InMux I__9965 (
            .O(N__43493),
            .I(N__43446));
    LocalMux I__9964 (
            .O(N__43490),
            .I(N__43443));
    LocalMux I__9963 (
            .O(N__43483),
            .I(N__43438));
    LocalMux I__9962 (
            .O(N__43474),
            .I(N__43438));
    InMux I__9961 (
            .O(N__43473),
            .I(N__43435));
    CascadeMux I__9960 (
            .O(N__43472),
            .I(N__43431));
    CascadeMux I__9959 (
            .O(N__43471),
            .I(N__43427));
    CascadeMux I__9958 (
            .O(N__43470),
            .I(N__43424));
    CascadeMux I__9957 (
            .O(N__43469),
            .I(N__43421));
    CascadeMux I__9956 (
            .O(N__43468),
            .I(N__43418));
    CascadeMux I__9955 (
            .O(N__43467),
            .I(N__43415));
    CascadeMux I__9954 (
            .O(N__43466),
            .I(N__43412));
    CascadeMux I__9953 (
            .O(N__43465),
            .I(N__43409));
    CascadeMux I__9952 (
            .O(N__43464),
            .I(N__43406));
    CascadeMux I__9951 (
            .O(N__43463),
            .I(N__43403));
    CascadeMux I__9950 (
            .O(N__43462),
            .I(N__43400));
    CascadeMux I__9949 (
            .O(N__43461),
            .I(N__43397));
    CascadeMux I__9948 (
            .O(N__43460),
            .I(N__43394));
    CascadeMux I__9947 (
            .O(N__43459),
            .I(N__43391));
    CascadeMux I__9946 (
            .O(N__43458),
            .I(N__43388));
    CascadeMux I__9945 (
            .O(N__43457),
            .I(N__43385));
    CascadeMux I__9944 (
            .O(N__43456),
            .I(N__43382));
    CascadeMux I__9943 (
            .O(N__43455),
            .I(N__43379));
    CascadeMux I__9942 (
            .O(N__43454),
            .I(N__43376));
    CascadeMux I__9941 (
            .O(N__43453),
            .I(N__43373));
    CascadeMux I__9940 (
            .O(N__43452),
            .I(N__43370));
    CascadeMux I__9939 (
            .O(N__43451),
            .I(N__43367));
    CascadeMux I__9938 (
            .O(N__43450),
            .I(N__43364));
    InMux I__9937 (
            .O(N__43449),
            .I(N__43354));
    LocalMux I__9936 (
            .O(N__43446),
            .I(N__43351));
    Span4Mux_h I__9935 (
            .O(N__43443),
            .I(N__43345));
    Span4Mux_v I__9934 (
            .O(N__43438),
            .I(N__43345));
    LocalMux I__9933 (
            .O(N__43435),
            .I(N__43342));
    CascadeMux I__9932 (
            .O(N__43434),
            .I(N__43331));
    InMux I__9931 (
            .O(N__43431),
            .I(N__43326));
    InMux I__9930 (
            .O(N__43430),
            .I(N__43326));
    InMux I__9929 (
            .O(N__43427),
            .I(N__43317));
    InMux I__9928 (
            .O(N__43424),
            .I(N__43317));
    InMux I__9927 (
            .O(N__43421),
            .I(N__43317));
    InMux I__9926 (
            .O(N__43418),
            .I(N__43317));
    InMux I__9925 (
            .O(N__43415),
            .I(N__43308));
    InMux I__9924 (
            .O(N__43412),
            .I(N__43308));
    InMux I__9923 (
            .O(N__43409),
            .I(N__43308));
    InMux I__9922 (
            .O(N__43406),
            .I(N__43308));
    InMux I__9921 (
            .O(N__43403),
            .I(N__43301));
    InMux I__9920 (
            .O(N__43400),
            .I(N__43301));
    InMux I__9919 (
            .O(N__43397),
            .I(N__43301));
    InMux I__9918 (
            .O(N__43394),
            .I(N__43294));
    InMux I__9917 (
            .O(N__43391),
            .I(N__43294));
    InMux I__9916 (
            .O(N__43388),
            .I(N__43294));
    InMux I__9915 (
            .O(N__43385),
            .I(N__43285));
    InMux I__9914 (
            .O(N__43382),
            .I(N__43285));
    InMux I__9913 (
            .O(N__43379),
            .I(N__43285));
    InMux I__9912 (
            .O(N__43376),
            .I(N__43285));
    InMux I__9911 (
            .O(N__43373),
            .I(N__43276));
    InMux I__9910 (
            .O(N__43370),
            .I(N__43276));
    InMux I__9909 (
            .O(N__43367),
            .I(N__43276));
    InMux I__9908 (
            .O(N__43364),
            .I(N__43276));
    CascadeMux I__9907 (
            .O(N__43363),
            .I(N__43273));
    CascadeMux I__9906 (
            .O(N__43362),
            .I(N__43270));
    CascadeMux I__9905 (
            .O(N__43361),
            .I(N__43267));
    CascadeMux I__9904 (
            .O(N__43360),
            .I(N__43264));
    CascadeMux I__9903 (
            .O(N__43359),
            .I(N__43261));
    CascadeMux I__9902 (
            .O(N__43358),
            .I(N__43258));
    CascadeMux I__9901 (
            .O(N__43357),
            .I(N__43255));
    LocalMux I__9900 (
            .O(N__43354),
            .I(N__43250));
    Span4Mux_s1_v I__9899 (
            .O(N__43351),
            .I(N__43250));
    InMux I__9898 (
            .O(N__43350),
            .I(N__43247));
    Span4Mux_v I__9897 (
            .O(N__43345),
            .I(N__43242));
    Span4Mux_v I__9896 (
            .O(N__43342),
            .I(N__43242));
    InMux I__9895 (
            .O(N__43341),
            .I(N__43235));
    InMux I__9894 (
            .O(N__43340),
            .I(N__43235));
    InMux I__9893 (
            .O(N__43339),
            .I(N__43235));
    InMux I__9892 (
            .O(N__43338),
            .I(N__43226));
    InMux I__9891 (
            .O(N__43337),
            .I(N__43226));
    InMux I__9890 (
            .O(N__43336),
            .I(N__43226));
    InMux I__9889 (
            .O(N__43335),
            .I(N__43226));
    InMux I__9888 (
            .O(N__43334),
            .I(N__43223));
    InMux I__9887 (
            .O(N__43331),
            .I(N__43220));
    LocalMux I__9886 (
            .O(N__43326),
            .I(N__43217));
    LocalMux I__9885 (
            .O(N__43317),
            .I(N__43212));
    LocalMux I__9884 (
            .O(N__43308),
            .I(N__43212));
    LocalMux I__9883 (
            .O(N__43301),
            .I(N__43203));
    LocalMux I__9882 (
            .O(N__43294),
            .I(N__43203));
    LocalMux I__9881 (
            .O(N__43285),
            .I(N__43203));
    LocalMux I__9880 (
            .O(N__43276),
            .I(N__43203));
    InMux I__9879 (
            .O(N__43273),
            .I(N__43196));
    InMux I__9878 (
            .O(N__43270),
            .I(N__43196));
    InMux I__9877 (
            .O(N__43267),
            .I(N__43196));
    InMux I__9876 (
            .O(N__43264),
            .I(N__43187));
    InMux I__9875 (
            .O(N__43261),
            .I(N__43187));
    InMux I__9874 (
            .O(N__43258),
            .I(N__43187));
    InMux I__9873 (
            .O(N__43255),
            .I(N__43187));
    Sp12to4 I__9872 (
            .O(N__43250),
            .I(N__43182));
    LocalMux I__9871 (
            .O(N__43247),
            .I(N__43182));
    Span4Mux_h I__9870 (
            .O(N__43242),
            .I(N__43179));
    LocalMux I__9869 (
            .O(N__43235),
            .I(N__43174));
    LocalMux I__9868 (
            .O(N__43226),
            .I(N__43174));
    LocalMux I__9867 (
            .O(N__43223),
            .I(N__43171));
    LocalMux I__9866 (
            .O(N__43220),
            .I(N__43166));
    Sp12to4 I__9865 (
            .O(N__43217),
            .I(N__43166));
    Span4Mux_v I__9864 (
            .O(N__43212),
            .I(N__43163));
    Span4Mux_v I__9863 (
            .O(N__43203),
            .I(N__43156));
    LocalMux I__9862 (
            .O(N__43196),
            .I(N__43156));
    LocalMux I__9861 (
            .O(N__43187),
            .I(N__43156));
    Span12Mux_s7_h I__9860 (
            .O(N__43182),
            .I(N__43153));
    Sp12to4 I__9859 (
            .O(N__43179),
            .I(N__43148));
    Span12Mux_s5_h I__9858 (
            .O(N__43174),
            .I(N__43148));
    Span12Mux_s10_h I__9857 (
            .O(N__43171),
            .I(N__43145));
    Span12Mux_v I__9856 (
            .O(N__43166),
            .I(N__43142));
    Span4Mux_h I__9855 (
            .O(N__43163),
            .I(N__43137));
    Span4Mux_h I__9854 (
            .O(N__43156),
            .I(N__43137));
    Span12Mux_v I__9853 (
            .O(N__43153),
            .I(N__43134));
    Span12Mux_h I__9852 (
            .O(N__43148),
            .I(N__43131));
    Span12Mux_v I__9851 (
            .O(N__43145),
            .I(N__43126));
    Span12Mux_h I__9850 (
            .O(N__43142),
            .I(N__43126));
    Span4Mux_v I__9849 (
            .O(N__43137),
            .I(N__43123));
    Odrv12 I__9848 (
            .O(N__43134),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__9847 (
            .O(N__43131),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__9846 (
            .O(N__43126),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__9845 (
            .O(N__43123),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__9844 (
            .O(N__43114),
            .I(N__43110));
    InMux I__9843 (
            .O(N__43113),
            .I(N__43107));
    InMux I__9842 (
            .O(N__43110),
            .I(N__43104));
    LocalMux I__9841 (
            .O(N__43107),
            .I(N__43098));
    LocalMux I__9840 (
            .O(N__43104),
            .I(N__43098));
    InMux I__9839 (
            .O(N__43103),
            .I(N__43095));
    Span4Mux_v I__9838 (
            .O(N__43098),
            .I(N__43092));
    LocalMux I__9837 (
            .O(N__43095),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__9836 (
            .O(N__43092),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__9835 (
            .O(N__43087),
            .I(bfn_17_13_0_));
    CascadeMux I__9834 (
            .O(N__43084),
            .I(N__43080));
    InMux I__9833 (
            .O(N__43083),
            .I(N__43077));
    InMux I__9832 (
            .O(N__43080),
            .I(N__43074));
    LocalMux I__9831 (
            .O(N__43077),
            .I(N__43068));
    LocalMux I__9830 (
            .O(N__43074),
            .I(N__43068));
    InMux I__9829 (
            .O(N__43073),
            .I(N__43065));
    Span4Mux_v I__9828 (
            .O(N__43068),
            .I(N__43062));
    LocalMux I__9827 (
            .O(N__43065),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__9826 (
            .O(N__43062),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__9825 (
            .O(N__43057),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    CascadeMux I__9824 (
            .O(N__43054),
            .I(N__43050));
    CascadeMux I__9823 (
            .O(N__43053),
            .I(N__43047));
    InMux I__9822 (
            .O(N__43050),
            .I(N__43041));
    InMux I__9821 (
            .O(N__43047),
            .I(N__43041));
    InMux I__9820 (
            .O(N__43046),
            .I(N__43038));
    LocalMux I__9819 (
            .O(N__43041),
            .I(N__43035));
    LocalMux I__9818 (
            .O(N__43038),
            .I(N__43030));
    Span4Mux_v I__9817 (
            .O(N__43035),
            .I(N__43030));
    Odrv4 I__9816 (
            .O(N__43030),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__9815 (
            .O(N__43027),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__9814 (
            .O(N__43024),
            .I(N__43020));
    InMux I__9813 (
            .O(N__43023),
            .I(N__43016));
    InMux I__9812 (
            .O(N__43020),
            .I(N__43013));
    InMux I__9811 (
            .O(N__43019),
            .I(N__43010));
    LocalMux I__9810 (
            .O(N__43016),
            .I(N__43005));
    LocalMux I__9809 (
            .O(N__43013),
            .I(N__43005));
    LocalMux I__9808 (
            .O(N__43010),
            .I(N__43000));
    Span4Mux_v I__9807 (
            .O(N__43005),
            .I(N__43000));
    Odrv4 I__9806 (
            .O(N__43000),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__9805 (
            .O(N__42997),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__9804 (
            .O(N__42994),
            .I(N__42988));
    InMux I__9803 (
            .O(N__42993),
            .I(N__42988));
    LocalMux I__9802 (
            .O(N__42988),
            .I(N__42984));
    InMux I__9801 (
            .O(N__42987),
            .I(N__42981));
    Span4Mux_v I__9800 (
            .O(N__42984),
            .I(N__42978));
    LocalMux I__9799 (
            .O(N__42981),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__9798 (
            .O(N__42978),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__9797 (
            .O(N__42973),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__9796 (
            .O(N__42970),
            .I(N__42966));
    CascadeMux I__9795 (
            .O(N__42969),
            .I(N__42963));
    InMux I__9794 (
            .O(N__42966),
            .I(N__42958));
    InMux I__9793 (
            .O(N__42963),
            .I(N__42958));
    LocalMux I__9792 (
            .O(N__42958),
            .I(N__42954));
    InMux I__9791 (
            .O(N__42957),
            .I(N__42951));
    Span4Mux_v I__9790 (
            .O(N__42954),
            .I(N__42948));
    LocalMux I__9789 (
            .O(N__42951),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__9788 (
            .O(N__42948),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__9787 (
            .O(N__42943),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__9786 (
            .O(N__42940),
            .I(N__42936));
    InMux I__9785 (
            .O(N__42939),
            .I(N__42933));
    InMux I__9784 (
            .O(N__42936),
            .I(N__42930));
    LocalMux I__9783 (
            .O(N__42933),
            .I(N__42924));
    LocalMux I__9782 (
            .O(N__42930),
            .I(N__42924));
    InMux I__9781 (
            .O(N__42929),
            .I(N__42921));
    Span4Mux_v I__9780 (
            .O(N__42924),
            .I(N__42918));
    LocalMux I__9779 (
            .O(N__42921),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__9778 (
            .O(N__42918),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__9777 (
            .O(N__42913),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__9776 (
            .O(N__42910),
            .I(N__42904));
    InMux I__9775 (
            .O(N__42909),
            .I(N__42904));
    LocalMux I__9774 (
            .O(N__42904),
            .I(N__42900));
    InMux I__9773 (
            .O(N__42903),
            .I(N__42897));
    Span4Mux_v I__9772 (
            .O(N__42900),
            .I(N__42894));
    LocalMux I__9771 (
            .O(N__42897),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__9770 (
            .O(N__42894),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__9769 (
            .O(N__42889),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    CascadeMux I__9768 (
            .O(N__42886),
            .I(N__42882));
    InMux I__9767 (
            .O(N__42885),
            .I(N__42879));
    InMux I__9766 (
            .O(N__42882),
            .I(N__42876));
    LocalMux I__9765 (
            .O(N__42879),
            .I(N__42870));
    LocalMux I__9764 (
            .O(N__42876),
            .I(N__42870));
    InMux I__9763 (
            .O(N__42875),
            .I(N__42867));
    Span4Mux_v I__9762 (
            .O(N__42870),
            .I(N__42864));
    LocalMux I__9761 (
            .O(N__42867),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__9760 (
            .O(N__42864),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    CascadeMux I__9759 (
            .O(N__42859),
            .I(N__42855));
    InMux I__9758 (
            .O(N__42858),
            .I(N__42852));
    InMux I__9757 (
            .O(N__42855),
            .I(N__42849));
    LocalMux I__9756 (
            .O(N__42852),
            .I(N__42843));
    LocalMux I__9755 (
            .O(N__42849),
            .I(N__42843));
    InMux I__9754 (
            .O(N__42848),
            .I(N__42840));
    Span4Mux_v I__9753 (
            .O(N__42843),
            .I(N__42837));
    LocalMux I__9752 (
            .O(N__42840),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__9751 (
            .O(N__42837),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__9750 (
            .O(N__42832),
            .I(bfn_17_12_0_));
    CascadeMux I__9749 (
            .O(N__42829),
            .I(N__42825));
    CascadeMux I__9748 (
            .O(N__42828),
            .I(N__42822));
    InMux I__9747 (
            .O(N__42825),
            .I(N__42819));
    InMux I__9746 (
            .O(N__42822),
            .I(N__42816));
    LocalMux I__9745 (
            .O(N__42819),
            .I(N__42810));
    LocalMux I__9744 (
            .O(N__42816),
            .I(N__42810));
    InMux I__9743 (
            .O(N__42815),
            .I(N__42807));
    Span4Mux_v I__9742 (
            .O(N__42810),
            .I(N__42804));
    LocalMux I__9741 (
            .O(N__42807),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__9740 (
            .O(N__42804),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__9739 (
            .O(N__42799),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__9738 (
            .O(N__42796),
            .I(N__42792));
    InMux I__9737 (
            .O(N__42795),
            .I(N__42788));
    InMux I__9736 (
            .O(N__42792),
            .I(N__42785));
    InMux I__9735 (
            .O(N__42791),
            .I(N__42782));
    LocalMux I__9734 (
            .O(N__42788),
            .I(N__42777));
    LocalMux I__9733 (
            .O(N__42785),
            .I(N__42777));
    LocalMux I__9732 (
            .O(N__42782),
            .I(N__42772));
    Span4Mux_v I__9731 (
            .O(N__42777),
            .I(N__42772));
    Odrv4 I__9730 (
            .O(N__42772),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__9729 (
            .O(N__42769),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__9728 (
            .O(N__42766),
            .I(N__42759));
    InMux I__9727 (
            .O(N__42765),
            .I(N__42759));
    InMux I__9726 (
            .O(N__42764),
            .I(N__42756));
    LocalMux I__9725 (
            .O(N__42759),
            .I(N__42753));
    LocalMux I__9724 (
            .O(N__42756),
            .I(N__42748));
    Span4Mux_v I__9723 (
            .O(N__42753),
            .I(N__42748));
    Odrv4 I__9722 (
            .O(N__42748),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__9721 (
            .O(N__42745),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    CascadeMux I__9720 (
            .O(N__42742),
            .I(N__42738));
    CascadeMux I__9719 (
            .O(N__42741),
            .I(N__42735));
    InMux I__9718 (
            .O(N__42738),
            .I(N__42730));
    InMux I__9717 (
            .O(N__42735),
            .I(N__42730));
    LocalMux I__9716 (
            .O(N__42730),
            .I(N__42726));
    InMux I__9715 (
            .O(N__42729),
            .I(N__42723));
    Span4Mux_v I__9714 (
            .O(N__42726),
            .I(N__42720));
    LocalMux I__9713 (
            .O(N__42723),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__9712 (
            .O(N__42720),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__9711 (
            .O(N__42715),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__9710 (
            .O(N__42712),
            .I(N__42708));
    CascadeMux I__9709 (
            .O(N__42711),
            .I(N__42705));
    InMux I__9708 (
            .O(N__42708),
            .I(N__42700));
    InMux I__9707 (
            .O(N__42705),
            .I(N__42700));
    LocalMux I__9706 (
            .O(N__42700),
            .I(N__42696));
    InMux I__9705 (
            .O(N__42699),
            .I(N__42693));
    Span4Mux_v I__9704 (
            .O(N__42696),
            .I(N__42690));
    LocalMux I__9703 (
            .O(N__42693),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__9702 (
            .O(N__42690),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__9701 (
            .O(N__42685),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__9700 (
            .O(N__42682),
            .I(N__42676));
    InMux I__9699 (
            .O(N__42681),
            .I(N__42676));
    LocalMux I__9698 (
            .O(N__42676),
            .I(N__42672));
    InMux I__9697 (
            .O(N__42675),
            .I(N__42669));
    Span4Mux_v I__9696 (
            .O(N__42672),
            .I(N__42666));
    LocalMux I__9695 (
            .O(N__42669),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__9694 (
            .O(N__42666),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__9693 (
            .O(N__42661),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__9692 (
            .O(N__42658),
            .I(N__42652));
    InMux I__9691 (
            .O(N__42657),
            .I(N__42652));
    LocalMux I__9690 (
            .O(N__42652),
            .I(N__42648));
    InMux I__9689 (
            .O(N__42651),
            .I(N__42645));
    Span4Mux_v I__9688 (
            .O(N__42648),
            .I(N__42642));
    LocalMux I__9687 (
            .O(N__42645),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__9686 (
            .O(N__42642),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__9685 (
            .O(N__42637),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__9684 (
            .O(N__42634),
            .I(N__42631));
    InMux I__9683 (
            .O(N__42631),
            .I(N__42623));
    InMux I__9682 (
            .O(N__42630),
            .I(N__42623));
    InMux I__9681 (
            .O(N__42629),
            .I(N__42618));
    InMux I__9680 (
            .O(N__42628),
            .I(N__42618));
    LocalMux I__9679 (
            .O(N__42623),
            .I(N__42615));
    LocalMux I__9678 (
            .O(N__42618),
            .I(N__42612));
    Span4Mux_v I__9677 (
            .O(N__42615),
            .I(N__42609));
    Span4Mux_v I__9676 (
            .O(N__42612),
            .I(N__42606));
    Odrv4 I__9675 (
            .O(N__42609),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    Odrv4 I__9674 (
            .O(N__42606),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    InMux I__9673 (
            .O(N__42601),
            .I(N__42595));
    InMux I__9672 (
            .O(N__42600),
            .I(N__42595));
    LocalMux I__9671 (
            .O(N__42595),
            .I(N__42592));
    Span4Mux_v I__9670 (
            .O(N__42592),
            .I(N__42585));
    InMux I__9669 (
            .O(N__42591),
            .I(N__42580));
    InMux I__9668 (
            .O(N__42590),
            .I(N__42580));
    InMux I__9667 (
            .O(N__42589),
            .I(N__42575));
    InMux I__9666 (
            .O(N__42588),
            .I(N__42575));
    Odrv4 I__9665 (
            .O(N__42585),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__9664 (
            .O(N__42580),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__9663 (
            .O(N__42575),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__9662 (
            .O(N__42568),
            .I(N__42564));
    CascadeMux I__9661 (
            .O(N__42567),
            .I(N__42561));
    LocalMux I__9660 (
            .O(N__42564),
            .I(N__42558));
    InMux I__9659 (
            .O(N__42561),
            .I(N__42555));
    Span4Mux_h I__9658 (
            .O(N__42558),
            .I(N__42549));
    LocalMux I__9657 (
            .O(N__42555),
            .I(N__42549));
    InMux I__9656 (
            .O(N__42554),
            .I(N__42546));
    Span4Mux_v I__9655 (
            .O(N__42549),
            .I(N__42543));
    LocalMux I__9654 (
            .O(N__42546),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__9653 (
            .O(N__42543),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__9652 (
            .O(N__42538),
            .I(bfn_17_11_0_));
    InMux I__9651 (
            .O(N__42535),
            .I(N__42532));
    LocalMux I__9650 (
            .O(N__42532),
            .I(N__42528));
    CascadeMux I__9649 (
            .O(N__42531),
            .I(N__42525));
    Span4Mux_h I__9648 (
            .O(N__42528),
            .I(N__42522));
    InMux I__9647 (
            .O(N__42525),
            .I(N__42519));
    Span4Mux_h I__9646 (
            .O(N__42522),
            .I(N__42513));
    LocalMux I__9645 (
            .O(N__42519),
            .I(N__42513));
    InMux I__9644 (
            .O(N__42518),
            .I(N__42510));
    Span4Mux_v I__9643 (
            .O(N__42513),
            .I(N__42507));
    LocalMux I__9642 (
            .O(N__42510),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__9641 (
            .O(N__42507),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__9640 (
            .O(N__42502),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__9639 (
            .O(N__42499),
            .I(N__42492));
    InMux I__9638 (
            .O(N__42498),
            .I(N__42492));
    InMux I__9637 (
            .O(N__42497),
            .I(N__42489));
    LocalMux I__9636 (
            .O(N__42492),
            .I(N__42486));
    LocalMux I__9635 (
            .O(N__42489),
            .I(N__42481));
    Span4Mux_v I__9634 (
            .O(N__42486),
            .I(N__42481));
    Odrv4 I__9633 (
            .O(N__42481),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__9632 (
            .O(N__42478),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__9631 (
            .O(N__42475),
            .I(N__42469));
    InMux I__9630 (
            .O(N__42474),
            .I(N__42469));
    LocalMux I__9629 (
            .O(N__42469),
            .I(N__42465));
    InMux I__9628 (
            .O(N__42468),
            .I(N__42462));
    Sp12to4 I__9627 (
            .O(N__42465),
            .I(N__42459));
    LocalMux I__9626 (
            .O(N__42462),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv12 I__9625 (
            .O(N__42459),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__9624 (
            .O(N__42454),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__9623 (
            .O(N__42451),
            .I(N__42447));
    CascadeMux I__9622 (
            .O(N__42450),
            .I(N__42444));
    InMux I__9621 (
            .O(N__42447),
            .I(N__42439));
    InMux I__9620 (
            .O(N__42444),
            .I(N__42439));
    LocalMux I__9619 (
            .O(N__42439),
            .I(N__42435));
    InMux I__9618 (
            .O(N__42438),
            .I(N__42432));
    Span4Mux_v I__9617 (
            .O(N__42435),
            .I(N__42429));
    LocalMux I__9616 (
            .O(N__42432),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__9615 (
            .O(N__42429),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__9614 (
            .O(N__42424),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__9613 (
            .O(N__42421),
            .I(N__42417));
    CascadeMux I__9612 (
            .O(N__42420),
            .I(N__42414));
    InMux I__9611 (
            .O(N__42417),
            .I(N__42409));
    InMux I__9610 (
            .O(N__42414),
            .I(N__42409));
    LocalMux I__9609 (
            .O(N__42409),
            .I(N__42405));
    InMux I__9608 (
            .O(N__42408),
            .I(N__42402));
    Span4Mux_v I__9607 (
            .O(N__42405),
            .I(N__42399));
    LocalMux I__9606 (
            .O(N__42402),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__9605 (
            .O(N__42399),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__9604 (
            .O(N__42394),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__9603 (
            .O(N__42391),
            .I(N__42385));
    InMux I__9602 (
            .O(N__42390),
            .I(N__42385));
    LocalMux I__9601 (
            .O(N__42385),
            .I(N__42381));
    InMux I__9600 (
            .O(N__42384),
            .I(N__42378));
    Span4Mux_v I__9599 (
            .O(N__42381),
            .I(N__42375));
    LocalMux I__9598 (
            .O(N__42378),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__9597 (
            .O(N__42375),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__9596 (
            .O(N__42370),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__9595 (
            .O(N__42367),
            .I(N__42361));
    InMux I__9594 (
            .O(N__42366),
            .I(N__42361));
    LocalMux I__9593 (
            .O(N__42361),
            .I(N__42357));
    InMux I__9592 (
            .O(N__42360),
            .I(N__42354));
    Span4Mux_v I__9591 (
            .O(N__42357),
            .I(N__42351));
    LocalMux I__9590 (
            .O(N__42354),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__9589 (
            .O(N__42351),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__9588 (
            .O(N__42346),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    InMux I__9587 (
            .O(N__42343),
            .I(N__42340));
    LocalMux I__9586 (
            .O(N__42340),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__9585 (
            .O(N__42337),
            .I(\phase_controller_slave.N_214_cascade_ ));
    CascadeMux I__9584 (
            .O(N__42334),
            .I(N__42328));
    CascadeMux I__9583 (
            .O(N__42333),
            .I(N__42325));
    CascadeMux I__9582 (
            .O(N__42332),
            .I(N__42322));
    CascadeMux I__9581 (
            .O(N__42331),
            .I(N__42319));
    InMux I__9580 (
            .O(N__42328),
            .I(N__42296));
    InMux I__9579 (
            .O(N__42325),
            .I(N__42296));
    InMux I__9578 (
            .O(N__42322),
            .I(N__42296));
    InMux I__9577 (
            .O(N__42319),
            .I(N__42296));
    InMux I__9576 (
            .O(N__42318),
            .I(N__42287));
    InMux I__9575 (
            .O(N__42317),
            .I(N__42287));
    InMux I__9574 (
            .O(N__42316),
            .I(N__42287));
    InMux I__9573 (
            .O(N__42315),
            .I(N__42287));
    InMux I__9572 (
            .O(N__42314),
            .I(N__42272));
    InMux I__9571 (
            .O(N__42313),
            .I(N__42272));
    InMux I__9570 (
            .O(N__42312),
            .I(N__42272));
    InMux I__9569 (
            .O(N__42311),
            .I(N__42272));
    InMux I__9568 (
            .O(N__42310),
            .I(N__42272));
    InMux I__9567 (
            .O(N__42309),
            .I(N__42272));
    InMux I__9566 (
            .O(N__42308),
            .I(N__42272));
    CascadeMux I__9565 (
            .O(N__42307),
            .I(N__42267));
    CascadeMux I__9564 (
            .O(N__42306),
            .I(N__42264));
    InMux I__9563 (
            .O(N__42305),
            .I(N__42261));
    LocalMux I__9562 (
            .O(N__42296),
            .I(N__42254));
    LocalMux I__9561 (
            .O(N__42287),
            .I(N__42254));
    LocalMux I__9560 (
            .O(N__42272),
            .I(N__42254));
    CascadeMux I__9559 (
            .O(N__42271),
            .I(N__42251));
    InMux I__9558 (
            .O(N__42270),
            .I(N__42247));
    InMux I__9557 (
            .O(N__42267),
            .I(N__42242));
    InMux I__9556 (
            .O(N__42264),
            .I(N__42242));
    LocalMux I__9555 (
            .O(N__42261),
            .I(N__42237));
    Span4Mux_v I__9554 (
            .O(N__42254),
            .I(N__42237));
    InMux I__9553 (
            .O(N__42251),
            .I(N__42232));
    InMux I__9552 (
            .O(N__42250),
            .I(N__42232));
    LocalMux I__9551 (
            .O(N__42247),
            .I(N__42227));
    LocalMux I__9550 (
            .O(N__42242),
            .I(N__42220));
    Span4Mux_h I__9549 (
            .O(N__42237),
            .I(N__42220));
    LocalMux I__9548 (
            .O(N__42232),
            .I(N__42220));
    InMux I__9547 (
            .O(N__42231),
            .I(N__42214));
    InMux I__9546 (
            .O(N__42230),
            .I(N__42214));
    Span4Mux_v I__9545 (
            .O(N__42227),
            .I(N__42211));
    Span4Mux_h I__9544 (
            .O(N__42220),
            .I(N__42208));
    InMux I__9543 (
            .O(N__42219),
            .I(N__42205));
    LocalMux I__9542 (
            .O(N__42214),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__9541 (
            .O(N__42211),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__9540 (
            .O(N__42208),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__9539 (
            .O(N__42205),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__9538 (
            .O(N__42196),
            .I(N__42192));
    CascadeMux I__9537 (
            .O(N__42195),
            .I(N__42184));
    InMux I__9536 (
            .O(N__42192),
            .I(N__42179));
    InMux I__9535 (
            .O(N__42191),
            .I(N__42179));
    CascadeMux I__9534 (
            .O(N__42190),
            .I(N__42169));
    CascadeMux I__9533 (
            .O(N__42189),
            .I(N__42166));
    CascadeMux I__9532 (
            .O(N__42188),
            .I(N__42163));
    CascadeMux I__9531 (
            .O(N__42187),
            .I(N__42160));
    InMux I__9530 (
            .O(N__42184),
            .I(N__42157));
    LocalMux I__9529 (
            .O(N__42179),
            .I(N__42154));
    CascadeMux I__9528 (
            .O(N__42178),
            .I(N__42147));
    CascadeMux I__9527 (
            .O(N__42177),
            .I(N__42144));
    CascadeMux I__9526 (
            .O(N__42176),
            .I(N__42141));
    CascadeMux I__9525 (
            .O(N__42175),
            .I(N__42138));
    InMux I__9524 (
            .O(N__42174),
            .I(N__42117));
    InMux I__9523 (
            .O(N__42173),
            .I(N__42117));
    InMux I__9522 (
            .O(N__42172),
            .I(N__42117));
    InMux I__9521 (
            .O(N__42169),
            .I(N__42117));
    InMux I__9520 (
            .O(N__42166),
            .I(N__42117));
    InMux I__9519 (
            .O(N__42163),
            .I(N__42117));
    InMux I__9518 (
            .O(N__42160),
            .I(N__42117));
    LocalMux I__9517 (
            .O(N__42157),
            .I(N__42114));
    Span4Mux_h I__9516 (
            .O(N__42154),
            .I(N__42111));
    InMux I__9515 (
            .O(N__42153),
            .I(N__42102));
    InMux I__9514 (
            .O(N__42152),
            .I(N__42102));
    InMux I__9513 (
            .O(N__42151),
            .I(N__42102));
    InMux I__9512 (
            .O(N__42150),
            .I(N__42102));
    InMux I__9511 (
            .O(N__42147),
            .I(N__42085));
    InMux I__9510 (
            .O(N__42144),
            .I(N__42085));
    InMux I__9509 (
            .O(N__42141),
            .I(N__42085));
    InMux I__9508 (
            .O(N__42138),
            .I(N__42085));
    InMux I__9507 (
            .O(N__42137),
            .I(N__42085));
    InMux I__9506 (
            .O(N__42136),
            .I(N__42085));
    InMux I__9505 (
            .O(N__42135),
            .I(N__42085));
    InMux I__9504 (
            .O(N__42134),
            .I(N__42085));
    InMux I__9503 (
            .O(N__42133),
            .I(N__42080));
    InMux I__9502 (
            .O(N__42132),
            .I(N__42080));
    LocalMux I__9501 (
            .O(N__42117),
            .I(N__42077));
    Span4Mux_v I__9500 (
            .O(N__42114),
            .I(N__42070));
    Span4Mux_v I__9499 (
            .O(N__42111),
            .I(N__42070));
    LocalMux I__9498 (
            .O(N__42102),
            .I(N__42070));
    LocalMux I__9497 (
            .O(N__42085),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    LocalMux I__9496 (
            .O(N__42080),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__9495 (
            .O(N__42077),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__9494 (
            .O(N__42070),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    CascadeMux I__9493 (
            .O(N__42061),
            .I(N__42058));
    InMux I__9492 (
            .O(N__42058),
            .I(N__42039));
    InMux I__9491 (
            .O(N__42057),
            .I(N__42024));
    InMux I__9490 (
            .O(N__42056),
            .I(N__42024));
    InMux I__9489 (
            .O(N__42055),
            .I(N__42024));
    InMux I__9488 (
            .O(N__42054),
            .I(N__42024));
    InMux I__9487 (
            .O(N__42053),
            .I(N__42024));
    InMux I__9486 (
            .O(N__42052),
            .I(N__42024));
    InMux I__9485 (
            .O(N__42051),
            .I(N__42024));
    InMux I__9484 (
            .O(N__42050),
            .I(N__42007));
    InMux I__9483 (
            .O(N__42049),
            .I(N__42007));
    InMux I__9482 (
            .O(N__42048),
            .I(N__42007));
    InMux I__9481 (
            .O(N__42047),
            .I(N__42007));
    InMux I__9480 (
            .O(N__42046),
            .I(N__42007));
    InMux I__9479 (
            .O(N__42045),
            .I(N__42007));
    InMux I__9478 (
            .O(N__42044),
            .I(N__42007));
    InMux I__9477 (
            .O(N__42043),
            .I(N__42007));
    InMux I__9476 (
            .O(N__42042),
            .I(N__41999));
    LocalMux I__9475 (
            .O(N__42039),
            .I(N__41994));
    LocalMux I__9474 (
            .O(N__42024),
            .I(N__41994));
    LocalMux I__9473 (
            .O(N__42007),
            .I(N__41991));
    InMux I__9472 (
            .O(N__42006),
            .I(N__41982));
    InMux I__9471 (
            .O(N__42005),
            .I(N__41982));
    InMux I__9470 (
            .O(N__42004),
            .I(N__41982));
    InMux I__9469 (
            .O(N__42003),
            .I(N__41982));
    CascadeMux I__9468 (
            .O(N__42002),
            .I(N__41979));
    LocalMux I__9467 (
            .O(N__41999),
            .I(N__41975));
    Span4Mux_v I__9466 (
            .O(N__41994),
            .I(N__41968));
    Span4Mux_v I__9465 (
            .O(N__41991),
            .I(N__41968));
    LocalMux I__9464 (
            .O(N__41982),
            .I(N__41968));
    InMux I__9463 (
            .O(N__41979),
            .I(N__41962));
    InMux I__9462 (
            .O(N__41978),
            .I(N__41962));
    Span4Mux_v I__9461 (
            .O(N__41975),
            .I(N__41959));
    Span4Mux_h I__9460 (
            .O(N__41968),
            .I(N__41956));
    InMux I__9459 (
            .O(N__41967),
            .I(N__41953));
    LocalMux I__9458 (
            .O(N__41962),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__9457 (
            .O(N__41959),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__9456 (
            .O(N__41956),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__9455 (
            .O(N__41953),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__9454 (
            .O(N__41944),
            .I(N__41941));
    InMux I__9453 (
            .O(N__41941),
            .I(N__41938));
    LocalMux I__9452 (
            .O(N__41938),
            .I(N__41935));
    Odrv4 I__9451 (
            .O(N__41935),
            .I(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ));
    CascadeMux I__9450 (
            .O(N__41932),
            .I(N__41928));
    InMux I__9449 (
            .O(N__41931),
            .I(N__41924));
    InMux I__9448 (
            .O(N__41928),
            .I(N__41921));
    InMux I__9447 (
            .O(N__41927),
            .I(N__41918));
    LocalMux I__9446 (
            .O(N__41924),
            .I(N__41913));
    LocalMux I__9445 (
            .O(N__41921),
            .I(N__41913));
    LocalMux I__9444 (
            .O(N__41918),
            .I(\current_shift_inst.timer_phase.counterZ0Z_27 ));
    Odrv4 I__9443 (
            .O(N__41913),
            .I(\current_shift_inst.timer_phase.counterZ0Z_27 ));
    CascadeMux I__9442 (
            .O(N__41908),
            .I(N__41905));
    InMux I__9441 (
            .O(N__41905),
            .I(N__41901));
    InMux I__9440 (
            .O(N__41904),
            .I(N__41898));
    LocalMux I__9439 (
            .O(N__41901),
            .I(N__41895));
    LocalMux I__9438 (
            .O(N__41898),
            .I(\current_shift_inst.timer_phase.counterZ0Z_29 ));
    Odrv4 I__9437 (
            .O(N__41895),
            .I(\current_shift_inst.timer_phase.counterZ0Z_29 ));
    InMux I__9436 (
            .O(N__41890),
            .I(N__41887));
    LocalMux I__9435 (
            .O(N__41887),
            .I(N__41883));
    InMux I__9434 (
            .O(N__41886),
            .I(N__41880));
    Span4Mux_h I__9433 (
            .O(N__41883),
            .I(N__41877));
    LocalMux I__9432 (
            .O(N__41880),
            .I(N__41874));
    Span4Mux_v I__9431 (
            .O(N__41877),
            .I(N__41870));
    Span12Mux_h I__9430 (
            .O(N__41874),
            .I(N__41867));
    InMux I__9429 (
            .O(N__41873),
            .I(N__41864));
    Odrv4 I__9428 (
            .O(N__41870),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    Odrv12 I__9427 (
            .O(N__41867),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    LocalMux I__9426 (
            .O(N__41864),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    InMux I__9425 (
            .O(N__41857),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ));
    InMux I__9424 (
            .O(N__41854),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__9423 (
            .O(N__41851),
            .I(N__41848));
    InMux I__9422 (
            .O(N__41848),
            .I(N__41844));
    CascadeMux I__9421 (
            .O(N__41847),
            .I(N__41841));
    LocalMux I__9420 (
            .O(N__41844),
            .I(N__41838));
    InMux I__9419 (
            .O(N__41841),
            .I(N__41835));
    Span4Mux_h I__9418 (
            .O(N__41838),
            .I(N__41832));
    LocalMux I__9417 (
            .O(N__41835),
            .I(N__41829));
    Span4Mux_v I__9416 (
            .O(N__41832),
            .I(N__41824));
    Span4Mux_h I__9415 (
            .O(N__41829),
            .I(N__41824));
    Odrv4 I__9414 (
            .O(N__41824),
            .I(\current_shift_inst.elapsed_time_ns_phase_31 ));
    CEMux I__9413 (
            .O(N__41821),
            .I(N__41806));
    CEMux I__9412 (
            .O(N__41820),
            .I(N__41806));
    CEMux I__9411 (
            .O(N__41819),
            .I(N__41806));
    CEMux I__9410 (
            .O(N__41818),
            .I(N__41806));
    CEMux I__9409 (
            .O(N__41817),
            .I(N__41806));
    GlobalMux I__9408 (
            .O(N__41806),
            .I(N__41803));
    gio2CtrlBuf I__9407 (
            .O(N__41803),
            .I(\current_shift_inst.timer_phase.N_188_i_g ));
    CascadeMux I__9406 (
            .O(N__41800),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_ ));
    InMux I__9405 (
            .O(N__41797),
            .I(N__41794));
    LocalMux I__9404 (
            .O(N__41794),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19 ));
    InMux I__9403 (
            .O(N__41791),
            .I(N__41788));
    LocalMux I__9402 (
            .O(N__41788),
            .I(N__41785));
    Odrv4 I__9401 (
            .O(N__41785),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19 ));
    InMux I__9400 (
            .O(N__41782),
            .I(N__41779));
    LocalMux I__9399 (
            .O(N__41779),
            .I(N__41776));
    Span4Mux_h I__9398 (
            .O(N__41776),
            .I(N__41773));
    Span4Mux_h I__9397 (
            .O(N__41773),
            .I(N__41770));
    Odrv4 I__9396 (
            .O(N__41770),
            .I(il_max_comp2_D1));
    InMux I__9395 (
            .O(N__41767),
            .I(N__41764));
    LocalMux I__9394 (
            .O(N__41764),
            .I(N__41761));
    Span4Mux_h I__9393 (
            .O(N__41761),
            .I(N__41758));
    Span4Mux_h I__9392 (
            .O(N__41758),
            .I(N__41755));
    Odrv4 I__9391 (
            .O(N__41755),
            .I(il_min_comp2_D1));
    CascadeMux I__9390 (
            .O(N__41752),
            .I(N__41747));
    InMux I__9389 (
            .O(N__41751),
            .I(N__41744));
    InMux I__9388 (
            .O(N__41750),
            .I(N__41741));
    InMux I__9387 (
            .O(N__41747),
            .I(N__41738));
    LocalMux I__9386 (
            .O(N__41744),
            .I(N__41731));
    LocalMux I__9385 (
            .O(N__41741),
            .I(N__41731));
    LocalMux I__9384 (
            .O(N__41738),
            .I(N__41731));
    Odrv4 I__9383 (
            .O(N__41731),
            .I(\current_shift_inst.timer_phase.counterZ0Z_19 ));
    InMux I__9382 (
            .O(N__41728),
            .I(N__41722));
    InMux I__9381 (
            .O(N__41727),
            .I(N__41722));
    LocalMux I__9380 (
            .O(N__41722),
            .I(N__41718));
    InMux I__9379 (
            .O(N__41721),
            .I(N__41715));
    Span4Mux_h I__9378 (
            .O(N__41718),
            .I(N__41712));
    LocalMux I__9377 (
            .O(N__41715),
            .I(N__41709));
    Span4Mux_v I__9376 (
            .O(N__41712),
            .I(N__41706));
    Span12Mux_v I__9375 (
            .O(N__41709),
            .I(N__41702));
    Span4Mux_h I__9374 (
            .O(N__41706),
            .I(N__41699));
    InMux I__9373 (
            .O(N__41705),
            .I(N__41696));
    Odrv12 I__9372 (
            .O(N__41702),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    Odrv4 I__9371 (
            .O(N__41699),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    LocalMux I__9370 (
            .O(N__41696),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    InMux I__9369 (
            .O(N__41689),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__9368 (
            .O(N__41686),
            .I(N__41682));
    CascadeMux I__9367 (
            .O(N__41685),
            .I(N__41679));
    InMux I__9366 (
            .O(N__41682),
            .I(N__41673));
    InMux I__9365 (
            .O(N__41679),
            .I(N__41673));
    InMux I__9364 (
            .O(N__41678),
            .I(N__41670));
    LocalMux I__9363 (
            .O(N__41673),
            .I(N__41667));
    LocalMux I__9362 (
            .O(N__41670),
            .I(\current_shift_inst.timer_phase.counterZ0Z_20 ));
    Odrv4 I__9361 (
            .O(N__41667),
            .I(\current_shift_inst.timer_phase.counterZ0Z_20 ));
    InMux I__9360 (
            .O(N__41662),
            .I(N__41658));
    CascadeMux I__9359 (
            .O(N__41661),
            .I(N__41655));
    LocalMux I__9358 (
            .O(N__41658),
            .I(N__41651));
    InMux I__9357 (
            .O(N__41655),
            .I(N__41648));
    InMux I__9356 (
            .O(N__41654),
            .I(N__41645));
    Span4Mux_h I__9355 (
            .O(N__41651),
            .I(N__41642));
    LocalMux I__9354 (
            .O(N__41648),
            .I(N__41639));
    LocalMux I__9353 (
            .O(N__41645),
            .I(N__41635));
    Span4Mux_v I__9352 (
            .O(N__41642),
            .I(N__41632));
    Span12Mux_h I__9351 (
            .O(N__41639),
            .I(N__41629));
    InMux I__9350 (
            .O(N__41638),
            .I(N__41626));
    Odrv12 I__9349 (
            .O(N__41635),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    Odrv4 I__9348 (
            .O(N__41632),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    Odrv12 I__9347 (
            .O(N__41629),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    LocalMux I__9346 (
            .O(N__41626),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    InMux I__9345 (
            .O(N__41617),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__9344 (
            .O(N__41614),
            .I(N__41610));
    CascadeMux I__9343 (
            .O(N__41613),
            .I(N__41607));
    InMux I__9342 (
            .O(N__41610),
            .I(N__41601));
    InMux I__9341 (
            .O(N__41607),
            .I(N__41601));
    InMux I__9340 (
            .O(N__41606),
            .I(N__41598));
    LocalMux I__9339 (
            .O(N__41601),
            .I(N__41595));
    LocalMux I__9338 (
            .O(N__41598),
            .I(\current_shift_inst.timer_phase.counterZ0Z_21 ));
    Odrv4 I__9337 (
            .O(N__41595),
            .I(\current_shift_inst.timer_phase.counterZ0Z_21 ));
    CascadeMux I__9336 (
            .O(N__41590),
            .I(N__41587));
    InMux I__9335 (
            .O(N__41587),
            .I(N__41584));
    LocalMux I__9334 (
            .O(N__41584),
            .I(N__41581));
    Span4Mux_h I__9333 (
            .O(N__41581),
            .I(N__41576));
    InMux I__9332 (
            .O(N__41580),
            .I(N__41571));
    InMux I__9331 (
            .O(N__41579),
            .I(N__41571));
    Span4Mux_v I__9330 (
            .O(N__41576),
            .I(N__41567));
    LocalMux I__9329 (
            .O(N__41571),
            .I(N__41564));
    InMux I__9328 (
            .O(N__41570),
            .I(N__41561));
    Odrv4 I__9327 (
            .O(N__41567),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    Odrv12 I__9326 (
            .O(N__41564),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    LocalMux I__9325 (
            .O(N__41561),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    InMux I__9324 (
            .O(N__41554),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__9323 (
            .O(N__41551),
            .I(N__41548));
    InMux I__9322 (
            .O(N__41548),
            .I(N__41543));
    InMux I__9321 (
            .O(N__41547),
            .I(N__41540));
    InMux I__9320 (
            .O(N__41546),
            .I(N__41537));
    LocalMux I__9319 (
            .O(N__41543),
            .I(N__41532));
    LocalMux I__9318 (
            .O(N__41540),
            .I(N__41532));
    LocalMux I__9317 (
            .O(N__41537),
            .I(\current_shift_inst.timer_phase.counterZ0Z_22 ));
    Odrv12 I__9316 (
            .O(N__41532),
            .I(\current_shift_inst.timer_phase.counterZ0Z_22 ));
    InMux I__9315 (
            .O(N__41527),
            .I(N__41521));
    InMux I__9314 (
            .O(N__41526),
            .I(N__41521));
    LocalMux I__9313 (
            .O(N__41521),
            .I(N__41517));
    InMux I__9312 (
            .O(N__41520),
            .I(N__41514));
    Span4Mux_h I__9311 (
            .O(N__41517),
            .I(N__41511));
    LocalMux I__9310 (
            .O(N__41514),
            .I(N__41507));
    Span4Mux_v I__9309 (
            .O(N__41511),
            .I(N__41504));
    InMux I__9308 (
            .O(N__41510),
            .I(N__41501));
    Odrv12 I__9307 (
            .O(N__41507),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    Odrv4 I__9306 (
            .O(N__41504),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    LocalMux I__9305 (
            .O(N__41501),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    InMux I__9304 (
            .O(N__41494),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ));
    InMux I__9303 (
            .O(N__41491),
            .I(N__41485));
    InMux I__9302 (
            .O(N__41490),
            .I(N__41485));
    LocalMux I__9301 (
            .O(N__41485),
            .I(N__41481));
    InMux I__9300 (
            .O(N__41484),
            .I(N__41478));
    Span4Mux_h I__9299 (
            .O(N__41481),
            .I(N__41475));
    LocalMux I__9298 (
            .O(N__41478),
            .I(\current_shift_inst.timer_phase.counterZ0Z_23 ));
    Odrv4 I__9297 (
            .O(N__41475),
            .I(\current_shift_inst.timer_phase.counterZ0Z_23 ));
    InMux I__9296 (
            .O(N__41470),
            .I(N__41465));
    InMux I__9295 (
            .O(N__41469),
            .I(N__41460));
    InMux I__9294 (
            .O(N__41468),
            .I(N__41460));
    LocalMux I__9293 (
            .O(N__41465),
            .I(N__41457));
    LocalMux I__9292 (
            .O(N__41460),
            .I(N__41454));
    Span4Mux_h I__9291 (
            .O(N__41457),
            .I(N__41451));
    Span12Mux_v I__9290 (
            .O(N__41454),
            .I(N__41447));
    Span4Mux_v I__9289 (
            .O(N__41451),
            .I(N__41444));
    InMux I__9288 (
            .O(N__41450),
            .I(N__41441));
    Odrv12 I__9287 (
            .O(N__41447),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    Odrv4 I__9286 (
            .O(N__41444),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    LocalMux I__9285 (
            .O(N__41441),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    InMux I__9284 (
            .O(N__41434),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ));
    InMux I__9283 (
            .O(N__41431),
            .I(N__41427));
    InMux I__9282 (
            .O(N__41430),
            .I(N__41423));
    LocalMux I__9281 (
            .O(N__41427),
            .I(N__41420));
    InMux I__9280 (
            .O(N__41426),
            .I(N__41417));
    LocalMux I__9279 (
            .O(N__41423),
            .I(N__41412));
    Span4Mux_v I__9278 (
            .O(N__41420),
            .I(N__41412));
    LocalMux I__9277 (
            .O(N__41417),
            .I(\current_shift_inst.timer_phase.counterZ0Z_24 ));
    Odrv4 I__9276 (
            .O(N__41412),
            .I(\current_shift_inst.timer_phase.counterZ0Z_24 ));
    InMux I__9275 (
            .O(N__41407),
            .I(N__41402));
    InMux I__9274 (
            .O(N__41406),
            .I(N__41397));
    InMux I__9273 (
            .O(N__41405),
            .I(N__41397));
    LocalMux I__9272 (
            .O(N__41402),
            .I(N__41394));
    LocalMux I__9271 (
            .O(N__41397),
            .I(N__41391));
    Span4Mux_v I__9270 (
            .O(N__41394),
            .I(N__41388));
    Span4Mux_h I__9269 (
            .O(N__41391),
            .I(N__41385));
    Span4Mux_v I__9268 (
            .O(N__41388),
            .I(N__41381));
    Span4Mux_v I__9267 (
            .O(N__41385),
            .I(N__41378));
    InMux I__9266 (
            .O(N__41384),
            .I(N__41375));
    Odrv4 I__9265 (
            .O(N__41381),
            .I(\current_shift_inst.elapsed_time_ns_phase_27 ));
    Odrv4 I__9264 (
            .O(N__41378),
            .I(\current_shift_inst.elapsed_time_ns_phase_27 ));
    LocalMux I__9263 (
            .O(N__41375),
            .I(\current_shift_inst.elapsed_time_ns_phase_27 ));
    InMux I__9262 (
            .O(N__41368),
            .I(bfn_16_25_0_));
    CascadeMux I__9261 (
            .O(N__41365),
            .I(N__41361));
    InMux I__9260 (
            .O(N__41364),
            .I(N__41358));
    InMux I__9259 (
            .O(N__41361),
            .I(N__41355));
    LocalMux I__9258 (
            .O(N__41358),
            .I(N__41349));
    LocalMux I__9257 (
            .O(N__41355),
            .I(N__41349));
    InMux I__9256 (
            .O(N__41354),
            .I(N__41346));
    Span4Mux_v I__9255 (
            .O(N__41349),
            .I(N__41343));
    LocalMux I__9254 (
            .O(N__41346),
            .I(\current_shift_inst.timer_phase.counterZ0Z_25 ));
    Odrv4 I__9253 (
            .O(N__41343),
            .I(\current_shift_inst.timer_phase.counterZ0Z_25 ));
    InMux I__9252 (
            .O(N__41338),
            .I(N__41333));
    InMux I__9251 (
            .O(N__41337),
            .I(N__41330));
    InMux I__9250 (
            .O(N__41336),
            .I(N__41327));
    LocalMux I__9249 (
            .O(N__41333),
            .I(N__41324));
    LocalMux I__9248 (
            .O(N__41330),
            .I(N__41321));
    LocalMux I__9247 (
            .O(N__41327),
            .I(N__41318));
    Span4Mux_h I__9246 (
            .O(N__41324),
            .I(N__41315));
    Span4Mux_h I__9245 (
            .O(N__41321),
            .I(N__41312));
    Span12Mux_v I__9244 (
            .O(N__41318),
            .I(N__41308));
    Span4Mux_v I__9243 (
            .O(N__41315),
            .I(N__41305));
    Span4Mux_v I__9242 (
            .O(N__41312),
            .I(N__41302));
    InMux I__9241 (
            .O(N__41311),
            .I(N__41299));
    Odrv12 I__9240 (
            .O(N__41308),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    Odrv4 I__9239 (
            .O(N__41305),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    Odrv4 I__9238 (
            .O(N__41302),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    LocalMux I__9237 (
            .O(N__41299),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    InMux I__9236 (
            .O(N__41290),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ));
    InMux I__9235 (
            .O(N__41287),
            .I(N__41283));
    InMux I__9234 (
            .O(N__41286),
            .I(N__41280));
    LocalMux I__9233 (
            .O(N__41283),
            .I(N__41277));
    LocalMux I__9232 (
            .O(N__41280),
            .I(\current_shift_inst.timer_phase.counterZ0Z_28 ));
    Odrv12 I__9231 (
            .O(N__41277),
            .I(\current_shift_inst.timer_phase.counterZ0Z_28 ));
    CascadeMux I__9230 (
            .O(N__41272),
            .I(N__41267));
    CascadeMux I__9229 (
            .O(N__41271),
            .I(N__41264));
    InMux I__9228 (
            .O(N__41270),
            .I(N__41261));
    InMux I__9227 (
            .O(N__41267),
            .I(N__41256));
    InMux I__9226 (
            .O(N__41264),
            .I(N__41256));
    LocalMux I__9225 (
            .O(N__41261),
            .I(N__41251));
    LocalMux I__9224 (
            .O(N__41256),
            .I(N__41251));
    Odrv4 I__9223 (
            .O(N__41251),
            .I(\current_shift_inst.timer_phase.counterZ0Z_26 ));
    InMux I__9222 (
            .O(N__41248),
            .I(N__41244));
    InMux I__9221 (
            .O(N__41247),
            .I(N__41241));
    LocalMux I__9220 (
            .O(N__41244),
            .I(N__41238));
    LocalMux I__9219 (
            .O(N__41241),
            .I(N__41235));
    Span4Mux_v I__9218 (
            .O(N__41238),
            .I(N__41232));
    Span12Mux_v I__9217 (
            .O(N__41235),
            .I(N__41228));
    Span4Mux_h I__9216 (
            .O(N__41232),
            .I(N__41225));
    InMux I__9215 (
            .O(N__41231),
            .I(N__41222));
    Odrv12 I__9214 (
            .O(N__41228),
            .I(\current_shift_inst.elapsed_time_ns_phase_29 ));
    Odrv4 I__9213 (
            .O(N__41225),
            .I(\current_shift_inst.elapsed_time_ns_phase_29 ));
    LocalMux I__9212 (
            .O(N__41222),
            .I(\current_shift_inst.elapsed_time_ns_phase_29 ));
    InMux I__9211 (
            .O(N__41215),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ));
    InMux I__9210 (
            .O(N__41212),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ));
    InMux I__9209 (
            .O(N__41209),
            .I(N__41202));
    InMux I__9208 (
            .O(N__41208),
            .I(N__41202));
    InMux I__9207 (
            .O(N__41207),
            .I(N__41199));
    LocalMux I__9206 (
            .O(N__41202),
            .I(N__41196));
    LocalMux I__9205 (
            .O(N__41199),
            .I(\current_shift_inst.timer_phase.counterZ0Z_12 ));
    Odrv12 I__9204 (
            .O(N__41196),
            .I(\current_shift_inst.timer_phase.counterZ0Z_12 ));
    InMux I__9203 (
            .O(N__41191),
            .I(N__41187));
    InMux I__9202 (
            .O(N__41190),
            .I(N__41184));
    LocalMux I__9201 (
            .O(N__41187),
            .I(N__41180));
    LocalMux I__9200 (
            .O(N__41184),
            .I(N__41177));
    InMux I__9199 (
            .O(N__41183),
            .I(N__41174));
    Span4Mux_v I__9198 (
            .O(N__41180),
            .I(N__41171));
    Span4Mux_h I__9197 (
            .O(N__41177),
            .I(N__41166));
    LocalMux I__9196 (
            .O(N__41174),
            .I(N__41166));
    Span4Mux_v I__9195 (
            .O(N__41171),
            .I(N__41163));
    Span4Mux_v I__9194 (
            .O(N__41166),
            .I(N__41160));
    Span4Mux_h I__9193 (
            .O(N__41163),
            .I(N__41156));
    Span4Mux_h I__9192 (
            .O(N__41160),
            .I(N__41153));
    InMux I__9191 (
            .O(N__41159),
            .I(N__41150));
    Odrv4 I__9190 (
            .O(N__41156),
            .I(\current_shift_inst.elapsed_time_ns_phase_15 ));
    Odrv4 I__9189 (
            .O(N__41153),
            .I(\current_shift_inst.elapsed_time_ns_phase_15 ));
    LocalMux I__9188 (
            .O(N__41150),
            .I(\current_shift_inst.elapsed_time_ns_phase_15 ));
    InMux I__9187 (
            .O(N__41143),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__9186 (
            .O(N__41140),
            .I(N__41136));
    CascadeMux I__9185 (
            .O(N__41139),
            .I(N__41133));
    InMux I__9184 (
            .O(N__41136),
            .I(N__41127));
    InMux I__9183 (
            .O(N__41133),
            .I(N__41127));
    InMux I__9182 (
            .O(N__41132),
            .I(N__41124));
    LocalMux I__9181 (
            .O(N__41127),
            .I(N__41121));
    LocalMux I__9180 (
            .O(N__41124),
            .I(\current_shift_inst.timer_phase.counterZ0Z_13 ));
    Odrv4 I__9179 (
            .O(N__41121),
            .I(\current_shift_inst.timer_phase.counterZ0Z_13 ));
    CascadeMux I__9178 (
            .O(N__41116),
            .I(N__41112));
    InMux I__9177 (
            .O(N__41115),
            .I(N__41108));
    InMux I__9176 (
            .O(N__41112),
            .I(N__41105));
    InMux I__9175 (
            .O(N__41111),
            .I(N__41102));
    LocalMux I__9174 (
            .O(N__41108),
            .I(N__41099));
    LocalMux I__9173 (
            .O(N__41105),
            .I(N__41094));
    LocalMux I__9172 (
            .O(N__41102),
            .I(N__41094));
    Span4Mux_h I__9171 (
            .O(N__41099),
            .I(N__41091));
    Span12Mux_h I__9170 (
            .O(N__41094),
            .I(N__41087));
    Span4Mux_v I__9169 (
            .O(N__41091),
            .I(N__41084));
    InMux I__9168 (
            .O(N__41090),
            .I(N__41081));
    Odrv12 I__9167 (
            .O(N__41087),
            .I(\current_shift_inst.elapsed_time_ns_phase_16 ));
    Odrv4 I__9166 (
            .O(N__41084),
            .I(\current_shift_inst.elapsed_time_ns_phase_16 ));
    LocalMux I__9165 (
            .O(N__41081),
            .I(\current_shift_inst.elapsed_time_ns_phase_16 ));
    InMux I__9164 (
            .O(N__41074),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__9163 (
            .O(N__41071),
            .I(N__41067));
    CascadeMux I__9162 (
            .O(N__41070),
            .I(N__41064));
    InMux I__9161 (
            .O(N__41067),
            .I(N__41058));
    InMux I__9160 (
            .O(N__41064),
            .I(N__41058));
    InMux I__9159 (
            .O(N__41063),
            .I(N__41055));
    LocalMux I__9158 (
            .O(N__41058),
            .I(N__41052));
    LocalMux I__9157 (
            .O(N__41055),
            .I(\current_shift_inst.timer_phase.counterZ0Z_14 ));
    Odrv12 I__9156 (
            .O(N__41052),
            .I(\current_shift_inst.timer_phase.counterZ0Z_14 ));
    InMux I__9155 (
            .O(N__41047),
            .I(N__41044));
    LocalMux I__9154 (
            .O(N__41044),
            .I(N__41040));
    InMux I__9153 (
            .O(N__41043),
            .I(N__41037));
    Span4Mux_h I__9152 (
            .O(N__41040),
            .I(N__41031));
    LocalMux I__9151 (
            .O(N__41037),
            .I(N__41031));
    InMux I__9150 (
            .O(N__41036),
            .I(N__41028));
    Span4Mux_h I__9149 (
            .O(N__41031),
            .I(N__41025));
    LocalMux I__9148 (
            .O(N__41028),
            .I(N__41022));
    Span4Mux_v I__9147 (
            .O(N__41025),
            .I(N__41018));
    Span12Mux_h I__9146 (
            .O(N__41022),
            .I(N__41015));
    InMux I__9145 (
            .O(N__41021),
            .I(N__41012));
    Odrv4 I__9144 (
            .O(N__41018),
            .I(\current_shift_inst.elapsed_time_ns_phase_17 ));
    Odrv12 I__9143 (
            .O(N__41015),
            .I(\current_shift_inst.elapsed_time_ns_phase_17 ));
    LocalMux I__9142 (
            .O(N__41012),
            .I(\current_shift_inst.elapsed_time_ns_phase_17 ));
    InMux I__9141 (
            .O(N__41005),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ));
    InMux I__9140 (
            .O(N__41002),
            .I(N__40995));
    InMux I__9139 (
            .O(N__41001),
            .I(N__40995));
    InMux I__9138 (
            .O(N__41000),
            .I(N__40992));
    LocalMux I__9137 (
            .O(N__40995),
            .I(N__40989));
    LocalMux I__9136 (
            .O(N__40992),
            .I(\current_shift_inst.timer_phase.counterZ0Z_15 ));
    Odrv12 I__9135 (
            .O(N__40989),
            .I(\current_shift_inst.timer_phase.counterZ0Z_15 ));
    InMux I__9134 (
            .O(N__40984),
            .I(N__40979));
    InMux I__9133 (
            .O(N__40983),
            .I(N__40974));
    InMux I__9132 (
            .O(N__40982),
            .I(N__40974));
    LocalMux I__9131 (
            .O(N__40979),
            .I(N__40971));
    LocalMux I__9130 (
            .O(N__40974),
            .I(N__40968));
    Span4Mux_h I__9129 (
            .O(N__40971),
            .I(N__40965));
    Span4Mux_h I__9128 (
            .O(N__40968),
            .I(N__40962));
    Span4Mux_v I__9127 (
            .O(N__40965),
            .I(N__40959));
    Span4Mux_v I__9126 (
            .O(N__40962),
            .I(N__40955));
    Span4Mux_h I__9125 (
            .O(N__40959),
            .I(N__40952));
    InMux I__9124 (
            .O(N__40958),
            .I(N__40949));
    Odrv4 I__9123 (
            .O(N__40955),
            .I(\current_shift_inst.elapsed_time_ns_phase_18 ));
    Odrv4 I__9122 (
            .O(N__40952),
            .I(\current_shift_inst.elapsed_time_ns_phase_18 ));
    LocalMux I__9121 (
            .O(N__40949),
            .I(\current_shift_inst.elapsed_time_ns_phase_18 ));
    InMux I__9120 (
            .O(N__40942),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ));
    InMux I__9119 (
            .O(N__40939),
            .I(N__40935));
    InMux I__9118 (
            .O(N__40938),
            .I(N__40932));
    LocalMux I__9117 (
            .O(N__40935),
            .I(N__40929));
    LocalMux I__9116 (
            .O(N__40932),
            .I(N__40923));
    Span4Mux_v I__9115 (
            .O(N__40929),
            .I(N__40923));
    InMux I__9114 (
            .O(N__40928),
            .I(N__40920));
    Span4Mux_h I__9113 (
            .O(N__40923),
            .I(N__40917));
    LocalMux I__9112 (
            .O(N__40920),
            .I(\current_shift_inst.timer_phase.counterZ0Z_16 ));
    Odrv4 I__9111 (
            .O(N__40917),
            .I(\current_shift_inst.timer_phase.counterZ0Z_16 ));
    InMux I__9110 (
            .O(N__40912),
            .I(N__40906));
    InMux I__9109 (
            .O(N__40911),
            .I(N__40906));
    LocalMux I__9108 (
            .O(N__40906),
            .I(N__40902));
    InMux I__9107 (
            .O(N__40905),
            .I(N__40899));
    Span4Mux_h I__9106 (
            .O(N__40902),
            .I(N__40894));
    LocalMux I__9105 (
            .O(N__40899),
            .I(N__40894));
    Span4Mux_v I__9104 (
            .O(N__40894),
            .I(N__40891));
    Span4Mux_v I__9103 (
            .O(N__40891),
            .I(N__40888));
    Span4Mux_h I__9102 (
            .O(N__40888),
            .I(N__40884));
    InMux I__9101 (
            .O(N__40887),
            .I(N__40881));
    Odrv4 I__9100 (
            .O(N__40884),
            .I(\current_shift_inst.elapsed_time_ns_phase_19 ));
    LocalMux I__9099 (
            .O(N__40881),
            .I(\current_shift_inst.elapsed_time_ns_phase_19 ));
    InMux I__9098 (
            .O(N__40876),
            .I(bfn_16_24_0_));
    CascadeMux I__9097 (
            .O(N__40873),
            .I(N__40870));
    InMux I__9096 (
            .O(N__40870),
            .I(N__40867));
    LocalMux I__9095 (
            .O(N__40867),
            .I(N__40863));
    InMux I__9094 (
            .O(N__40866),
            .I(N__40859));
    Span4Mux_v I__9093 (
            .O(N__40863),
            .I(N__40856));
    InMux I__9092 (
            .O(N__40862),
            .I(N__40853));
    LocalMux I__9091 (
            .O(N__40859),
            .I(N__40848));
    Span4Mux_h I__9090 (
            .O(N__40856),
            .I(N__40848));
    LocalMux I__9089 (
            .O(N__40853),
            .I(\current_shift_inst.timer_phase.counterZ0Z_17 ));
    Odrv4 I__9088 (
            .O(N__40848),
            .I(\current_shift_inst.timer_phase.counterZ0Z_17 ));
    InMux I__9087 (
            .O(N__40843),
            .I(N__40839));
    InMux I__9086 (
            .O(N__40842),
            .I(N__40835));
    LocalMux I__9085 (
            .O(N__40839),
            .I(N__40832));
    InMux I__9084 (
            .O(N__40838),
            .I(N__40829));
    LocalMux I__9083 (
            .O(N__40835),
            .I(N__40826));
    Span4Mux_h I__9082 (
            .O(N__40832),
            .I(N__40821));
    LocalMux I__9081 (
            .O(N__40829),
            .I(N__40821));
    Sp12to4 I__9080 (
            .O(N__40826),
            .I(N__40818));
    Span4Mux_h I__9079 (
            .O(N__40821),
            .I(N__40815));
    Span12Mux_v I__9078 (
            .O(N__40818),
            .I(N__40811));
    Span4Mux_v I__9077 (
            .O(N__40815),
            .I(N__40808));
    InMux I__9076 (
            .O(N__40814),
            .I(N__40805));
    Odrv12 I__9075 (
            .O(N__40811),
            .I(\current_shift_inst.elapsed_time_ns_phase_20 ));
    Odrv4 I__9074 (
            .O(N__40808),
            .I(\current_shift_inst.elapsed_time_ns_phase_20 ));
    LocalMux I__9073 (
            .O(N__40805),
            .I(\current_shift_inst.elapsed_time_ns_phase_20 ));
    InMux I__9072 (
            .O(N__40798),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__9071 (
            .O(N__40795),
            .I(N__40790));
    InMux I__9070 (
            .O(N__40794),
            .I(N__40787));
    InMux I__9069 (
            .O(N__40793),
            .I(N__40784));
    InMux I__9068 (
            .O(N__40790),
            .I(N__40781));
    LocalMux I__9067 (
            .O(N__40787),
            .I(N__40774));
    LocalMux I__9066 (
            .O(N__40784),
            .I(N__40774));
    LocalMux I__9065 (
            .O(N__40781),
            .I(N__40774));
    Odrv4 I__9064 (
            .O(N__40774),
            .I(\current_shift_inst.timer_phase.counterZ0Z_18 ));
    InMux I__9063 (
            .O(N__40771),
            .I(N__40765));
    InMux I__9062 (
            .O(N__40770),
            .I(N__40765));
    LocalMux I__9061 (
            .O(N__40765),
            .I(N__40761));
    InMux I__9060 (
            .O(N__40764),
            .I(N__40758));
    Span4Mux_h I__9059 (
            .O(N__40761),
            .I(N__40755));
    LocalMux I__9058 (
            .O(N__40758),
            .I(N__40752));
    Span4Mux_v I__9057 (
            .O(N__40755),
            .I(N__40749));
    Span12Mux_h I__9056 (
            .O(N__40752),
            .I(N__40745));
    Span4Mux_h I__9055 (
            .O(N__40749),
            .I(N__40742));
    InMux I__9054 (
            .O(N__40748),
            .I(N__40739));
    Odrv12 I__9053 (
            .O(N__40745),
            .I(\current_shift_inst.elapsed_time_ns_phase_21 ));
    Odrv4 I__9052 (
            .O(N__40742),
            .I(\current_shift_inst.elapsed_time_ns_phase_21 ));
    LocalMux I__9051 (
            .O(N__40739),
            .I(\current_shift_inst.elapsed_time_ns_phase_21 ));
    InMux I__9050 (
            .O(N__40732),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__9049 (
            .O(N__40729),
            .I(N__40725));
    CascadeMux I__9048 (
            .O(N__40728),
            .I(N__40722));
    InMux I__9047 (
            .O(N__40725),
            .I(N__40716));
    InMux I__9046 (
            .O(N__40722),
            .I(N__40716));
    InMux I__9045 (
            .O(N__40721),
            .I(N__40713));
    LocalMux I__9044 (
            .O(N__40716),
            .I(N__40710));
    LocalMux I__9043 (
            .O(N__40713),
            .I(\current_shift_inst.timer_phase.counterZ0Z_4 ));
    Odrv4 I__9042 (
            .O(N__40710),
            .I(\current_shift_inst.timer_phase.counterZ0Z_4 ));
    CascadeMux I__9041 (
            .O(N__40705),
            .I(N__40702));
    InMux I__9040 (
            .O(N__40702),
            .I(N__40698));
    CascadeMux I__9039 (
            .O(N__40701),
            .I(N__40694));
    LocalMux I__9038 (
            .O(N__40698),
            .I(N__40691));
    InMux I__9037 (
            .O(N__40697),
            .I(N__40686));
    InMux I__9036 (
            .O(N__40694),
            .I(N__40686));
    Span4Mux_v I__9035 (
            .O(N__40691),
            .I(N__40683));
    LocalMux I__9034 (
            .O(N__40686),
            .I(N__40680));
    Span4Mux_h I__9033 (
            .O(N__40683),
            .I(N__40676));
    Sp12to4 I__9032 (
            .O(N__40680),
            .I(N__40673));
    InMux I__9031 (
            .O(N__40679),
            .I(N__40670));
    Odrv4 I__9030 (
            .O(N__40676),
            .I(\current_shift_inst.elapsed_time_ns_phase_7 ));
    Odrv12 I__9029 (
            .O(N__40673),
            .I(\current_shift_inst.elapsed_time_ns_phase_7 ));
    LocalMux I__9028 (
            .O(N__40670),
            .I(\current_shift_inst.elapsed_time_ns_phase_7 ));
    InMux I__9027 (
            .O(N__40663),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__9026 (
            .O(N__40660),
            .I(N__40656));
    CascadeMux I__9025 (
            .O(N__40659),
            .I(N__40653));
    InMux I__9024 (
            .O(N__40656),
            .I(N__40647));
    InMux I__9023 (
            .O(N__40653),
            .I(N__40647));
    InMux I__9022 (
            .O(N__40652),
            .I(N__40644));
    LocalMux I__9021 (
            .O(N__40647),
            .I(N__40641));
    LocalMux I__9020 (
            .O(N__40644),
            .I(\current_shift_inst.timer_phase.counterZ0Z_5 ));
    Odrv4 I__9019 (
            .O(N__40641),
            .I(\current_shift_inst.timer_phase.counterZ0Z_5 ));
    CascadeMux I__9018 (
            .O(N__40636),
            .I(N__40633));
    InMux I__9017 (
            .O(N__40633),
            .I(N__40629));
    InMux I__9016 (
            .O(N__40632),
            .I(N__40625));
    LocalMux I__9015 (
            .O(N__40629),
            .I(N__40622));
    InMux I__9014 (
            .O(N__40628),
            .I(N__40619));
    LocalMux I__9013 (
            .O(N__40625),
            .I(N__40616));
    Span4Mux_v I__9012 (
            .O(N__40622),
            .I(N__40613));
    LocalMux I__9011 (
            .O(N__40619),
            .I(N__40610));
    Span4Mux_h I__9010 (
            .O(N__40616),
            .I(N__40607));
    Span4Mux_h I__9009 (
            .O(N__40613),
            .I(N__40603));
    Span4Mux_h I__9008 (
            .O(N__40610),
            .I(N__40600));
    Span4Mux_v I__9007 (
            .O(N__40607),
            .I(N__40597));
    InMux I__9006 (
            .O(N__40606),
            .I(N__40594));
    Odrv4 I__9005 (
            .O(N__40603),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    Odrv4 I__9004 (
            .O(N__40600),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    Odrv4 I__9003 (
            .O(N__40597),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    LocalMux I__9002 (
            .O(N__40594),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    InMux I__9001 (
            .O(N__40585),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ));
    InMux I__9000 (
            .O(N__40582),
            .I(N__40575));
    InMux I__8999 (
            .O(N__40581),
            .I(N__40575));
    InMux I__8998 (
            .O(N__40580),
            .I(N__40572));
    LocalMux I__8997 (
            .O(N__40575),
            .I(N__40569));
    LocalMux I__8996 (
            .O(N__40572),
            .I(\current_shift_inst.timer_phase.counterZ0Z_6 ));
    Odrv12 I__8995 (
            .O(N__40569),
            .I(\current_shift_inst.timer_phase.counterZ0Z_6 ));
    InMux I__8994 (
            .O(N__40564),
            .I(N__40557));
    InMux I__8993 (
            .O(N__40563),
            .I(N__40557));
    InMux I__8992 (
            .O(N__40562),
            .I(N__40554));
    LocalMux I__8991 (
            .O(N__40557),
            .I(N__40551));
    LocalMux I__8990 (
            .O(N__40554),
            .I(N__40548));
    Span4Mux_h I__8989 (
            .O(N__40551),
            .I(N__40545));
    Span4Mux_h I__8988 (
            .O(N__40548),
            .I(N__40542));
    Span4Mux_h I__8987 (
            .O(N__40545),
            .I(N__40538));
    Span4Mux_h I__8986 (
            .O(N__40542),
            .I(N__40535));
    InMux I__8985 (
            .O(N__40541),
            .I(N__40532));
    Odrv4 I__8984 (
            .O(N__40538),
            .I(\current_shift_inst.elapsed_time_ns_phase_9 ));
    Odrv4 I__8983 (
            .O(N__40535),
            .I(\current_shift_inst.elapsed_time_ns_phase_9 ));
    LocalMux I__8982 (
            .O(N__40532),
            .I(\current_shift_inst.elapsed_time_ns_phase_9 ));
    InMux I__8981 (
            .O(N__40525),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ));
    InMux I__8980 (
            .O(N__40522),
            .I(N__40515));
    InMux I__8979 (
            .O(N__40521),
            .I(N__40515));
    InMux I__8978 (
            .O(N__40520),
            .I(N__40512));
    LocalMux I__8977 (
            .O(N__40515),
            .I(N__40509));
    LocalMux I__8976 (
            .O(N__40512),
            .I(\current_shift_inst.timer_phase.counterZ0Z_7 ));
    Odrv12 I__8975 (
            .O(N__40509),
            .I(\current_shift_inst.timer_phase.counterZ0Z_7 ));
    InMux I__8974 (
            .O(N__40504),
            .I(N__40499));
    InMux I__8973 (
            .O(N__40503),
            .I(N__40496));
    InMux I__8972 (
            .O(N__40502),
            .I(N__40493));
    LocalMux I__8971 (
            .O(N__40499),
            .I(N__40490));
    LocalMux I__8970 (
            .O(N__40496),
            .I(N__40487));
    LocalMux I__8969 (
            .O(N__40493),
            .I(N__40484));
    Span4Mux_h I__8968 (
            .O(N__40490),
            .I(N__40481));
    Span4Mux_h I__8967 (
            .O(N__40487),
            .I(N__40478));
    Span4Mux_v I__8966 (
            .O(N__40484),
            .I(N__40473));
    Span4Mux_v I__8965 (
            .O(N__40481),
            .I(N__40473));
    Span4Mux_h I__8964 (
            .O(N__40478),
            .I(N__40469));
    Span4Mux_h I__8963 (
            .O(N__40473),
            .I(N__40466));
    InMux I__8962 (
            .O(N__40472),
            .I(N__40463));
    Odrv4 I__8961 (
            .O(N__40469),
            .I(\current_shift_inst.elapsed_time_ns_phase_10 ));
    Odrv4 I__8960 (
            .O(N__40466),
            .I(\current_shift_inst.elapsed_time_ns_phase_10 ));
    LocalMux I__8959 (
            .O(N__40463),
            .I(\current_shift_inst.elapsed_time_ns_phase_10 ));
    InMux I__8958 (
            .O(N__40456),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__8957 (
            .O(N__40453),
            .I(N__40450));
    InMux I__8956 (
            .O(N__40450),
            .I(N__40447));
    LocalMux I__8955 (
            .O(N__40447),
            .I(N__40443));
    InMux I__8954 (
            .O(N__40446),
            .I(N__40439));
    Span4Mux_v I__8953 (
            .O(N__40443),
            .I(N__40436));
    InMux I__8952 (
            .O(N__40442),
            .I(N__40433));
    LocalMux I__8951 (
            .O(N__40439),
            .I(N__40428));
    Span4Mux_h I__8950 (
            .O(N__40436),
            .I(N__40428));
    LocalMux I__8949 (
            .O(N__40433),
            .I(\current_shift_inst.timer_phase.counterZ0Z_8 ));
    Odrv4 I__8948 (
            .O(N__40428),
            .I(\current_shift_inst.timer_phase.counterZ0Z_8 ));
    CascadeMux I__8947 (
            .O(N__40423),
            .I(N__40420));
    InMux I__8946 (
            .O(N__40420),
            .I(N__40416));
    InMux I__8945 (
            .O(N__40419),
            .I(N__40413));
    LocalMux I__8944 (
            .O(N__40416),
            .I(N__40409));
    LocalMux I__8943 (
            .O(N__40413),
            .I(N__40406));
    InMux I__8942 (
            .O(N__40412),
            .I(N__40403));
    Span4Mux_h I__8941 (
            .O(N__40409),
            .I(N__40400));
    Span4Mux_h I__8940 (
            .O(N__40406),
            .I(N__40397));
    LocalMux I__8939 (
            .O(N__40403),
            .I(N__40394));
    Span4Mux_v I__8938 (
            .O(N__40400),
            .I(N__40390));
    Span4Mux_h I__8937 (
            .O(N__40397),
            .I(N__40387));
    Span12Mux_h I__8936 (
            .O(N__40394),
            .I(N__40384));
    InMux I__8935 (
            .O(N__40393),
            .I(N__40381));
    Odrv4 I__8934 (
            .O(N__40390),
            .I(\current_shift_inst.elapsed_time_ns_phase_11 ));
    Odrv4 I__8933 (
            .O(N__40387),
            .I(\current_shift_inst.elapsed_time_ns_phase_11 ));
    Odrv12 I__8932 (
            .O(N__40384),
            .I(\current_shift_inst.elapsed_time_ns_phase_11 ));
    LocalMux I__8931 (
            .O(N__40381),
            .I(\current_shift_inst.elapsed_time_ns_phase_11 ));
    InMux I__8930 (
            .O(N__40372),
            .I(bfn_16_23_0_));
    CascadeMux I__8929 (
            .O(N__40369),
            .I(N__40365));
    InMux I__8928 (
            .O(N__40368),
            .I(N__40362));
    InMux I__8927 (
            .O(N__40365),
            .I(N__40359));
    LocalMux I__8926 (
            .O(N__40362),
            .I(N__40353));
    LocalMux I__8925 (
            .O(N__40359),
            .I(N__40353));
    InMux I__8924 (
            .O(N__40358),
            .I(N__40350));
    Span4Mux_v I__8923 (
            .O(N__40353),
            .I(N__40347));
    LocalMux I__8922 (
            .O(N__40350),
            .I(\current_shift_inst.timer_phase.counterZ0Z_9 ));
    Odrv4 I__8921 (
            .O(N__40347),
            .I(\current_shift_inst.timer_phase.counterZ0Z_9 ));
    InMux I__8920 (
            .O(N__40342),
            .I(N__40337));
    InMux I__8919 (
            .O(N__40341),
            .I(N__40332));
    InMux I__8918 (
            .O(N__40340),
            .I(N__40332));
    LocalMux I__8917 (
            .O(N__40337),
            .I(N__40329));
    LocalMux I__8916 (
            .O(N__40332),
            .I(N__40326));
    Span4Mux_h I__8915 (
            .O(N__40329),
            .I(N__40323));
    Span4Mux_h I__8914 (
            .O(N__40326),
            .I(N__40320));
    Span4Mux_h I__8913 (
            .O(N__40323),
            .I(N__40316));
    Span4Mux_v I__8912 (
            .O(N__40320),
            .I(N__40313));
    InMux I__8911 (
            .O(N__40319),
            .I(N__40310));
    Odrv4 I__8910 (
            .O(N__40316),
            .I(\current_shift_inst.elapsed_time_ns_phase_12 ));
    Odrv4 I__8909 (
            .O(N__40313),
            .I(\current_shift_inst.elapsed_time_ns_phase_12 ));
    LocalMux I__8908 (
            .O(N__40310),
            .I(\current_shift_inst.elapsed_time_ns_phase_12 ));
    InMux I__8907 (
            .O(N__40303),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__8906 (
            .O(N__40300),
            .I(N__40295));
    CascadeMux I__8905 (
            .O(N__40299),
            .I(N__40292));
    InMux I__8904 (
            .O(N__40298),
            .I(N__40289));
    InMux I__8903 (
            .O(N__40295),
            .I(N__40284));
    InMux I__8902 (
            .O(N__40292),
            .I(N__40284));
    LocalMux I__8901 (
            .O(N__40289),
            .I(N__40279));
    LocalMux I__8900 (
            .O(N__40284),
            .I(N__40279));
    Odrv4 I__8899 (
            .O(N__40279),
            .I(\current_shift_inst.timer_phase.counterZ0Z_10 ));
    CascadeMux I__8898 (
            .O(N__40276),
            .I(N__40273));
    InMux I__8897 (
            .O(N__40273),
            .I(N__40270));
    LocalMux I__8896 (
            .O(N__40270),
            .I(N__40266));
    InMux I__8895 (
            .O(N__40269),
            .I(N__40262));
    Span4Mux_h I__8894 (
            .O(N__40266),
            .I(N__40259));
    InMux I__8893 (
            .O(N__40265),
            .I(N__40256));
    LocalMux I__8892 (
            .O(N__40262),
            .I(N__40253));
    Span4Mux_h I__8891 (
            .O(N__40259),
            .I(N__40250));
    LocalMux I__8890 (
            .O(N__40256),
            .I(N__40247));
    Span4Mux_h I__8889 (
            .O(N__40253),
            .I(N__40244));
    Sp12to4 I__8888 (
            .O(N__40250),
            .I(N__40240));
    Span12Mux_h I__8887 (
            .O(N__40247),
            .I(N__40237));
    Span4Mux_v I__8886 (
            .O(N__40244),
            .I(N__40234));
    InMux I__8885 (
            .O(N__40243),
            .I(N__40231));
    Odrv12 I__8884 (
            .O(N__40240),
            .I(\current_shift_inst.elapsed_time_ns_phase_13 ));
    Odrv12 I__8883 (
            .O(N__40237),
            .I(\current_shift_inst.elapsed_time_ns_phase_13 ));
    Odrv4 I__8882 (
            .O(N__40234),
            .I(\current_shift_inst.elapsed_time_ns_phase_13 ));
    LocalMux I__8881 (
            .O(N__40231),
            .I(\current_shift_inst.elapsed_time_ns_phase_13 ));
    InMux I__8880 (
            .O(N__40222),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__8879 (
            .O(N__40219),
            .I(N__40214));
    InMux I__8878 (
            .O(N__40218),
            .I(N__40211));
    InMux I__8877 (
            .O(N__40217),
            .I(N__40208));
    InMux I__8876 (
            .O(N__40214),
            .I(N__40205));
    LocalMux I__8875 (
            .O(N__40211),
            .I(N__40198));
    LocalMux I__8874 (
            .O(N__40208),
            .I(N__40198));
    LocalMux I__8873 (
            .O(N__40205),
            .I(N__40198));
    Odrv4 I__8872 (
            .O(N__40198),
            .I(\current_shift_inst.timer_phase.counterZ0Z_11 ));
    InMux I__8871 (
            .O(N__40195),
            .I(N__40190));
    InMux I__8870 (
            .O(N__40194),
            .I(N__40187));
    InMux I__8869 (
            .O(N__40193),
            .I(N__40184));
    LocalMux I__8868 (
            .O(N__40190),
            .I(N__40181));
    LocalMux I__8867 (
            .O(N__40187),
            .I(N__40178));
    LocalMux I__8866 (
            .O(N__40184),
            .I(N__40175));
    Span4Mux_h I__8865 (
            .O(N__40181),
            .I(N__40170));
    Span4Mux_v I__8864 (
            .O(N__40178),
            .I(N__40170));
    Span4Mux_v I__8863 (
            .O(N__40175),
            .I(N__40167));
    Span4Mux_v I__8862 (
            .O(N__40170),
            .I(N__40164));
    Span4Mux_v I__8861 (
            .O(N__40167),
            .I(N__40160));
    Span4Mux_h I__8860 (
            .O(N__40164),
            .I(N__40157));
    InMux I__8859 (
            .O(N__40163),
            .I(N__40154));
    Odrv4 I__8858 (
            .O(N__40160),
            .I(\current_shift_inst.elapsed_time_ns_phase_14 ));
    Odrv4 I__8857 (
            .O(N__40157),
            .I(\current_shift_inst.elapsed_time_ns_phase_14 ));
    LocalMux I__8856 (
            .O(N__40154),
            .I(\current_shift_inst.elapsed_time_ns_phase_14 ));
    InMux I__8855 (
            .O(N__40147),
            .I(N__40144));
    LocalMux I__8854 (
            .O(N__40144),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5 ));
    CascadeMux I__8853 (
            .O(N__40141),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4_cascade_ ));
    InMux I__8852 (
            .O(N__40138),
            .I(N__40135));
    LocalMux I__8851 (
            .O(N__40135),
            .I(N__40132));
    Odrv4 I__8850 (
            .O(N__40132),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6 ));
    InMux I__8849 (
            .O(N__40129),
            .I(N__40126));
    LocalMux I__8848 (
            .O(N__40126),
            .I(N__40122));
    InMux I__8847 (
            .O(N__40125),
            .I(N__40119));
    Span4Mux_h I__8846 (
            .O(N__40122),
            .I(N__40115));
    LocalMux I__8845 (
            .O(N__40119),
            .I(N__40112));
    InMux I__8844 (
            .O(N__40118),
            .I(N__40109));
    Odrv4 I__8843 (
            .O(N__40115),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    Odrv4 I__8842 (
            .O(N__40112),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    LocalMux I__8841 (
            .O(N__40109),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    InMux I__8840 (
            .O(N__40102),
            .I(N__40096));
    InMux I__8839 (
            .O(N__40101),
            .I(N__40096));
    LocalMux I__8838 (
            .O(N__40096),
            .I(N__40092));
    InMux I__8837 (
            .O(N__40095),
            .I(N__40089));
    Odrv4 I__8836 (
            .O(N__40092),
            .I(\current_shift_inst.elapsed_time_ns_phase_3 ));
    LocalMux I__8835 (
            .O(N__40089),
            .I(\current_shift_inst.elapsed_time_ns_phase_3 ));
    InMux I__8834 (
            .O(N__40084),
            .I(N__40079));
    InMux I__8833 (
            .O(N__40083),
            .I(N__40076));
    InMux I__8832 (
            .O(N__40082),
            .I(N__40073));
    LocalMux I__8831 (
            .O(N__40079),
            .I(N__40070));
    LocalMux I__8830 (
            .O(N__40076),
            .I(N__40065));
    LocalMux I__8829 (
            .O(N__40073),
            .I(N__40065));
    Odrv4 I__8828 (
            .O(N__40070),
            .I(\current_shift_inst.timer_phase.counterZ0Z_1 ));
    Odrv4 I__8827 (
            .O(N__40065),
            .I(\current_shift_inst.timer_phase.counterZ0Z_1 ));
    InMux I__8826 (
            .O(N__40060),
            .I(N__40053));
    InMux I__8825 (
            .O(N__40059),
            .I(N__40053));
    InMux I__8824 (
            .O(N__40058),
            .I(N__40050));
    LocalMux I__8823 (
            .O(N__40053),
            .I(N__40047));
    LocalMux I__8822 (
            .O(N__40050),
            .I(N__40044));
    Span4Mux_h I__8821 (
            .O(N__40047),
            .I(N__40041));
    Span4Mux_h I__8820 (
            .O(N__40044),
            .I(N__40038));
    Span4Mux_h I__8819 (
            .O(N__40041),
            .I(N__40034));
    Span4Mux_h I__8818 (
            .O(N__40038),
            .I(N__40031));
    InMux I__8817 (
            .O(N__40037),
            .I(N__40028));
    Odrv4 I__8816 (
            .O(N__40034),
            .I(\current_shift_inst.elapsed_time_ns_phase_4 ));
    Odrv4 I__8815 (
            .O(N__40031),
            .I(\current_shift_inst.elapsed_time_ns_phase_4 ));
    LocalMux I__8814 (
            .O(N__40028),
            .I(\current_shift_inst.elapsed_time_ns_phase_4 ));
    InMux I__8813 (
            .O(N__40021),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__8812 (
            .O(N__40018),
            .I(N__40013));
    InMux I__8811 (
            .O(N__40017),
            .I(N__40010));
    InMux I__8810 (
            .O(N__40016),
            .I(N__40007));
    InMux I__8809 (
            .O(N__40013),
            .I(N__40004));
    LocalMux I__8808 (
            .O(N__40010),
            .I(N__39997));
    LocalMux I__8807 (
            .O(N__40007),
            .I(N__39997));
    LocalMux I__8806 (
            .O(N__40004),
            .I(N__39997));
    Odrv4 I__8805 (
            .O(N__39997),
            .I(\current_shift_inst.timer_phase.counterZ0Z_2 ));
    InMux I__8804 (
            .O(N__39994),
            .I(N__39991));
    LocalMux I__8803 (
            .O(N__39991),
            .I(N__39986));
    InMux I__8802 (
            .O(N__39990),
            .I(N__39983));
    InMux I__8801 (
            .O(N__39989),
            .I(N__39980));
    Span4Mux_v I__8800 (
            .O(N__39986),
            .I(N__39975));
    LocalMux I__8799 (
            .O(N__39983),
            .I(N__39975));
    LocalMux I__8798 (
            .O(N__39980),
            .I(N__39972));
    Sp12to4 I__8797 (
            .O(N__39975),
            .I(N__39966));
    Span12Mux_v I__8796 (
            .O(N__39972),
            .I(N__39966));
    InMux I__8795 (
            .O(N__39971),
            .I(N__39963));
    Odrv12 I__8794 (
            .O(N__39966),
            .I(\current_shift_inst.elapsed_time_ns_phase_5 ));
    LocalMux I__8793 (
            .O(N__39963),
            .I(\current_shift_inst.elapsed_time_ns_phase_5 ));
    InMux I__8792 (
            .O(N__39958),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__8791 (
            .O(N__39955),
            .I(N__39950));
    InMux I__8790 (
            .O(N__39954),
            .I(N__39947));
    InMux I__8789 (
            .O(N__39953),
            .I(N__39944));
    InMux I__8788 (
            .O(N__39950),
            .I(N__39941));
    LocalMux I__8787 (
            .O(N__39947),
            .I(N__39934));
    LocalMux I__8786 (
            .O(N__39944),
            .I(N__39934));
    LocalMux I__8785 (
            .O(N__39941),
            .I(N__39934));
    Odrv4 I__8784 (
            .O(N__39934),
            .I(\current_shift_inst.timer_phase.counterZ0Z_3 ));
    InMux I__8783 (
            .O(N__39931),
            .I(N__39926));
    InMux I__8782 (
            .O(N__39930),
            .I(N__39921));
    InMux I__8781 (
            .O(N__39929),
            .I(N__39921));
    LocalMux I__8780 (
            .O(N__39926),
            .I(N__39918));
    LocalMux I__8779 (
            .O(N__39921),
            .I(N__39914));
    Span4Mux_h I__8778 (
            .O(N__39918),
            .I(N__39911));
    InMux I__8777 (
            .O(N__39917),
            .I(N__39908));
    Odrv12 I__8776 (
            .O(N__39914),
            .I(\current_shift_inst.elapsed_time_ns_phase_6 ));
    Odrv4 I__8775 (
            .O(N__39911),
            .I(\current_shift_inst.elapsed_time_ns_phase_6 ));
    LocalMux I__8774 (
            .O(N__39908),
            .I(\current_shift_inst.elapsed_time_ns_phase_6 ));
    InMux I__8773 (
            .O(N__39901),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ));
    InMux I__8772 (
            .O(N__39898),
            .I(N__39895));
    LocalMux I__8771 (
            .O(N__39895),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ));
    InMux I__8770 (
            .O(N__39892),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__8769 (
            .O(N__39889),
            .I(N__39886));
    LocalMux I__8768 (
            .O(N__39886),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ));
    InMux I__8767 (
            .O(N__39883),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    CEMux I__8766 (
            .O(N__39880),
            .I(N__39862));
    CEMux I__8765 (
            .O(N__39879),
            .I(N__39862));
    CEMux I__8764 (
            .O(N__39878),
            .I(N__39862));
    CEMux I__8763 (
            .O(N__39877),
            .I(N__39862));
    CEMux I__8762 (
            .O(N__39876),
            .I(N__39862));
    CEMux I__8761 (
            .O(N__39875),
            .I(N__39862));
    GlobalMux I__8760 (
            .O(N__39862),
            .I(N__39859));
    gio2CtrlBuf I__8759 (
            .O(N__39859),
            .I(\current_shift_inst.timer_s1.N_187_i_g ));
    InMux I__8758 (
            .O(N__39856),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__8757 (
            .O(N__39853),
            .I(N__39850));
    LocalMux I__8756 (
            .O(N__39850),
            .I(N__39846));
    InMux I__8755 (
            .O(N__39849),
            .I(N__39843));
    Span4Mux_v I__8754 (
            .O(N__39846),
            .I(N__39838));
    LocalMux I__8753 (
            .O(N__39843),
            .I(N__39838));
    Span4Mux_v I__8752 (
            .O(N__39838),
            .I(N__39835));
    Odrv4 I__8751 (
            .O(N__39835),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__8750 (
            .O(N__39832),
            .I(N__39828));
    InMux I__8749 (
            .O(N__39831),
            .I(N__39825));
    LocalMux I__8748 (
            .O(N__39828),
            .I(N__39821));
    LocalMux I__8747 (
            .O(N__39825),
            .I(N__39818));
    InMux I__8746 (
            .O(N__39824),
            .I(N__39815));
    Span4Mux_v I__8745 (
            .O(N__39821),
            .I(N__39811));
    Span12Mux_v I__8744 (
            .O(N__39818),
            .I(N__39806));
    LocalMux I__8743 (
            .O(N__39815),
            .I(N__39806));
    InMux I__8742 (
            .O(N__39814),
            .I(N__39803));
    Span4Mux_h I__8741 (
            .O(N__39811),
            .I(N__39800));
    Span12Mux_v I__8740 (
            .O(N__39806),
            .I(N__39797));
    LocalMux I__8739 (
            .O(N__39803),
            .I(N__39794));
    Odrv4 I__8738 (
            .O(N__39800),
            .I(measured_delay_tr_18));
    Odrv12 I__8737 (
            .O(N__39797),
            .I(measured_delay_tr_18));
    Odrv4 I__8736 (
            .O(N__39794),
            .I(measured_delay_tr_18));
    InMux I__8735 (
            .O(N__39787),
            .I(N__39783));
    InMux I__8734 (
            .O(N__39786),
            .I(N__39779));
    LocalMux I__8733 (
            .O(N__39783),
            .I(N__39776));
    InMux I__8732 (
            .O(N__39782),
            .I(N__39773));
    LocalMux I__8731 (
            .O(N__39779),
            .I(N__39770));
    Span4Mux_v I__8730 (
            .O(N__39776),
            .I(N__39767));
    LocalMux I__8729 (
            .O(N__39773),
            .I(N__39764));
    Span4Mux_v I__8728 (
            .O(N__39770),
            .I(N__39760));
    Span4Mux_v I__8727 (
            .O(N__39767),
            .I(N__39755));
    Span4Mux_v I__8726 (
            .O(N__39764),
            .I(N__39755));
    InMux I__8725 (
            .O(N__39763),
            .I(N__39752));
    Odrv4 I__8724 (
            .O(N__39760),
            .I(measured_delay_tr_17));
    Odrv4 I__8723 (
            .O(N__39755),
            .I(measured_delay_tr_17));
    LocalMux I__8722 (
            .O(N__39752),
            .I(measured_delay_tr_17));
    CascadeMux I__8721 (
            .O(N__39745),
            .I(N__39742));
    InMux I__8720 (
            .O(N__39742),
            .I(N__39737));
    InMux I__8719 (
            .O(N__39741),
            .I(N__39733));
    InMux I__8718 (
            .O(N__39740),
            .I(N__39730));
    LocalMux I__8717 (
            .O(N__39737),
            .I(N__39727));
    CascadeMux I__8716 (
            .O(N__39736),
            .I(N__39724));
    LocalMux I__8715 (
            .O(N__39733),
            .I(N__39721));
    LocalMux I__8714 (
            .O(N__39730),
            .I(N__39718));
    Span4Mux_v I__8713 (
            .O(N__39727),
            .I(N__39715));
    InMux I__8712 (
            .O(N__39724),
            .I(N__39712));
    Span12Mux_h I__8711 (
            .O(N__39721),
            .I(N__39709));
    Span4Mux_v I__8710 (
            .O(N__39718),
            .I(N__39706));
    Span4Mux_h I__8709 (
            .O(N__39715),
            .I(N__39701));
    LocalMux I__8708 (
            .O(N__39712),
            .I(N__39701));
    Odrv12 I__8707 (
            .O(N__39709),
            .I(measured_delay_tr_19));
    Odrv4 I__8706 (
            .O(N__39706),
            .I(measured_delay_tr_19));
    Odrv4 I__8705 (
            .O(N__39701),
            .I(measured_delay_tr_19));
    InMux I__8704 (
            .O(N__39694),
            .I(N__39691));
    LocalMux I__8703 (
            .O(N__39691),
            .I(N__39687));
    InMux I__8702 (
            .O(N__39690),
            .I(N__39684));
    Span4Mux_h I__8701 (
            .O(N__39687),
            .I(N__39680));
    LocalMux I__8700 (
            .O(N__39684),
            .I(N__39677));
    CascadeMux I__8699 (
            .O(N__39683),
            .I(N__39674));
    Span4Mux_v I__8698 (
            .O(N__39680),
            .I(N__39670));
    Span4Mux_h I__8697 (
            .O(N__39677),
            .I(N__39667));
    InMux I__8696 (
            .O(N__39674),
            .I(N__39663));
    InMux I__8695 (
            .O(N__39673),
            .I(N__39660));
    Span4Mux_v I__8694 (
            .O(N__39670),
            .I(N__39655));
    Span4Mux_h I__8693 (
            .O(N__39667),
            .I(N__39655));
    InMux I__8692 (
            .O(N__39666),
            .I(N__39652));
    LocalMux I__8691 (
            .O(N__39663),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__8690 (
            .O(N__39660),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__8689 (
            .O(N__39655),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__8688 (
            .O(N__39652),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    InMux I__8687 (
            .O(N__39643),
            .I(N__39639));
    InMux I__8686 (
            .O(N__39642),
            .I(N__39636));
    LocalMux I__8685 (
            .O(N__39639),
            .I(N__39632));
    LocalMux I__8684 (
            .O(N__39636),
            .I(N__39628));
    InMux I__8683 (
            .O(N__39635),
            .I(N__39625));
    Sp12to4 I__8682 (
            .O(N__39632),
            .I(N__39622));
    InMux I__8681 (
            .O(N__39631),
            .I(N__39619));
    Span12Mux_v I__8680 (
            .O(N__39628),
            .I(N__39616));
    LocalMux I__8679 (
            .O(N__39625),
            .I(N__39611));
    Span12Mux_s11_h I__8678 (
            .O(N__39622),
            .I(N__39611));
    LocalMux I__8677 (
            .O(N__39619),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv12 I__8676 (
            .O(N__39616),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv12 I__8675 (
            .O(N__39611),
            .I(\phase_controller_inst1.tr_time_passed ));
    CascadeMux I__8674 (
            .O(N__39604),
            .I(N__39601));
    InMux I__8673 (
            .O(N__39601),
            .I(N__39598));
    LocalMux I__8672 (
            .O(N__39598),
            .I(N__39594));
    InMux I__8671 (
            .O(N__39597),
            .I(N__39591));
    Span4Mux_h I__8670 (
            .O(N__39594),
            .I(N__39588));
    LocalMux I__8669 (
            .O(N__39591),
            .I(N__39585));
    Span4Mux_h I__8668 (
            .O(N__39588),
            .I(N__39580));
    Span4Mux_h I__8667 (
            .O(N__39585),
            .I(N__39576));
    InMux I__8666 (
            .O(N__39584),
            .I(N__39573));
    InMux I__8665 (
            .O(N__39583),
            .I(N__39570));
    Span4Mux_v I__8664 (
            .O(N__39580),
            .I(N__39567));
    InMux I__8663 (
            .O(N__39579),
            .I(N__39564));
    Odrv4 I__8662 (
            .O(N__39576),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__8661 (
            .O(N__39573),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__8660 (
            .O(N__39570),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    Odrv4 I__8659 (
            .O(N__39567),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__8658 (
            .O(N__39564),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    InMux I__8657 (
            .O(N__39553),
            .I(N__39550));
    LocalMux I__8656 (
            .O(N__39550),
            .I(N__39546));
    InMux I__8655 (
            .O(N__39549),
            .I(N__39542));
    Span4Mux_h I__8654 (
            .O(N__39546),
            .I(N__39539));
    InMux I__8653 (
            .O(N__39545),
            .I(N__39536));
    LocalMux I__8652 (
            .O(N__39542),
            .I(N__39533));
    Span4Mux_h I__8651 (
            .O(N__39539),
            .I(N__39530));
    LocalMux I__8650 (
            .O(N__39536),
            .I(N__39525));
    Span4Mux_v I__8649 (
            .O(N__39533),
            .I(N__39525));
    Odrv4 I__8648 (
            .O(N__39530),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    Odrv4 I__8647 (
            .O(N__39525),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    CEMux I__8646 (
            .O(N__39520),
            .I(N__39517));
    LocalMux I__8645 (
            .O(N__39517),
            .I(N__39514));
    Span4Mux_v I__8644 (
            .O(N__39514),
            .I(N__39511));
    Span4Mux_h I__8643 (
            .O(N__39511),
            .I(N__39508));
    Odrv4 I__8642 (
            .O(N__39508),
            .I(\phase_controller_inst1.N_221_0 ));
    CascadeMux I__8641 (
            .O(N__39505),
            .I(\delay_measurement_inst.delay_tr_timer.N_424_cascade_ ));
    InMux I__8640 (
            .O(N__39502),
            .I(N__39499));
    LocalMux I__8639 (
            .O(N__39499),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ));
    InMux I__8638 (
            .O(N__39496),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__8637 (
            .O(N__39493),
            .I(N__39490));
    LocalMux I__8636 (
            .O(N__39490),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ));
    InMux I__8635 (
            .O(N__39487),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__8634 (
            .O(N__39484),
            .I(N__39481));
    LocalMux I__8633 (
            .O(N__39481),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ));
    InMux I__8632 (
            .O(N__39478),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__8631 (
            .O(N__39475),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__8630 (
            .O(N__39472),
            .I(N__39469));
    LocalMux I__8629 (
            .O(N__39469),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ));
    InMux I__8628 (
            .O(N__39466),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__8627 (
            .O(N__39463),
            .I(N__39460));
    LocalMux I__8626 (
            .O(N__39460),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ));
    InMux I__8625 (
            .O(N__39457),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__8624 (
            .O(N__39454),
            .I(N__39451));
    LocalMux I__8623 (
            .O(N__39451),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ));
    InMux I__8622 (
            .O(N__39448),
            .I(bfn_16_18_0_));
    InMux I__8621 (
            .O(N__39445),
            .I(N__39442));
    LocalMux I__8620 (
            .O(N__39442),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ));
    InMux I__8619 (
            .O(N__39439),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__8618 (
            .O(N__39436),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__8617 (
            .O(N__39433),
            .I(N__39430));
    LocalMux I__8616 (
            .O(N__39430),
            .I(N__39427));
    Odrv4 I__8615 (
            .O(N__39427),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ));
    InMux I__8614 (
            .O(N__39424),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__8613 (
            .O(N__39421),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__8612 (
            .O(N__39418),
            .I(N__39415));
    LocalMux I__8611 (
            .O(N__39415),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ));
    InMux I__8610 (
            .O(N__39412),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__8609 (
            .O(N__39409),
            .I(N__39406));
    LocalMux I__8608 (
            .O(N__39406),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ));
    InMux I__8607 (
            .O(N__39403),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__8606 (
            .O(N__39400),
            .I(N__39397));
    LocalMux I__8605 (
            .O(N__39397),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ));
    InMux I__8604 (
            .O(N__39394),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__8603 (
            .O(N__39391),
            .I(N__39388));
    LocalMux I__8602 (
            .O(N__39388),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ));
    InMux I__8601 (
            .O(N__39385),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__8600 (
            .O(N__39382),
            .I(N__39379));
    LocalMux I__8599 (
            .O(N__39379),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ));
    InMux I__8598 (
            .O(N__39376),
            .I(bfn_16_17_0_));
    InMux I__8597 (
            .O(N__39373),
            .I(N__39370));
    LocalMux I__8596 (
            .O(N__39370),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ));
    InMux I__8595 (
            .O(N__39367),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__8594 (
            .O(N__39364),
            .I(N__39361));
    LocalMux I__8593 (
            .O(N__39361),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ));
    InMux I__8592 (
            .O(N__39358),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__8591 (
            .O(N__39355),
            .I(N__39352));
    LocalMux I__8590 (
            .O(N__39352),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ));
    InMux I__8589 (
            .O(N__39349),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__8588 (
            .O(N__39346),
            .I(N__39343));
    LocalMux I__8587 (
            .O(N__39343),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ));
    InMux I__8586 (
            .O(N__39340),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__8585 (
            .O(N__39337),
            .I(N__39334));
    LocalMux I__8584 (
            .O(N__39334),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ));
    InMux I__8583 (
            .O(N__39331),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__8582 (
            .O(N__39328),
            .I(N__39325));
    LocalMux I__8581 (
            .O(N__39325),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ));
    InMux I__8580 (
            .O(N__39322),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__8579 (
            .O(N__39319),
            .I(N__39316));
    LocalMux I__8578 (
            .O(N__39316),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ));
    InMux I__8577 (
            .O(N__39313),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__8576 (
            .O(N__39310),
            .I(N__39307));
    LocalMux I__8575 (
            .O(N__39307),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ));
    InMux I__8574 (
            .O(N__39304),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__8573 (
            .O(N__39301),
            .I(N__39298));
    LocalMux I__8572 (
            .O(N__39298),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ));
    InMux I__8571 (
            .O(N__39295),
            .I(bfn_16_16_0_));
    InMux I__8570 (
            .O(N__39292),
            .I(N__39289));
    LocalMux I__8569 (
            .O(N__39289),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ));
    InMux I__8568 (
            .O(N__39286),
            .I(N__39283));
    LocalMux I__8567 (
            .O(N__39283),
            .I(N__39280));
    Span4Mux_v I__8566 (
            .O(N__39280),
            .I(N__39276));
    InMux I__8565 (
            .O(N__39279),
            .I(N__39273));
    Odrv4 I__8564 (
            .O(N__39276),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ));
    LocalMux I__8563 (
            .O(N__39273),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ));
    CascadeMux I__8562 (
            .O(N__39268),
            .I(N__39265));
    InMux I__8561 (
            .O(N__39265),
            .I(N__39262));
    LocalMux I__8560 (
            .O(N__39262),
            .I(N__39258));
    CascadeMux I__8559 (
            .O(N__39261),
            .I(N__39255));
    Span4Mux_h I__8558 (
            .O(N__39258),
            .I(N__39252));
    InMux I__8557 (
            .O(N__39255),
            .I(N__39249));
    Odrv4 I__8556 (
            .O(N__39252),
            .I(measured_delay_tr_1));
    LocalMux I__8555 (
            .O(N__39249),
            .I(measured_delay_tr_1));
    CascadeMux I__8554 (
            .O(N__39244),
            .I(N__39241));
    InMux I__8553 (
            .O(N__39241),
            .I(N__39238));
    LocalMux I__8552 (
            .O(N__39238),
            .I(N__39235));
    Odrv4 I__8551 (
            .O(N__39235),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__8550 (
            .O(N__39232),
            .I(N__39229));
    InMux I__8549 (
            .O(N__39229),
            .I(N__39226));
    LocalMux I__8548 (
            .O(N__39226),
            .I(N__39223));
    Odrv4 I__8547 (
            .O(N__39223),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__8546 (
            .O(N__39220),
            .I(N__39216));
    CascadeMux I__8545 (
            .O(N__39219),
            .I(N__39211));
    InMux I__8544 (
            .O(N__39216),
            .I(N__39208));
    InMux I__8543 (
            .O(N__39215),
            .I(N__39205));
    InMux I__8542 (
            .O(N__39214),
            .I(N__39200));
    InMux I__8541 (
            .O(N__39211),
            .I(N__39200));
    LocalMux I__8540 (
            .O(N__39208),
            .I(N__39197));
    LocalMux I__8539 (
            .O(N__39205),
            .I(N__39192));
    LocalMux I__8538 (
            .O(N__39200),
            .I(N__39192));
    Span4Mux_v I__8537 (
            .O(N__39197),
            .I(N__39189));
    Span4Mux_v I__8536 (
            .O(N__39192),
            .I(N__39186));
    Odrv4 I__8535 (
            .O(N__39189),
            .I(measured_delay_tr_9));
    Odrv4 I__8534 (
            .O(N__39186),
            .I(measured_delay_tr_9));
    InMux I__8533 (
            .O(N__39181),
            .I(N__39178));
    LocalMux I__8532 (
            .O(N__39178),
            .I(N__39175));
    Span4Mux_v I__8531 (
            .O(N__39175),
            .I(N__39172));
    Span4Mux_h I__8530 (
            .O(N__39172),
            .I(N__39169));
    Odrv4 I__8529 (
            .O(N__39169),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3 ));
    InMux I__8528 (
            .O(N__39166),
            .I(N__39161));
    InMux I__8527 (
            .O(N__39165),
            .I(N__39156));
    InMux I__8526 (
            .O(N__39164),
            .I(N__39156));
    LocalMux I__8525 (
            .O(N__39161),
            .I(N__39151));
    LocalMux I__8524 (
            .O(N__39156),
            .I(N__39151));
    Span4Mux_v I__8523 (
            .O(N__39151),
            .I(N__39147));
    CascadeMux I__8522 (
            .O(N__39150),
            .I(N__39143));
    Span4Mux_h I__8521 (
            .O(N__39147),
            .I(N__39140));
    InMux I__8520 (
            .O(N__39146),
            .I(N__39135));
    InMux I__8519 (
            .O(N__39143),
            .I(N__39135));
    Odrv4 I__8518 (
            .O(N__39140),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ));
    LocalMux I__8517 (
            .O(N__39135),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ));
    InMux I__8516 (
            .O(N__39130),
            .I(N__39124));
    InMux I__8515 (
            .O(N__39129),
            .I(N__39124));
    LocalMux I__8514 (
            .O(N__39124),
            .I(N__39119));
    InMux I__8513 (
            .O(N__39123),
            .I(N__39116));
    CascadeMux I__8512 (
            .O(N__39122),
            .I(N__39113));
    Span4Mux_v I__8511 (
            .O(N__39119),
            .I(N__39107));
    LocalMux I__8510 (
            .O(N__39116),
            .I(N__39107));
    InMux I__8509 (
            .O(N__39113),
            .I(N__39102));
    InMux I__8508 (
            .O(N__39112),
            .I(N__39102));
    Span4Mux_h I__8507 (
            .O(N__39107),
            .I(N__39099));
    LocalMux I__8506 (
            .O(N__39102),
            .I(measured_delay_tr_3));
    Odrv4 I__8505 (
            .O(N__39099),
            .I(measured_delay_tr_3));
    CascadeMux I__8504 (
            .O(N__39094),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_ ));
    InMux I__8503 (
            .O(N__39091),
            .I(N__39082));
    InMux I__8502 (
            .O(N__39090),
            .I(N__39082));
    InMux I__8501 (
            .O(N__39089),
            .I(N__39082));
    LocalMux I__8500 (
            .O(N__39082),
            .I(N__39076));
    InMux I__8499 (
            .O(N__39081),
            .I(N__39069));
    InMux I__8498 (
            .O(N__39080),
            .I(N__39069));
    InMux I__8497 (
            .O(N__39079),
            .I(N__39069));
    Span12Mux_h I__8496 (
            .O(N__39076),
            .I(N__39066));
    LocalMux I__8495 (
            .O(N__39069),
            .I(N__39063));
    Odrv12 I__8494 (
            .O(N__39066),
            .I(\phase_controller_inst1.stoper_tr.N_20_li ));
    Odrv12 I__8493 (
            .O(N__39063),
            .I(\phase_controller_inst1.stoper_tr.N_20_li ));
    CascadeMux I__8492 (
            .O(N__39058),
            .I(N__39055));
    InMux I__8491 (
            .O(N__39055),
            .I(N__39052));
    LocalMux I__8490 (
            .O(N__39052),
            .I(N__39049));
    Odrv12 I__8489 (
            .O(N__39049),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ));
    InMux I__8488 (
            .O(N__39046),
            .I(N__39042));
    InMux I__8487 (
            .O(N__39045),
            .I(N__39039));
    LocalMux I__8486 (
            .O(N__39042),
            .I(N__39034));
    LocalMux I__8485 (
            .O(N__39039),
            .I(N__39031));
    CascadeMux I__8484 (
            .O(N__39038),
            .I(N__39028));
    InMux I__8483 (
            .O(N__39037),
            .I(N__39025));
    Span4Mux_v I__8482 (
            .O(N__39034),
            .I(N__39022));
    Span4Mux_h I__8481 (
            .O(N__39031),
            .I(N__39019));
    InMux I__8480 (
            .O(N__39028),
            .I(N__39016));
    LocalMux I__8479 (
            .O(N__39025),
            .I(N__39011));
    Span4Mux_h I__8478 (
            .O(N__39022),
            .I(N__39011));
    Odrv4 I__8477 (
            .O(N__39019),
            .I(measured_delay_tr_8));
    LocalMux I__8476 (
            .O(N__39016),
            .I(measured_delay_tr_8));
    Odrv4 I__8475 (
            .O(N__39011),
            .I(measured_delay_tr_8));
    InMux I__8474 (
            .O(N__39004),
            .I(N__38999));
    InMux I__8473 (
            .O(N__39003),
            .I(N__38995));
    InMux I__8472 (
            .O(N__39002),
            .I(N__38992));
    LocalMux I__8471 (
            .O(N__38999),
            .I(N__38989));
    CascadeMux I__8470 (
            .O(N__38998),
            .I(N__38986));
    LocalMux I__8469 (
            .O(N__38995),
            .I(N__38983));
    LocalMux I__8468 (
            .O(N__38992),
            .I(N__38980));
    Span4Mux_v I__8467 (
            .O(N__38989),
            .I(N__38977));
    InMux I__8466 (
            .O(N__38986),
            .I(N__38974));
    Span4Mux_v I__8465 (
            .O(N__38983),
            .I(N__38969));
    Span4Mux_h I__8464 (
            .O(N__38980),
            .I(N__38969));
    Odrv4 I__8463 (
            .O(N__38977),
            .I(measured_delay_tr_7));
    LocalMux I__8462 (
            .O(N__38974),
            .I(measured_delay_tr_7));
    Odrv4 I__8461 (
            .O(N__38969),
            .I(measured_delay_tr_7));
    InMux I__8460 (
            .O(N__38962),
            .I(N__38959));
    LocalMux I__8459 (
            .O(N__38959),
            .I(N__38956));
    Span4Mux_v I__8458 (
            .O(N__38956),
            .I(N__38951));
    InMux I__8457 (
            .O(N__38955),
            .I(N__38948));
    InMux I__8456 (
            .O(N__38954),
            .I(N__38945));
    Span4Mux_h I__8455 (
            .O(N__38951),
            .I(N__38942));
    LocalMux I__8454 (
            .O(N__38948),
            .I(N__38937));
    LocalMux I__8453 (
            .O(N__38945),
            .I(N__38937));
    Sp12to4 I__8452 (
            .O(N__38942),
            .I(N__38934));
    Span4Mux_v I__8451 (
            .O(N__38937),
            .I(N__38931));
    Odrv12 I__8450 (
            .O(N__38934),
            .I(measured_delay_tr_6));
    Odrv4 I__8449 (
            .O(N__38931),
            .I(measured_delay_tr_6));
    CascadeMux I__8448 (
            .O(N__38926),
            .I(N__38923));
    InMux I__8447 (
            .O(N__38923),
            .I(N__38920));
    LocalMux I__8446 (
            .O(N__38920),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6 ));
    CascadeMux I__8445 (
            .O(N__38917),
            .I(N__38914));
    InMux I__8444 (
            .O(N__38914),
            .I(N__38909));
    InMux I__8443 (
            .O(N__38913),
            .I(N__38906));
    CascadeMux I__8442 (
            .O(N__38912),
            .I(N__38903));
    LocalMux I__8441 (
            .O(N__38909),
            .I(N__38898));
    LocalMux I__8440 (
            .O(N__38906),
            .I(N__38898));
    InMux I__8439 (
            .O(N__38903),
            .I(N__38893));
    Span4Mux_v I__8438 (
            .O(N__38898),
            .I(N__38890));
    InMux I__8437 (
            .O(N__38897),
            .I(N__38885));
    InMux I__8436 (
            .O(N__38896),
            .I(N__38885));
    LocalMux I__8435 (
            .O(N__38893),
            .I(N__38876));
    Span4Mux_h I__8434 (
            .O(N__38890),
            .I(N__38876));
    LocalMux I__8433 (
            .O(N__38885),
            .I(N__38876));
    InMux I__8432 (
            .O(N__38884),
            .I(N__38873));
    CascadeMux I__8431 (
            .O(N__38883),
            .I(N__38870));
    Span4Mux_h I__8430 (
            .O(N__38876),
            .I(N__38864));
    LocalMux I__8429 (
            .O(N__38873),
            .I(N__38861));
    InMux I__8428 (
            .O(N__38870),
            .I(N__38858));
    InMux I__8427 (
            .O(N__38869),
            .I(N__38851));
    InMux I__8426 (
            .O(N__38868),
            .I(N__38851));
    InMux I__8425 (
            .O(N__38867),
            .I(N__38851));
    Span4Mux_v I__8424 (
            .O(N__38864),
            .I(N__38848));
    Span4Mux_h I__8423 (
            .O(N__38861),
            .I(N__38845));
    LocalMux I__8422 (
            .O(N__38858),
            .I(measured_delay_tr_15));
    LocalMux I__8421 (
            .O(N__38851),
            .I(measured_delay_tr_15));
    Odrv4 I__8420 (
            .O(N__38848),
            .I(measured_delay_tr_15));
    Odrv4 I__8419 (
            .O(N__38845),
            .I(measured_delay_tr_15));
    CascadeMux I__8418 (
            .O(N__38836),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_ ));
    InMux I__8417 (
            .O(N__38833),
            .I(N__38830));
    LocalMux I__8416 (
            .O(N__38830),
            .I(N__38827));
    Span4Mux_h I__8415 (
            .O(N__38827),
            .I(N__38820));
    InMux I__8414 (
            .O(N__38826),
            .I(N__38815));
    InMux I__8413 (
            .O(N__38825),
            .I(N__38815));
    InMux I__8412 (
            .O(N__38824),
            .I(N__38810));
    InMux I__8411 (
            .O(N__38823),
            .I(N__38810));
    Span4Mux_v I__8410 (
            .O(N__38820),
            .I(N__38805));
    LocalMux I__8409 (
            .O(N__38815),
            .I(N__38805));
    LocalMux I__8408 (
            .O(N__38810),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ));
    Odrv4 I__8407 (
            .O(N__38805),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ));
    InMux I__8406 (
            .O(N__38800),
            .I(N__38795));
    CascadeMux I__8405 (
            .O(N__38799),
            .I(N__38792));
    CascadeMux I__8404 (
            .O(N__38798),
            .I(N__38789));
    LocalMux I__8403 (
            .O(N__38795),
            .I(N__38786));
    InMux I__8402 (
            .O(N__38792),
            .I(N__38783));
    InMux I__8401 (
            .O(N__38789),
            .I(N__38780));
    Span4Mux_v I__8400 (
            .O(N__38786),
            .I(N__38777));
    LocalMux I__8399 (
            .O(N__38783),
            .I(N__38772));
    LocalMux I__8398 (
            .O(N__38780),
            .I(N__38772));
    Span4Mux_h I__8397 (
            .O(N__38777),
            .I(N__38769));
    Span4Mux_h I__8396 (
            .O(N__38772),
            .I(N__38766));
    Odrv4 I__8395 (
            .O(N__38769),
            .I(measured_delay_tr_5));
    Odrv4 I__8394 (
            .O(N__38766),
            .I(measured_delay_tr_5));
    CascadeMux I__8393 (
            .O(N__38761),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_ ));
    CascadeMux I__8392 (
            .O(N__38758),
            .I(N__38755));
    InMux I__8391 (
            .O(N__38755),
            .I(N__38752));
    LocalMux I__8390 (
            .O(N__38752),
            .I(N__38749));
    Span4Mux_h I__8389 (
            .O(N__38749),
            .I(N__38746));
    Odrv4 I__8388 (
            .O(N__38746),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ));
    InMux I__8387 (
            .O(N__38743),
            .I(N__38740));
    LocalMux I__8386 (
            .O(N__38740),
            .I(N__38737));
    Odrv12 I__8385 (
            .O(N__38737),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ));
    InMux I__8384 (
            .O(N__38734),
            .I(N__38730));
    InMux I__8383 (
            .O(N__38733),
            .I(N__38727));
    LocalMux I__8382 (
            .O(N__38730),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__8381 (
            .O(N__38727),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__8380 (
            .O(N__38722),
            .I(N__38719));
    InMux I__8379 (
            .O(N__38719),
            .I(N__38716));
    LocalMux I__8378 (
            .O(N__38716),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ));
    InMux I__8377 (
            .O(N__38713),
            .I(N__38709));
    InMux I__8376 (
            .O(N__38712),
            .I(N__38706));
    LocalMux I__8375 (
            .O(N__38709),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__8374 (
            .O(N__38706),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__8373 (
            .O(N__38701),
            .I(N__38698));
    LocalMux I__8372 (
            .O(N__38698),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ));
    CascadeMux I__8371 (
            .O(N__38695),
            .I(N__38692));
    InMux I__8370 (
            .O(N__38692),
            .I(N__38688));
    InMux I__8369 (
            .O(N__38691),
            .I(N__38685));
    LocalMux I__8368 (
            .O(N__38688),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__8367 (
            .O(N__38685),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__8366 (
            .O(N__38680),
            .I(N__38677));
    LocalMux I__8365 (
            .O(N__38677),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ));
    InMux I__8364 (
            .O(N__38674),
            .I(N__38670));
    InMux I__8363 (
            .O(N__38673),
            .I(N__38667));
    LocalMux I__8362 (
            .O(N__38670),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__8361 (
            .O(N__38667),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__8360 (
            .O(N__38662),
            .I(N__38659));
    LocalMux I__8359 (
            .O(N__38659),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ));
    InMux I__8358 (
            .O(N__38656),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__8357 (
            .O(N__38653),
            .I(N__38650));
    InMux I__8356 (
            .O(N__38650),
            .I(N__38647));
    LocalMux I__8355 (
            .O(N__38647),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__8354 (
            .O(N__38644),
            .I(N__38641));
    InMux I__8353 (
            .O(N__38641),
            .I(N__38638));
    LocalMux I__8352 (
            .O(N__38638),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__8351 (
            .O(N__38635),
            .I(N__38632));
    InMux I__8350 (
            .O(N__38632),
            .I(N__38629));
    LocalMux I__8349 (
            .O(N__38629),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ));
    InMux I__8348 (
            .O(N__38626),
            .I(N__38623));
    LocalMux I__8347 (
            .O(N__38623),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__8346 (
            .O(N__38620),
            .I(N__38617));
    InMux I__8345 (
            .O(N__38617),
            .I(N__38614));
    LocalMux I__8344 (
            .O(N__38614),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ));
    InMux I__8343 (
            .O(N__38611),
            .I(N__38607));
    InMux I__8342 (
            .O(N__38610),
            .I(N__38604));
    LocalMux I__8341 (
            .O(N__38607),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__8340 (
            .O(N__38604),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__8339 (
            .O(N__38599),
            .I(N__38596));
    LocalMux I__8338 (
            .O(N__38596),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__8337 (
            .O(N__38593),
            .I(N__38590));
    InMux I__8336 (
            .O(N__38590),
            .I(N__38587));
    LocalMux I__8335 (
            .O(N__38587),
            .I(N__38584));
    Odrv4 I__8334 (
            .O(N__38584),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__8333 (
            .O(N__38581),
            .I(N__38578));
    InMux I__8332 (
            .O(N__38578),
            .I(N__38574));
    InMux I__8331 (
            .O(N__38577),
            .I(N__38571));
    LocalMux I__8330 (
            .O(N__38574),
            .I(N__38568));
    LocalMux I__8329 (
            .O(N__38571),
            .I(N__38565));
    Odrv4 I__8328 (
            .O(N__38568),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__8327 (
            .O(N__38565),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__8326 (
            .O(N__38560),
            .I(N__38557));
    LocalMux I__8325 (
            .O(N__38557),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__8324 (
            .O(N__38554),
            .I(N__38551));
    InMux I__8323 (
            .O(N__38551),
            .I(N__38548));
    LocalMux I__8322 (
            .O(N__38548),
            .I(N__38545));
    Odrv4 I__8321 (
            .O(N__38545),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ));
    InMux I__8320 (
            .O(N__38542),
            .I(N__38539));
    LocalMux I__8319 (
            .O(N__38539),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__8318 (
            .O(N__38536),
            .I(N__38533));
    InMux I__8317 (
            .O(N__38533),
            .I(N__38530));
    LocalMux I__8316 (
            .O(N__38530),
            .I(N__38527));
    Odrv4 I__8315 (
            .O(N__38527),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ));
    InMux I__8314 (
            .O(N__38524),
            .I(N__38520));
    InMux I__8313 (
            .O(N__38523),
            .I(N__38517));
    LocalMux I__8312 (
            .O(N__38520),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__8311 (
            .O(N__38517),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__8310 (
            .O(N__38512),
            .I(N__38509));
    LocalMux I__8309 (
            .O(N__38509),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__8308 (
            .O(N__38506),
            .I(N__38503));
    InMux I__8307 (
            .O(N__38503),
            .I(N__38499));
    InMux I__8306 (
            .O(N__38502),
            .I(N__38496));
    LocalMux I__8305 (
            .O(N__38499),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__8304 (
            .O(N__38496),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__8303 (
            .O(N__38491),
            .I(N__38488));
    InMux I__8302 (
            .O(N__38488),
            .I(N__38485));
    LocalMux I__8301 (
            .O(N__38485),
            .I(N__38482));
    Span4Mux_v I__8300 (
            .O(N__38482),
            .I(N__38479));
    Odrv4 I__8299 (
            .O(N__38479),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ));
    InMux I__8298 (
            .O(N__38476),
            .I(N__38473));
    LocalMux I__8297 (
            .O(N__38473),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__8296 (
            .O(N__38470),
            .I(N__38467));
    InMux I__8295 (
            .O(N__38467),
            .I(N__38464));
    LocalMux I__8294 (
            .O(N__38464),
            .I(N__38461));
    Odrv4 I__8293 (
            .O(N__38461),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ));
    InMux I__8292 (
            .O(N__38458),
            .I(N__38454));
    InMux I__8291 (
            .O(N__38457),
            .I(N__38451));
    LocalMux I__8290 (
            .O(N__38454),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__8289 (
            .O(N__38451),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__8288 (
            .O(N__38446),
            .I(N__38443));
    LocalMux I__8287 (
            .O(N__38443),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__8286 (
            .O(N__38440),
            .I(N__38437));
    InMux I__8285 (
            .O(N__38437),
            .I(N__38434));
    LocalMux I__8284 (
            .O(N__38434),
            .I(N__38431));
    Span4Mux_v I__8283 (
            .O(N__38431),
            .I(N__38428));
    Odrv4 I__8282 (
            .O(N__38428),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ));
    InMux I__8281 (
            .O(N__38425),
            .I(N__38421));
    InMux I__8280 (
            .O(N__38424),
            .I(N__38418));
    LocalMux I__8279 (
            .O(N__38421),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__8278 (
            .O(N__38418),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__8277 (
            .O(N__38413),
            .I(N__38410));
    LocalMux I__8276 (
            .O(N__38410),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__8275 (
            .O(N__38407),
            .I(N__38403));
    InMux I__8274 (
            .O(N__38406),
            .I(N__38399));
    InMux I__8273 (
            .O(N__38403),
            .I(N__38396));
    InMux I__8272 (
            .O(N__38402),
            .I(N__38393));
    LocalMux I__8271 (
            .O(N__38399),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__8270 (
            .O(N__38396),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__8269 (
            .O(N__38393),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__8268 (
            .O(N__38386),
            .I(N__38383));
    LocalMux I__8267 (
            .O(N__38383),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ));
    InMux I__8266 (
            .O(N__38380),
            .I(N__38376));
    InMux I__8265 (
            .O(N__38379),
            .I(N__38373));
    LocalMux I__8264 (
            .O(N__38376),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__8263 (
            .O(N__38373),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__8262 (
            .O(N__38368),
            .I(N__38365));
    LocalMux I__8261 (
            .O(N__38365),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__8260 (
            .O(N__38362),
            .I(N__38359));
    InMux I__8259 (
            .O(N__38359),
            .I(N__38355));
    InMux I__8258 (
            .O(N__38358),
            .I(N__38352));
    LocalMux I__8257 (
            .O(N__38355),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__8256 (
            .O(N__38352),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__8255 (
            .O(N__38347),
            .I(N__38344));
    LocalMux I__8254 (
            .O(N__38344),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__8253 (
            .O(N__38341),
            .I(N__38338));
    InMux I__8252 (
            .O(N__38338),
            .I(N__38335));
    LocalMux I__8251 (
            .O(N__38335),
            .I(N__38332));
    Odrv4 I__8250 (
            .O(N__38332),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ));
    InMux I__8249 (
            .O(N__38329),
            .I(N__38325));
    InMux I__8248 (
            .O(N__38328),
            .I(N__38322));
    LocalMux I__8247 (
            .O(N__38325),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__8246 (
            .O(N__38322),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__8245 (
            .O(N__38317),
            .I(N__38314));
    LocalMux I__8244 (
            .O(N__38314),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ));
    InMux I__8243 (
            .O(N__38311),
            .I(N__38307));
    InMux I__8242 (
            .O(N__38310),
            .I(N__38304));
    LocalMux I__8241 (
            .O(N__38307),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__8240 (
            .O(N__38304),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__8239 (
            .O(N__38299),
            .I(N__38296));
    LocalMux I__8238 (
            .O(N__38296),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__8237 (
            .O(N__38293),
            .I(N__38290));
    InMux I__8236 (
            .O(N__38290),
            .I(N__38287));
    LocalMux I__8235 (
            .O(N__38287),
            .I(N__38284));
    Odrv4 I__8234 (
            .O(N__38284),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ));
    InMux I__8233 (
            .O(N__38281),
            .I(N__38277));
    InMux I__8232 (
            .O(N__38280),
            .I(N__38274));
    LocalMux I__8231 (
            .O(N__38277),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__8230 (
            .O(N__38274),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__8229 (
            .O(N__38269),
            .I(N__38266));
    LocalMux I__8228 (
            .O(N__38266),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__8227 (
            .O(N__38263),
            .I(N__38260));
    InMux I__8226 (
            .O(N__38260),
            .I(N__38257));
    LocalMux I__8225 (
            .O(N__38257),
            .I(N__38254));
    Odrv4 I__8224 (
            .O(N__38254),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ));
    InMux I__8223 (
            .O(N__38251),
            .I(N__38247));
    InMux I__8222 (
            .O(N__38250),
            .I(N__38244));
    LocalMux I__8221 (
            .O(N__38247),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__8220 (
            .O(N__38244),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__8219 (
            .O(N__38239),
            .I(N__38236));
    LocalMux I__8218 (
            .O(N__38236),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__8217 (
            .O(N__38233),
            .I(N__38230));
    InMux I__8216 (
            .O(N__38230),
            .I(N__38227));
    LocalMux I__8215 (
            .O(N__38227),
            .I(N__38224));
    Span4Mux_h I__8214 (
            .O(N__38224),
            .I(N__38221));
    Odrv4 I__8213 (
            .O(N__38221),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ));
    InMux I__8212 (
            .O(N__38218),
            .I(N__38214));
    InMux I__8211 (
            .O(N__38217),
            .I(N__38211));
    LocalMux I__8210 (
            .O(N__38214),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__8209 (
            .O(N__38211),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__8208 (
            .O(N__38206),
            .I(N__38203));
    InMux I__8207 (
            .O(N__38203),
            .I(N__38200));
    LocalMux I__8206 (
            .O(N__38200),
            .I(N__38197));
    Odrv4 I__8205 (
            .O(N__38197),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ));
    InMux I__8204 (
            .O(N__38194),
            .I(N__38191));
    LocalMux I__8203 (
            .O(N__38191),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__8202 (
            .O(N__38188),
            .I(N__38185));
    InMux I__8201 (
            .O(N__38185),
            .I(N__38182));
    LocalMux I__8200 (
            .O(N__38182),
            .I(N__38179));
    Odrv12 I__8199 (
            .O(N__38179),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ));
    InMux I__8198 (
            .O(N__38176),
            .I(N__38173));
    LocalMux I__8197 (
            .O(N__38173),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ));
    CascadeMux I__8196 (
            .O(N__38170),
            .I(N__38167));
    InMux I__8195 (
            .O(N__38167),
            .I(N__38164));
    LocalMux I__8194 (
            .O(N__38164),
            .I(N__38161));
    Odrv4 I__8193 (
            .O(N__38161),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ));
    InMux I__8192 (
            .O(N__38158),
            .I(N__38155));
    LocalMux I__8191 (
            .O(N__38155),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ));
    CascadeMux I__8190 (
            .O(N__38152),
            .I(N__38149));
    InMux I__8189 (
            .O(N__38149),
            .I(N__38146));
    LocalMux I__8188 (
            .O(N__38146),
            .I(N__38143));
    Odrv4 I__8187 (
            .O(N__38143),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ));
    InMux I__8186 (
            .O(N__38140),
            .I(N__38137));
    LocalMux I__8185 (
            .O(N__38137),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ));
    CascadeMux I__8184 (
            .O(N__38134),
            .I(N__38131));
    InMux I__8183 (
            .O(N__38131),
            .I(N__38128));
    LocalMux I__8182 (
            .O(N__38128),
            .I(N__38125));
    Span4Mux_h I__8181 (
            .O(N__38125),
            .I(N__38122));
    Odrv4 I__8180 (
            .O(N__38122),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ));
    InMux I__8179 (
            .O(N__38119),
            .I(N__38116));
    LocalMux I__8178 (
            .O(N__38116),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ));
    InMux I__8177 (
            .O(N__38113),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__8176 (
            .O(N__38110),
            .I(N__38107));
    InMux I__8175 (
            .O(N__38107),
            .I(N__38104));
    LocalMux I__8174 (
            .O(N__38104),
            .I(N__38101));
    Odrv4 I__8173 (
            .O(N__38101),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ));
    InMux I__8172 (
            .O(N__38098),
            .I(N__38095));
    LocalMux I__8171 (
            .O(N__38095),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__8170 (
            .O(N__38092),
            .I(N__38089));
    InMux I__8169 (
            .O(N__38089),
            .I(N__38086));
    LocalMux I__8168 (
            .O(N__38086),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ));
    InMux I__8167 (
            .O(N__38083),
            .I(N__38080));
    LocalMux I__8166 (
            .O(N__38080),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__8165 (
            .O(N__38077),
            .I(N__38074));
    InMux I__8164 (
            .O(N__38074),
            .I(N__38071));
    LocalMux I__8163 (
            .O(N__38071),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ));
    InMux I__8162 (
            .O(N__38068),
            .I(N__38065));
    LocalMux I__8161 (
            .O(N__38065),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__8160 (
            .O(N__38062),
            .I(N__38059));
    InMux I__8159 (
            .O(N__38059),
            .I(N__38056));
    LocalMux I__8158 (
            .O(N__38056),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ));
    InMux I__8157 (
            .O(N__38053),
            .I(N__38050));
    LocalMux I__8156 (
            .O(N__38050),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__8155 (
            .O(N__38047),
            .I(N__38044));
    InMux I__8154 (
            .O(N__38044),
            .I(N__38041));
    LocalMux I__8153 (
            .O(N__38041),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ));
    InMux I__8152 (
            .O(N__38038),
            .I(N__38035));
    LocalMux I__8151 (
            .O(N__38035),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__8150 (
            .O(N__38032),
            .I(N__38029));
    InMux I__8149 (
            .O(N__38029),
            .I(N__38026));
    LocalMux I__8148 (
            .O(N__38026),
            .I(N__38023));
    Odrv12 I__8147 (
            .O(N__38023),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ));
    InMux I__8146 (
            .O(N__38020),
            .I(N__38017));
    LocalMux I__8145 (
            .O(N__38017),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__8144 (
            .O(N__38014),
            .I(N__38011));
    InMux I__8143 (
            .O(N__38011),
            .I(N__38008));
    LocalMux I__8142 (
            .O(N__38008),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ));
    InMux I__8141 (
            .O(N__38005),
            .I(N__38002));
    LocalMux I__8140 (
            .O(N__38002),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__8139 (
            .O(N__37999),
            .I(N__37996));
    InMux I__8138 (
            .O(N__37996),
            .I(N__37993));
    LocalMux I__8137 (
            .O(N__37993),
            .I(N__37990));
    Span4Mux_v I__8136 (
            .O(N__37990),
            .I(N__37987));
    Span4Mux_h I__8135 (
            .O(N__37987),
            .I(N__37984));
    Odrv4 I__8134 (
            .O(N__37984),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ));
    InMux I__8133 (
            .O(N__37981),
            .I(N__37978));
    LocalMux I__8132 (
            .O(N__37978),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ));
    InMux I__8131 (
            .O(N__37975),
            .I(N__37972));
    LocalMux I__8130 (
            .O(N__37972),
            .I(N__37969));
    Odrv4 I__8129 (
            .O(N__37969),
            .I(delay_hc_input_c));
    InMux I__8128 (
            .O(N__37966),
            .I(N__37963));
    LocalMux I__8127 (
            .O(N__37963),
            .I(N__37960));
    Odrv12 I__8126 (
            .O(N__37960),
            .I(delay_hc_d1));
    CascadeMux I__8125 (
            .O(N__37957),
            .I(N__37954));
    InMux I__8124 (
            .O(N__37954),
            .I(N__37951));
    LocalMux I__8123 (
            .O(N__37951),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_0 ));
    InMux I__8122 (
            .O(N__37948),
            .I(N__37945));
    LocalMux I__8121 (
            .O(N__37945),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__8120 (
            .O(N__37942),
            .I(N__37939));
    InMux I__8119 (
            .O(N__37939),
            .I(N__37936));
    LocalMux I__8118 (
            .O(N__37936),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__8117 (
            .O(N__37933),
            .I(N__37930));
    InMux I__8116 (
            .O(N__37930),
            .I(N__37927));
    LocalMux I__8115 (
            .O(N__37927),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ));
    InMux I__8114 (
            .O(N__37924),
            .I(N__37921));
    LocalMux I__8113 (
            .O(N__37921),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__8112 (
            .O(N__37918),
            .I(N__37915));
    InMux I__8111 (
            .O(N__37915),
            .I(N__37912));
    LocalMux I__8110 (
            .O(N__37912),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ));
    InMux I__8109 (
            .O(N__37909),
            .I(N__37906));
    LocalMux I__8108 (
            .O(N__37906),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__8107 (
            .O(N__37903),
            .I(N__37900));
    InMux I__8106 (
            .O(N__37900),
            .I(N__37897));
    LocalMux I__8105 (
            .O(N__37897),
            .I(N__37894));
    Odrv4 I__8104 (
            .O(N__37894),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ));
    InMux I__8103 (
            .O(N__37891),
            .I(N__37888));
    LocalMux I__8102 (
            .O(N__37888),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__8101 (
            .O(N__37885),
            .I(N__37882));
    InMux I__8100 (
            .O(N__37882),
            .I(N__37879));
    LocalMux I__8099 (
            .O(N__37879),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ));
    InMux I__8098 (
            .O(N__37876),
            .I(N__37873));
    LocalMux I__8097 (
            .O(N__37873),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__8096 (
            .O(N__37870),
            .I(N__37867));
    InMux I__8095 (
            .O(N__37867),
            .I(N__37864));
    LocalMux I__8094 (
            .O(N__37864),
            .I(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ));
    InMux I__8093 (
            .O(N__37861),
            .I(N__37858));
    LocalMux I__8092 (
            .O(N__37858),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__8091 (
            .O(N__37855),
            .I(N__37852));
    InMux I__8090 (
            .O(N__37852),
            .I(N__37849));
    LocalMux I__8089 (
            .O(N__37849),
            .I(N__37846));
    Span4Mux_v I__8088 (
            .O(N__37846),
            .I(N__37843));
    Odrv4 I__8087 (
            .O(N__37843),
            .I(\current_shift_inst.z_5_23 ));
    InMux I__8086 (
            .O(N__37840),
            .I(\current_shift_inst.z_5_cry_22 ));
    CascadeMux I__8085 (
            .O(N__37837),
            .I(N__37834));
    InMux I__8084 (
            .O(N__37834),
            .I(N__37831));
    LocalMux I__8083 (
            .O(N__37831),
            .I(N__37828));
    Span4Mux_h I__8082 (
            .O(N__37828),
            .I(N__37825));
    Odrv4 I__8081 (
            .O(N__37825),
            .I(\current_shift_inst.z_5_24 ));
    InMux I__8080 (
            .O(N__37822),
            .I(\current_shift_inst.z_5_cry_23 ));
    InMux I__8079 (
            .O(N__37819),
            .I(N__37816));
    LocalMux I__8078 (
            .O(N__37816),
            .I(N__37813));
    Span4Mux_v I__8077 (
            .O(N__37813),
            .I(N__37810));
    Odrv4 I__8076 (
            .O(N__37810),
            .I(\current_shift_inst.z_5_25 ));
    InMux I__8075 (
            .O(N__37807),
            .I(bfn_15_24_0_));
    CascadeMux I__8074 (
            .O(N__37804),
            .I(N__37801));
    InMux I__8073 (
            .O(N__37801),
            .I(N__37798));
    LocalMux I__8072 (
            .O(N__37798),
            .I(N__37795));
    Span4Mux_h I__8071 (
            .O(N__37795),
            .I(N__37792));
    Odrv4 I__8070 (
            .O(N__37792),
            .I(\current_shift_inst.z_5_26 ));
    InMux I__8069 (
            .O(N__37789),
            .I(\current_shift_inst.z_5_cry_25 ));
    CascadeMux I__8068 (
            .O(N__37786),
            .I(N__37783));
    InMux I__8067 (
            .O(N__37783),
            .I(N__37780));
    LocalMux I__8066 (
            .O(N__37780),
            .I(N__37777));
    Span4Mux_h I__8065 (
            .O(N__37777),
            .I(N__37774));
    Odrv4 I__8064 (
            .O(N__37774),
            .I(\current_shift_inst.z_5_27 ));
    InMux I__8063 (
            .O(N__37771),
            .I(\current_shift_inst.z_5_cry_26 ));
    InMux I__8062 (
            .O(N__37768),
            .I(N__37765));
    LocalMux I__8061 (
            .O(N__37765),
            .I(N__37762));
    Span4Mux_v I__8060 (
            .O(N__37762),
            .I(N__37759));
    Odrv4 I__8059 (
            .O(N__37759),
            .I(\current_shift_inst.z_5_28 ));
    InMux I__8058 (
            .O(N__37756),
            .I(\current_shift_inst.z_5_cry_27 ));
    CascadeMux I__8057 (
            .O(N__37753),
            .I(N__37750));
    InMux I__8056 (
            .O(N__37750),
            .I(N__37747));
    LocalMux I__8055 (
            .O(N__37747),
            .I(N__37744));
    Span4Mux_v I__8054 (
            .O(N__37744),
            .I(N__37741));
    Odrv4 I__8053 (
            .O(N__37741),
            .I(\current_shift_inst.z_5_29 ));
    InMux I__8052 (
            .O(N__37738),
            .I(\current_shift_inst.z_5_cry_28 ));
    InMux I__8051 (
            .O(N__37735),
            .I(N__37732));
    LocalMux I__8050 (
            .O(N__37732),
            .I(N__37729));
    Span4Mux_v I__8049 (
            .O(N__37729),
            .I(N__37726));
    Odrv4 I__8048 (
            .O(N__37726),
            .I(\current_shift_inst.z_5_30 ));
    InMux I__8047 (
            .O(N__37723),
            .I(\current_shift_inst.z_5_cry_29 ));
    InMux I__8046 (
            .O(N__37720),
            .I(\current_shift_inst.z_5_cry_30 ));
    InMux I__8045 (
            .O(N__37717),
            .I(N__37714));
    LocalMux I__8044 (
            .O(N__37714),
            .I(N__37711));
    Span4Mux_v I__8043 (
            .O(N__37711),
            .I(N__37708));
    Odrv4 I__8042 (
            .O(N__37708),
            .I(\current_shift_inst.z_5_cry_30_THRU_CO ));
    CascadeMux I__8041 (
            .O(N__37705),
            .I(N__37702));
    InMux I__8040 (
            .O(N__37702),
            .I(N__37699));
    LocalMux I__8039 (
            .O(N__37699),
            .I(N__37696));
    Span4Mux_v I__8038 (
            .O(N__37696),
            .I(N__37693));
    Odrv4 I__8037 (
            .O(N__37693),
            .I(\current_shift_inst.z_5_15 ));
    InMux I__8036 (
            .O(N__37690),
            .I(\current_shift_inst.z_5_cry_14 ));
    CascadeMux I__8035 (
            .O(N__37687),
            .I(N__37684));
    InMux I__8034 (
            .O(N__37684),
            .I(N__37681));
    LocalMux I__8033 (
            .O(N__37681),
            .I(N__37678));
    Span4Mux_h I__8032 (
            .O(N__37678),
            .I(N__37675));
    Odrv4 I__8031 (
            .O(N__37675),
            .I(\current_shift_inst.z_5_16 ));
    InMux I__8030 (
            .O(N__37672),
            .I(\current_shift_inst.z_5_cry_15 ));
    InMux I__8029 (
            .O(N__37669),
            .I(N__37666));
    LocalMux I__8028 (
            .O(N__37666),
            .I(N__37663));
    Span4Mux_v I__8027 (
            .O(N__37663),
            .I(N__37660));
    Odrv4 I__8026 (
            .O(N__37660),
            .I(\current_shift_inst.z_5_17 ));
    InMux I__8025 (
            .O(N__37657),
            .I(bfn_15_23_0_));
    CascadeMux I__8024 (
            .O(N__37654),
            .I(N__37651));
    InMux I__8023 (
            .O(N__37651),
            .I(N__37648));
    LocalMux I__8022 (
            .O(N__37648),
            .I(N__37645));
    Span4Mux_h I__8021 (
            .O(N__37645),
            .I(N__37642));
    Odrv4 I__8020 (
            .O(N__37642),
            .I(\current_shift_inst.z_5_18 ));
    InMux I__8019 (
            .O(N__37639),
            .I(\current_shift_inst.z_5_cry_17 ));
    InMux I__8018 (
            .O(N__37636),
            .I(N__37633));
    LocalMux I__8017 (
            .O(N__37633),
            .I(N__37630));
    Odrv4 I__8016 (
            .O(N__37630),
            .I(\current_shift_inst.z_5_19 ));
    InMux I__8015 (
            .O(N__37627),
            .I(\current_shift_inst.z_5_cry_18 ));
    InMux I__8014 (
            .O(N__37624),
            .I(N__37621));
    LocalMux I__8013 (
            .O(N__37621),
            .I(N__37618));
    Span4Mux_h I__8012 (
            .O(N__37618),
            .I(N__37615));
    Odrv4 I__8011 (
            .O(N__37615),
            .I(\current_shift_inst.z_5_20 ));
    InMux I__8010 (
            .O(N__37612),
            .I(\current_shift_inst.z_5_cry_19 ));
    InMux I__8009 (
            .O(N__37609),
            .I(N__37606));
    LocalMux I__8008 (
            .O(N__37606),
            .I(N__37603));
    Odrv4 I__8007 (
            .O(N__37603),
            .I(\current_shift_inst.z_5_21 ));
    InMux I__8006 (
            .O(N__37600),
            .I(\current_shift_inst.z_5_cry_20 ));
    InMux I__8005 (
            .O(N__37597),
            .I(N__37594));
    LocalMux I__8004 (
            .O(N__37594),
            .I(N__37591));
    Span4Mux_v I__8003 (
            .O(N__37591),
            .I(N__37588));
    Odrv4 I__8002 (
            .O(N__37588),
            .I(\current_shift_inst.z_5_22 ));
    InMux I__8001 (
            .O(N__37585),
            .I(\current_shift_inst.z_5_cry_21 ));
    CascadeMux I__8000 (
            .O(N__37582),
            .I(N__37579));
    InMux I__7999 (
            .O(N__37579),
            .I(N__37576));
    LocalMux I__7998 (
            .O(N__37576),
            .I(N__37573));
    Span4Mux_v I__7997 (
            .O(N__37573),
            .I(N__37570));
    Odrv4 I__7996 (
            .O(N__37570),
            .I(\current_shift_inst.z_5_7 ));
    InMux I__7995 (
            .O(N__37567),
            .I(\current_shift_inst.z_5_cry_6 ));
    InMux I__7994 (
            .O(N__37564),
            .I(N__37561));
    LocalMux I__7993 (
            .O(N__37561),
            .I(N__37558));
    Span4Mux_h I__7992 (
            .O(N__37558),
            .I(N__37555));
    Odrv4 I__7991 (
            .O(N__37555),
            .I(\current_shift_inst.z_5_8 ));
    InMux I__7990 (
            .O(N__37552),
            .I(\current_shift_inst.z_5_cry_7 ));
    CascadeMux I__7989 (
            .O(N__37549),
            .I(N__37546));
    InMux I__7988 (
            .O(N__37546),
            .I(N__37543));
    LocalMux I__7987 (
            .O(N__37543),
            .I(N__37540));
    Odrv4 I__7986 (
            .O(N__37540),
            .I(\current_shift_inst.z_5_9 ));
    InMux I__7985 (
            .O(N__37537),
            .I(bfn_15_22_0_));
    InMux I__7984 (
            .O(N__37534),
            .I(N__37531));
    LocalMux I__7983 (
            .O(N__37531),
            .I(N__37528));
    Odrv4 I__7982 (
            .O(N__37528),
            .I(\current_shift_inst.z_5_10 ));
    InMux I__7981 (
            .O(N__37525),
            .I(\current_shift_inst.z_5_cry_9 ));
    InMux I__7980 (
            .O(N__37522),
            .I(N__37519));
    LocalMux I__7979 (
            .O(N__37519),
            .I(N__37516));
    Odrv4 I__7978 (
            .O(N__37516),
            .I(\current_shift_inst.z_5_11 ));
    InMux I__7977 (
            .O(N__37513),
            .I(\current_shift_inst.z_5_cry_10 ));
    CascadeMux I__7976 (
            .O(N__37510),
            .I(N__37507));
    InMux I__7975 (
            .O(N__37507),
            .I(N__37504));
    LocalMux I__7974 (
            .O(N__37504),
            .I(N__37501));
    Odrv4 I__7973 (
            .O(N__37501),
            .I(\current_shift_inst.z_5_12 ));
    InMux I__7972 (
            .O(N__37498),
            .I(\current_shift_inst.z_5_cry_11 ));
    InMux I__7971 (
            .O(N__37495),
            .I(N__37492));
    LocalMux I__7970 (
            .O(N__37492),
            .I(N__37489));
    Odrv4 I__7969 (
            .O(N__37489),
            .I(\current_shift_inst.z_5_13 ));
    InMux I__7968 (
            .O(N__37486),
            .I(\current_shift_inst.z_5_cry_12 ));
    CascadeMux I__7967 (
            .O(N__37483),
            .I(N__37480));
    InMux I__7966 (
            .O(N__37480),
            .I(N__37477));
    LocalMux I__7965 (
            .O(N__37477),
            .I(N__37474));
    Span4Mux_v I__7964 (
            .O(N__37474),
            .I(N__37471));
    Odrv4 I__7963 (
            .O(N__37471),
            .I(\current_shift_inst.z_5_14 ));
    InMux I__7962 (
            .O(N__37468),
            .I(\current_shift_inst.z_5_cry_13 ));
    InMux I__7961 (
            .O(N__37465),
            .I(N__37462));
    LocalMux I__7960 (
            .O(N__37462),
            .I(N__37459));
    Span4Mux_h I__7959 (
            .O(N__37459),
            .I(N__37456));
    Span4Mux_h I__7958 (
            .O(N__37456),
            .I(N__37453));
    Odrv4 I__7957 (
            .O(N__37453),
            .I(\current_shift_inst.N_1742_i ));
    CascadeMux I__7956 (
            .O(N__37450),
            .I(N__37445));
    CascadeMux I__7955 (
            .O(N__37449),
            .I(N__37440));
    InMux I__7954 (
            .O(N__37448),
            .I(N__37437));
    InMux I__7953 (
            .O(N__37445),
            .I(N__37432));
    InMux I__7952 (
            .O(N__37444),
            .I(N__37432));
    CascadeMux I__7951 (
            .O(N__37443),
            .I(N__37428));
    InMux I__7950 (
            .O(N__37440),
            .I(N__37424));
    LocalMux I__7949 (
            .O(N__37437),
            .I(N__37421));
    LocalMux I__7948 (
            .O(N__37432),
            .I(N__37418));
    InMux I__7947 (
            .O(N__37431),
            .I(N__37413));
    InMux I__7946 (
            .O(N__37428),
            .I(N__37413));
    InMux I__7945 (
            .O(N__37427),
            .I(N__37410));
    LocalMux I__7944 (
            .O(N__37424),
            .I(N__37405));
    Span4Mux_v I__7943 (
            .O(N__37421),
            .I(N__37402));
    Span4Mux_v I__7942 (
            .O(N__37418),
            .I(N__37399));
    LocalMux I__7941 (
            .O(N__37413),
            .I(N__37394));
    LocalMux I__7940 (
            .O(N__37410),
            .I(N__37394));
    InMux I__7939 (
            .O(N__37409),
            .I(N__37391));
    InMux I__7938 (
            .O(N__37408),
            .I(N__37388));
    Span4Mux_v I__7937 (
            .O(N__37405),
            .I(N__37381));
    Span4Mux_h I__7936 (
            .O(N__37402),
            .I(N__37381));
    Span4Mux_h I__7935 (
            .O(N__37399),
            .I(N__37381));
    Span4Mux_v I__7934 (
            .O(N__37394),
            .I(N__37376));
    LocalMux I__7933 (
            .O(N__37391),
            .I(N__37376));
    LocalMux I__7932 (
            .O(N__37388),
            .I(N__37373));
    Span4Mux_v I__7931 (
            .O(N__37381),
            .I(N__37368));
    Span4Mux_v I__7930 (
            .O(N__37376),
            .I(N__37368));
    Odrv4 I__7929 (
            .O(N__37373),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__7928 (
            .O(N__37368),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__7927 (
            .O(N__37363),
            .I(N__37359));
    InMux I__7926 (
            .O(N__37362),
            .I(N__37356));
    InMux I__7925 (
            .O(N__37359),
            .I(N__37353));
    LocalMux I__7924 (
            .O(N__37356),
            .I(N__37350));
    LocalMux I__7923 (
            .O(N__37353),
            .I(N__37347));
    Span4Mux_v I__7922 (
            .O(N__37350),
            .I(N__37344));
    Span4Mux_v I__7921 (
            .O(N__37347),
            .I(N__37341));
    Span4Mux_h I__7920 (
            .O(N__37344),
            .I(N__37338));
    Sp12to4 I__7919 (
            .O(N__37341),
            .I(N__37335));
    Odrv4 I__7918 (
            .O(N__37338),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ));
    Odrv12 I__7917 (
            .O(N__37335),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ));
    InMux I__7916 (
            .O(N__37330),
            .I(N__37323));
    InMux I__7915 (
            .O(N__37329),
            .I(N__37323));
    InMux I__7914 (
            .O(N__37328),
            .I(N__37318));
    LocalMux I__7913 (
            .O(N__37323),
            .I(N__37314));
    InMux I__7912 (
            .O(N__37322),
            .I(N__37309));
    InMux I__7911 (
            .O(N__37321),
            .I(N__37309));
    LocalMux I__7910 (
            .O(N__37318),
            .I(N__37306));
    InMux I__7909 (
            .O(N__37317),
            .I(N__37303));
    Odrv12 I__7908 (
            .O(N__37314),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    LocalMux I__7907 (
            .O(N__37309),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    Odrv4 I__7906 (
            .O(N__37306),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    LocalMux I__7905 (
            .O(N__37303),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    InMux I__7904 (
            .O(N__37294),
            .I(N__37290));
    CascadeMux I__7903 (
            .O(N__37293),
            .I(N__37287));
    LocalMux I__7902 (
            .O(N__37290),
            .I(N__37282));
    InMux I__7901 (
            .O(N__37287),
            .I(N__37277));
    InMux I__7900 (
            .O(N__37286),
            .I(N__37277));
    InMux I__7899 (
            .O(N__37285),
            .I(N__37274));
    Odrv12 I__7898 (
            .O(N__37282),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    LocalMux I__7897 (
            .O(N__37277),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    LocalMux I__7896 (
            .O(N__37274),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    InMux I__7895 (
            .O(N__37267),
            .I(N__37264));
    LocalMux I__7894 (
            .O(N__37264),
            .I(N__37261));
    Odrv4 I__7893 (
            .O(N__37261),
            .I(\current_shift_inst.z_5_2 ));
    InMux I__7892 (
            .O(N__37258),
            .I(\current_shift_inst.z_5_cry_1 ));
    InMux I__7891 (
            .O(N__37255),
            .I(N__37252));
    LocalMux I__7890 (
            .O(N__37252),
            .I(N__37249));
    Odrv4 I__7889 (
            .O(N__37249),
            .I(\current_shift_inst.z_5_3 ));
    InMux I__7888 (
            .O(N__37246),
            .I(\current_shift_inst.z_5_cry_2 ));
    CascadeMux I__7887 (
            .O(N__37243),
            .I(N__37240));
    InMux I__7886 (
            .O(N__37240),
            .I(N__37237));
    LocalMux I__7885 (
            .O(N__37237),
            .I(N__37234));
    Odrv4 I__7884 (
            .O(N__37234),
            .I(\current_shift_inst.z_5_4 ));
    InMux I__7883 (
            .O(N__37231),
            .I(\current_shift_inst.z_5_cry_3 ));
    InMux I__7882 (
            .O(N__37228),
            .I(N__37225));
    LocalMux I__7881 (
            .O(N__37225),
            .I(N__37222));
    Odrv4 I__7880 (
            .O(N__37222),
            .I(\current_shift_inst.z_5_5 ));
    InMux I__7879 (
            .O(N__37219),
            .I(\current_shift_inst.z_5_cry_4 ));
    CascadeMux I__7878 (
            .O(N__37216),
            .I(N__37213));
    InMux I__7877 (
            .O(N__37213),
            .I(N__37210));
    LocalMux I__7876 (
            .O(N__37210),
            .I(N__37207));
    Odrv4 I__7875 (
            .O(N__37207),
            .I(\current_shift_inst.z_5_6 ));
    InMux I__7874 (
            .O(N__37204),
            .I(\current_shift_inst.z_5_cry_5 ));
    InMux I__7873 (
            .O(N__37201),
            .I(N__37198));
    LocalMux I__7872 (
            .O(N__37198),
            .I(N__37195));
    Odrv4 I__7871 (
            .O(N__37195),
            .I(\current_shift_inst.un4_control_input_axb_21 ));
    InMux I__7870 (
            .O(N__37192),
            .I(N__37189));
    LocalMux I__7869 (
            .O(N__37189),
            .I(N__37186));
    Span4Mux_h I__7868 (
            .O(N__37186),
            .I(N__37183));
    Odrv4 I__7867 (
            .O(N__37183),
            .I(\current_shift_inst.un4_control_input_axb_13 ));
    InMux I__7866 (
            .O(N__37180),
            .I(N__37176));
    InMux I__7865 (
            .O(N__37179),
            .I(N__37173));
    LocalMux I__7864 (
            .O(N__37176),
            .I(N__37169));
    LocalMux I__7863 (
            .O(N__37173),
            .I(N__37166));
    InMux I__7862 (
            .O(N__37172),
            .I(N__37163));
    Span4Mux_v I__7861 (
            .O(N__37169),
            .I(N__37158));
    Span4Mux_h I__7860 (
            .O(N__37166),
            .I(N__37158));
    LocalMux I__7859 (
            .O(N__37163),
            .I(measured_delay_tr_12));
    Odrv4 I__7858 (
            .O(N__37158),
            .I(measured_delay_tr_12));
    CascadeMux I__7857 (
            .O(N__37153),
            .I(N__37149));
    InMux I__7856 (
            .O(N__37152),
            .I(N__37145));
    InMux I__7855 (
            .O(N__37149),
            .I(N__37142));
    InMux I__7854 (
            .O(N__37148),
            .I(N__37139));
    LocalMux I__7853 (
            .O(N__37145),
            .I(N__37134));
    LocalMux I__7852 (
            .O(N__37142),
            .I(N__37134));
    LocalMux I__7851 (
            .O(N__37139),
            .I(measured_delay_tr_13));
    Odrv12 I__7850 (
            .O(N__37134),
            .I(measured_delay_tr_13));
    InMux I__7849 (
            .O(N__37129),
            .I(N__37124));
    InMux I__7848 (
            .O(N__37128),
            .I(N__37121));
    InMux I__7847 (
            .O(N__37127),
            .I(N__37118));
    LocalMux I__7846 (
            .O(N__37124),
            .I(N__37113));
    LocalMux I__7845 (
            .O(N__37121),
            .I(N__37113));
    LocalMux I__7844 (
            .O(N__37118),
            .I(measured_delay_tr_11));
    Odrv12 I__7843 (
            .O(N__37113),
            .I(measured_delay_tr_11));
    InMux I__7842 (
            .O(N__37108),
            .I(N__37103));
    InMux I__7841 (
            .O(N__37107),
            .I(N__37100));
    InMux I__7840 (
            .O(N__37106),
            .I(N__37097));
    LocalMux I__7839 (
            .O(N__37103),
            .I(N__37092));
    LocalMux I__7838 (
            .O(N__37100),
            .I(N__37092));
    LocalMux I__7837 (
            .O(N__37097),
            .I(measured_delay_tr_10));
    Odrv12 I__7836 (
            .O(N__37092),
            .I(measured_delay_tr_10));
    InMux I__7835 (
            .O(N__37087),
            .I(N__37084));
    LocalMux I__7834 (
            .O(N__37084),
            .I(\current_shift_inst.un4_control_input_axb_30 ));
    InMux I__7833 (
            .O(N__37081),
            .I(N__37078));
    LocalMux I__7832 (
            .O(N__37078),
            .I(\current_shift_inst.un4_control_input_axb_26 ));
    InMux I__7831 (
            .O(N__37075),
            .I(N__37072));
    LocalMux I__7830 (
            .O(N__37072),
            .I(\current_shift_inst.un4_control_input_axb_29 ));
    InMux I__7829 (
            .O(N__37069),
            .I(N__37066));
    LocalMux I__7828 (
            .O(N__37066),
            .I(\current_shift_inst.un4_control_input_axb_28 ));
    InMux I__7827 (
            .O(N__37063),
            .I(N__37060));
    LocalMux I__7826 (
            .O(N__37060),
            .I(\current_shift_inst.un4_control_input_axb_25 ));
    CascadeMux I__7825 (
            .O(N__37057),
            .I(N__37054));
    InMux I__7824 (
            .O(N__37054),
            .I(N__37051));
    LocalMux I__7823 (
            .O(N__37051),
            .I(N__37048));
    Span4Mux_v I__7822 (
            .O(N__37048),
            .I(N__37045));
    Odrv4 I__7821 (
            .O(N__37045),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__7820 (
            .O(N__37042),
            .I(N__37039));
    InMux I__7819 (
            .O(N__37039),
            .I(N__37036));
    LocalMux I__7818 (
            .O(N__37036),
            .I(N__37033));
    Span4Mux_v I__7817 (
            .O(N__37033),
            .I(N__37030));
    Odrv4 I__7816 (
            .O(N__37030),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__7815 (
            .O(N__37027),
            .I(N__37024));
    InMux I__7814 (
            .O(N__37024),
            .I(N__37021));
    LocalMux I__7813 (
            .O(N__37021),
            .I(N__37018));
    Span4Mux_v I__7812 (
            .O(N__37018),
            .I(N__37015));
    Odrv4 I__7811 (
            .O(N__37015),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__7810 (
            .O(N__37012),
            .I(N__37006));
    InMux I__7809 (
            .O(N__37011),
            .I(N__37002));
    InMux I__7808 (
            .O(N__37010),
            .I(N__36993));
    InMux I__7807 (
            .O(N__37009),
            .I(N__36993));
    InMux I__7806 (
            .O(N__37006),
            .I(N__36993));
    InMux I__7805 (
            .O(N__37005),
            .I(N__36993));
    LocalMux I__7804 (
            .O(N__37002),
            .I(N__36986));
    LocalMux I__7803 (
            .O(N__36993),
            .I(N__36983));
    InMux I__7802 (
            .O(N__36992),
            .I(N__36974));
    InMux I__7801 (
            .O(N__36991),
            .I(N__36974));
    InMux I__7800 (
            .O(N__36990),
            .I(N__36974));
    InMux I__7799 (
            .O(N__36989),
            .I(N__36974));
    Span4Mux_v I__7798 (
            .O(N__36986),
            .I(N__36966));
    Span4Mux_v I__7797 (
            .O(N__36983),
            .I(N__36966));
    LocalMux I__7796 (
            .O(N__36974),
            .I(N__36966));
    InMux I__7795 (
            .O(N__36973),
            .I(N__36963));
    Span4Mux_v I__7794 (
            .O(N__36966),
            .I(N__36958));
    LocalMux I__7793 (
            .O(N__36963),
            .I(N__36958));
    Span4Mux_h I__7792 (
            .O(N__36958),
            .I(N__36955));
    Odrv4 I__7791 (
            .O(N__36955),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ));
    CascadeMux I__7790 (
            .O(N__36952),
            .I(N__36949));
    InMux I__7789 (
            .O(N__36949),
            .I(N__36946));
    LocalMux I__7788 (
            .O(N__36946),
            .I(N__36943));
    Span4Mux_h I__7787 (
            .O(N__36943),
            .I(N__36940));
    Span4Mux_v I__7786 (
            .O(N__36940),
            .I(N__36937));
    Odrv4 I__7785 (
            .O(N__36937),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__7784 (
            .O(N__36934),
            .I(N__36931));
    LocalMux I__7783 (
            .O(N__36931),
            .I(\current_shift_inst.un4_control_input_axb_12 ));
    InMux I__7782 (
            .O(N__36928),
            .I(N__36925));
    LocalMux I__7781 (
            .O(N__36925),
            .I(\current_shift_inst.un4_control_input_axb_19 ));
    InMux I__7780 (
            .O(N__36922),
            .I(N__36919));
    LocalMux I__7779 (
            .O(N__36919),
            .I(\current_shift_inst.un4_control_input_axb_17 ));
    CascadeMux I__7778 (
            .O(N__36916),
            .I(N__36913));
    InMux I__7777 (
            .O(N__36913),
            .I(N__36910));
    LocalMux I__7776 (
            .O(N__36910),
            .I(\current_shift_inst.un4_control_input_axb_15 ));
    CascadeMux I__7775 (
            .O(N__36907),
            .I(N__36904));
    InMux I__7774 (
            .O(N__36904),
            .I(N__36901));
    LocalMux I__7773 (
            .O(N__36901),
            .I(\current_shift_inst.un4_control_input_axb_16 ));
    InMux I__7772 (
            .O(N__36898),
            .I(N__36895));
    LocalMux I__7771 (
            .O(N__36895),
            .I(\current_shift_inst.un4_control_input_axb_18 ));
    InMux I__7770 (
            .O(N__36892),
            .I(N__36889));
    LocalMux I__7769 (
            .O(N__36889),
            .I(\current_shift_inst.un4_control_input_axb_23 ));
    InMux I__7768 (
            .O(N__36886),
            .I(N__36883));
    LocalMux I__7767 (
            .O(N__36883),
            .I(\current_shift_inst.un4_control_input_axb_27 ));
    InMux I__7766 (
            .O(N__36880),
            .I(N__36877));
    LocalMux I__7765 (
            .O(N__36877),
            .I(\current_shift_inst.un4_control_input_axb_20 ));
    InMux I__7764 (
            .O(N__36874),
            .I(N__36871));
    LocalMux I__7763 (
            .O(N__36871),
            .I(\current_shift_inst.un4_control_input_axb_6 ));
    InMux I__7762 (
            .O(N__36868),
            .I(N__36865));
    LocalMux I__7761 (
            .O(N__36865),
            .I(\current_shift_inst.un4_control_input_axb_7 ));
    InMux I__7760 (
            .O(N__36862),
            .I(N__36859));
    LocalMux I__7759 (
            .O(N__36859),
            .I(\current_shift_inst.un4_control_input_axb_8 ));
    InMux I__7758 (
            .O(N__36856),
            .I(N__36853));
    LocalMux I__7757 (
            .O(N__36853),
            .I(\current_shift_inst.un4_control_input_axb_9 ));
    InMux I__7756 (
            .O(N__36850),
            .I(N__36847));
    LocalMux I__7755 (
            .O(N__36847),
            .I(\current_shift_inst.un4_control_input_axb_10 ));
    InMux I__7754 (
            .O(N__36844),
            .I(N__36841));
    LocalMux I__7753 (
            .O(N__36841),
            .I(\current_shift_inst.un4_control_input_axb_11 ));
    InMux I__7752 (
            .O(N__36838),
            .I(N__36835));
    LocalMux I__7751 (
            .O(N__36835),
            .I(\current_shift_inst.un4_control_input_axb_22 ));
    CascadeMux I__7750 (
            .O(N__36832),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_ ));
    InMux I__7749 (
            .O(N__36829),
            .I(N__36823));
    InMux I__7748 (
            .O(N__36828),
            .I(N__36823));
    LocalMux I__7747 (
            .O(N__36823),
            .I(N__36818));
    InMux I__7746 (
            .O(N__36822),
            .I(N__36815));
    CascadeMux I__7745 (
            .O(N__36821),
            .I(N__36812));
    Span4Mux_h I__7744 (
            .O(N__36818),
            .I(N__36808));
    LocalMux I__7743 (
            .O(N__36815),
            .I(N__36805));
    InMux I__7742 (
            .O(N__36812),
            .I(N__36802));
    InMux I__7741 (
            .O(N__36811),
            .I(N__36799));
    Span4Mux_v I__7740 (
            .O(N__36808),
            .I(N__36796));
    Span4Mux_h I__7739 (
            .O(N__36805),
            .I(N__36793));
    LocalMux I__7738 (
            .O(N__36802),
            .I(measured_delay_tr_14));
    LocalMux I__7737 (
            .O(N__36799),
            .I(measured_delay_tr_14));
    Odrv4 I__7736 (
            .O(N__36796),
            .I(measured_delay_tr_14));
    Odrv4 I__7735 (
            .O(N__36793),
            .I(measured_delay_tr_14));
    InMux I__7734 (
            .O(N__36784),
            .I(N__36781));
    LocalMux I__7733 (
            .O(N__36781),
            .I(\current_shift_inst.un4_control_input_axb_4 ));
    InMux I__7732 (
            .O(N__36778),
            .I(N__36775));
    LocalMux I__7731 (
            .O(N__36775),
            .I(\current_shift_inst.un4_control_input_axb_5 ));
    InMux I__7730 (
            .O(N__36772),
            .I(N__36769));
    LocalMux I__7729 (
            .O(N__36769),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ));
    CascadeMux I__7728 (
            .O(N__36766),
            .I(N__36763));
    InMux I__7727 (
            .O(N__36763),
            .I(N__36760));
    LocalMux I__7726 (
            .O(N__36760),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ));
    InMux I__7725 (
            .O(N__36757),
            .I(N__36754));
    LocalMux I__7724 (
            .O(N__36754),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ));
    CascadeMux I__7723 (
            .O(N__36751),
            .I(N__36748));
    InMux I__7722 (
            .O(N__36748),
            .I(N__36745));
    LocalMux I__7721 (
            .O(N__36745),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ));
    InMux I__7720 (
            .O(N__36742),
            .I(N__36739));
    LocalMux I__7719 (
            .O(N__36739),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ));
    InMux I__7718 (
            .O(N__36736),
            .I(N__36733));
    LocalMux I__7717 (
            .O(N__36733),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ));
    CascadeMux I__7716 (
            .O(N__36730),
            .I(N__36727));
    InMux I__7715 (
            .O(N__36727),
            .I(N__36724));
    LocalMux I__7714 (
            .O(N__36724),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ));
    InMux I__7713 (
            .O(N__36721),
            .I(N__36718));
    LocalMux I__7712 (
            .O(N__36718),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ));
    CascadeMux I__7711 (
            .O(N__36715),
            .I(N__36712));
    InMux I__7710 (
            .O(N__36712),
            .I(N__36709));
    LocalMux I__7709 (
            .O(N__36709),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ));
    InMux I__7708 (
            .O(N__36706),
            .I(N__36703));
    LocalMux I__7707 (
            .O(N__36703),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ));
    CascadeMux I__7706 (
            .O(N__36700),
            .I(N__36697));
    InMux I__7705 (
            .O(N__36697),
            .I(N__36694));
    LocalMux I__7704 (
            .O(N__36694),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ));
    CascadeMux I__7703 (
            .O(N__36691),
            .I(N__36688));
    InMux I__7702 (
            .O(N__36688),
            .I(N__36685));
    LocalMux I__7701 (
            .O(N__36685),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ));
    InMux I__7700 (
            .O(N__36682),
            .I(N__36679));
    LocalMux I__7699 (
            .O(N__36679),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ));
    CascadeMux I__7698 (
            .O(N__36676),
            .I(N__36673));
    InMux I__7697 (
            .O(N__36673),
            .I(N__36670));
    LocalMux I__7696 (
            .O(N__36670),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ));
    InMux I__7695 (
            .O(N__36667),
            .I(N__36643));
    InMux I__7694 (
            .O(N__36666),
            .I(N__36630));
    InMux I__7693 (
            .O(N__36665),
            .I(N__36630));
    InMux I__7692 (
            .O(N__36664),
            .I(N__36630));
    InMux I__7691 (
            .O(N__36663),
            .I(N__36630));
    InMux I__7690 (
            .O(N__36662),
            .I(N__36630));
    InMux I__7689 (
            .O(N__36661),
            .I(N__36630));
    InMux I__7688 (
            .O(N__36660),
            .I(N__36615));
    InMux I__7687 (
            .O(N__36659),
            .I(N__36615));
    InMux I__7686 (
            .O(N__36658),
            .I(N__36615));
    InMux I__7685 (
            .O(N__36657),
            .I(N__36615));
    InMux I__7684 (
            .O(N__36656),
            .I(N__36615));
    InMux I__7683 (
            .O(N__36655),
            .I(N__36615));
    InMux I__7682 (
            .O(N__36654),
            .I(N__36615));
    InMux I__7681 (
            .O(N__36653),
            .I(N__36596));
    InMux I__7680 (
            .O(N__36652),
            .I(N__36596));
    InMux I__7679 (
            .O(N__36651),
            .I(N__36596));
    InMux I__7678 (
            .O(N__36650),
            .I(N__36596));
    InMux I__7677 (
            .O(N__36649),
            .I(N__36596));
    InMux I__7676 (
            .O(N__36648),
            .I(N__36596));
    InMux I__7675 (
            .O(N__36647),
            .I(N__36596));
    InMux I__7674 (
            .O(N__36646),
            .I(N__36593));
    LocalMux I__7673 (
            .O(N__36643),
            .I(N__36588));
    LocalMux I__7672 (
            .O(N__36630),
            .I(N__36588));
    LocalMux I__7671 (
            .O(N__36615),
            .I(N__36581));
    InMux I__7670 (
            .O(N__36614),
            .I(N__36572));
    InMux I__7669 (
            .O(N__36613),
            .I(N__36572));
    InMux I__7668 (
            .O(N__36612),
            .I(N__36572));
    InMux I__7667 (
            .O(N__36611),
            .I(N__36572));
    LocalMux I__7666 (
            .O(N__36596),
            .I(N__36567));
    LocalMux I__7665 (
            .O(N__36593),
            .I(N__36567));
    Span4Mux_v I__7664 (
            .O(N__36588),
            .I(N__36558));
    InMux I__7663 (
            .O(N__36587),
            .I(N__36549));
    InMux I__7662 (
            .O(N__36586),
            .I(N__36549));
    InMux I__7661 (
            .O(N__36585),
            .I(N__36549));
    InMux I__7660 (
            .O(N__36584),
            .I(N__36549));
    Span4Mux_v I__7659 (
            .O(N__36581),
            .I(N__36544));
    LocalMux I__7658 (
            .O(N__36572),
            .I(N__36544));
    Span4Mux_h I__7657 (
            .O(N__36567),
            .I(N__36541));
    InMux I__7656 (
            .O(N__36566),
            .I(N__36534));
    InMux I__7655 (
            .O(N__36565),
            .I(N__36534));
    InMux I__7654 (
            .O(N__36564),
            .I(N__36534));
    InMux I__7653 (
            .O(N__36563),
            .I(N__36527));
    InMux I__7652 (
            .O(N__36562),
            .I(N__36527));
    InMux I__7651 (
            .O(N__36561),
            .I(N__36527));
    Sp12to4 I__7650 (
            .O(N__36558),
            .I(N__36520));
    LocalMux I__7649 (
            .O(N__36549),
            .I(N__36520));
    Span4Mux_h I__7648 (
            .O(N__36544),
            .I(N__36517));
    Span4Mux_h I__7647 (
            .O(N__36541),
            .I(N__36510));
    LocalMux I__7646 (
            .O(N__36534),
            .I(N__36510));
    LocalMux I__7645 (
            .O(N__36527),
            .I(N__36510));
    InMux I__7644 (
            .O(N__36526),
            .I(N__36505));
    InMux I__7643 (
            .O(N__36525),
            .I(N__36505));
    Odrv12 I__7642 (
            .O(N__36520),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv4 I__7641 (
            .O(N__36517),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv4 I__7640 (
            .O(N__36510),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    LocalMux I__7639 (
            .O(N__36505),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    InMux I__7638 (
            .O(N__36496),
            .I(N__36492));
    CascadeMux I__7637 (
            .O(N__36495),
            .I(N__36487));
    LocalMux I__7636 (
            .O(N__36492),
            .I(N__36484));
    InMux I__7635 (
            .O(N__36491),
            .I(N__36481));
    InMux I__7634 (
            .O(N__36490),
            .I(N__36478));
    InMux I__7633 (
            .O(N__36487),
            .I(N__36474));
    Span4Mux_h I__7632 (
            .O(N__36484),
            .I(N__36471));
    LocalMux I__7631 (
            .O(N__36481),
            .I(N__36468));
    LocalMux I__7630 (
            .O(N__36478),
            .I(N__36465));
    InMux I__7629 (
            .O(N__36477),
            .I(N__36462));
    LocalMux I__7628 (
            .O(N__36474),
            .I(measured_delay_hc_8));
    Odrv4 I__7627 (
            .O(N__36471),
            .I(measured_delay_hc_8));
    Odrv12 I__7626 (
            .O(N__36468),
            .I(measured_delay_hc_8));
    Odrv4 I__7625 (
            .O(N__36465),
            .I(measured_delay_hc_8));
    LocalMux I__7624 (
            .O(N__36462),
            .I(measured_delay_hc_8));
    CascadeMux I__7623 (
            .O(N__36451),
            .I(N__36446));
    CascadeMux I__7622 (
            .O(N__36450),
            .I(N__36434));
    CascadeMux I__7621 (
            .O(N__36449),
            .I(N__36431));
    InMux I__7620 (
            .O(N__36446),
            .I(N__36422));
    InMux I__7619 (
            .O(N__36445),
            .I(N__36422));
    InMux I__7618 (
            .O(N__36444),
            .I(N__36422));
    InMux I__7617 (
            .O(N__36443),
            .I(N__36422));
    CascadeMux I__7616 (
            .O(N__36442),
            .I(N__36414));
    InMux I__7615 (
            .O(N__36441),
            .I(N__36399));
    InMux I__7614 (
            .O(N__36440),
            .I(N__36399));
    InMux I__7613 (
            .O(N__36439),
            .I(N__36399));
    InMux I__7612 (
            .O(N__36438),
            .I(N__36399));
    InMux I__7611 (
            .O(N__36437),
            .I(N__36399));
    InMux I__7610 (
            .O(N__36434),
            .I(N__36399));
    InMux I__7609 (
            .O(N__36431),
            .I(N__36399));
    LocalMux I__7608 (
            .O(N__36422),
            .I(N__36393));
    InMux I__7607 (
            .O(N__36421),
            .I(N__36386));
    InMux I__7606 (
            .O(N__36420),
            .I(N__36386));
    InMux I__7605 (
            .O(N__36419),
            .I(N__36386));
    InMux I__7604 (
            .O(N__36418),
            .I(N__36379));
    InMux I__7603 (
            .O(N__36417),
            .I(N__36379));
    InMux I__7602 (
            .O(N__36414),
            .I(N__36379));
    LocalMux I__7601 (
            .O(N__36399),
            .I(N__36376));
    InMux I__7600 (
            .O(N__36398),
            .I(N__36369));
    InMux I__7599 (
            .O(N__36397),
            .I(N__36369));
    InMux I__7598 (
            .O(N__36396),
            .I(N__36369));
    Span4Mux_h I__7597 (
            .O(N__36393),
            .I(N__36362));
    LocalMux I__7596 (
            .O(N__36386),
            .I(N__36362));
    LocalMux I__7595 (
            .O(N__36379),
            .I(N__36354));
    Span4Mux_h I__7594 (
            .O(N__36376),
            .I(N__36349));
    LocalMux I__7593 (
            .O(N__36369),
            .I(N__36349));
    CascadeMux I__7592 (
            .O(N__36368),
            .I(N__36345));
    CascadeMux I__7591 (
            .O(N__36367),
            .I(N__36341));
    Span4Mux_v I__7590 (
            .O(N__36362),
            .I(N__36336));
    CascadeMux I__7589 (
            .O(N__36361),
            .I(N__36332));
    CascadeMux I__7588 (
            .O(N__36360),
            .I(N__36329));
    CascadeMux I__7587 (
            .O(N__36359),
            .I(N__36326));
    CascadeMux I__7586 (
            .O(N__36358),
            .I(N__36322));
    CascadeMux I__7585 (
            .O(N__36357),
            .I(N__36311));
    Span4Mux_v I__7584 (
            .O(N__36354),
            .I(N__36306));
    Span4Mux_h I__7583 (
            .O(N__36349),
            .I(N__36306));
    InMux I__7582 (
            .O(N__36348),
            .I(N__36295));
    InMux I__7581 (
            .O(N__36345),
            .I(N__36295));
    InMux I__7580 (
            .O(N__36344),
            .I(N__36295));
    InMux I__7579 (
            .O(N__36341),
            .I(N__36295));
    InMux I__7578 (
            .O(N__36340),
            .I(N__36295));
    InMux I__7577 (
            .O(N__36339),
            .I(N__36292));
    Span4Mux_h I__7576 (
            .O(N__36336),
            .I(N__36289));
    InMux I__7575 (
            .O(N__36335),
            .I(N__36286));
    InMux I__7574 (
            .O(N__36332),
            .I(N__36271));
    InMux I__7573 (
            .O(N__36329),
            .I(N__36271));
    InMux I__7572 (
            .O(N__36326),
            .I(N__36271));
    InMux I__7571 (
            .O(N__36325),
            .I(N__36271));
    InMux I__7570 (
            .O(N__36322),
            .I(N__36271));
    InMux I__7569 (
            .O(N__36321),
            .I(N__36271));
    InMux I__7568 (
            .O(N__36320),
            .I(N__36271));
    InMux I__7567 (
            .O(N__36319),
            .I(N__36268));
    InMux I__7566 (
            .O(N__36318),
            .I(N__36255));
    InMux I__7565 (
            .O(N__36317),
            .I(N__36255));
    InMux I__7564 (
            .O(N__36316),
            .I(N__36255));
    InMux I__7563 (
            .O(N__36315),
            .I(N__36255));
    InMux I__7562 (
            .O(N__36314),
            .I(N__36255));
    InMux I__7561 (
            .O(N__36311),
            .I(N__36255));
    Span4Mux_h I__7560 (
            .O(N__36306),
            .I(N__36250));
    LocalMux I__7559 (
            .O(N__36295),
            .I(N__36250));
    LocalMux I__7558 (
            .O(N__36292),
            .I(measured_delay_hc_31));
    Odrv4 I__7557 (
            .O(N__36289),
            .I(measured_delay_hc_31));
    LocalMux I__7556 (
            .O(N__36286),
            .I(measured_delay_hc_31));
    LocalMux I__7555 (
            .O(N__36271),
            .I(measured_delay_hc_31));
    LocalMux I__7554 (
            .O(N__36268),
            .I(measured_delay_hc_31));
    LocalMux I__7553 (
            .O(N__36255),
            .I(measured_delay_hc_31));
    Odrv4 I__7552 (
            .O(N__36250),
            .I(measured_delay_hc_31));
    CascadeMux I__7551 (
            .O(N__36235),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    CEMux I__7550 (
            .O(N__36232),
            .I(N__36228));
    CEMux I__7549 (
            .O(N__36231),
            .I(N__36223));
    LocalMux I__7548 (
            .O(N__36228),
            .I(N__36219));
    CEMux I__7547 (
            .O(N__36227),
            .I(N__36216));
    CEMux I__7546 (
            .O(N__36226),
            .I(N__36213));
    LocalMux I__7545 (
            .O(N__36223),
            .I(N__36210));
    CEMux I__7544 (
            .O(N__36222),
            .I(N__36207));
    Span4Mux_v I__7543 (
            .O(N__36219),
            .I(N__36202));
    LocalMux I__7542 (
            .O(N__36216),
            .I(N__36202));
    LocalMux I__7541 (
            .O(N__36213),
            .I(N__36199));
    Span4Mux_v I__7540 (
            .O(N__36210),
            .I(N__36196));
    LocalMux I__7539 (
            .O(N__36207),
            .I(N__36193));
    Span4Mux_h I__7538 (
            .O(N__36202),
            .I(N__36190));
    Span4Mux_v I__7537 (
            .O(N__36199),
            .I(N__36185));
    Span4Mux_h I__7536 (
            .O(N__36196),
            .I(N__36185));
    Odrv12 I__7535 (
            .O(N__36193),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__7534 (
            .O(N__36190),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__7533 (
            .O(N__36185),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__7532 (
            .O(N__36178),
            .I(N__36175));
    LocalMux I__7531 (
            .O(N__36175),
            .I(N__36172));
    Odrv4 I__7530 (
            .O(N__36172),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ));
    InMux I__7529 (
            .O(N__36169),
            .I(N__36166));
    LocalMux I__7528 (
            .O(N__36166),
            .I(N__36163));
    Odrv4 I__7527 (
            .O(N__36163),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ));
    CascadeMux I__7526 (
            .O(N__36160),
            .I(N__36157));
    InMux I__7525 (
            .O(N__36157),
            .I(N__36154));
    LocalMux I__7524 (
            .O(N__36154),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ));
    InMux I__7523 (
            .O(N__36151),
            .I(N__36146));
    InMux I__7522 (
            .O(N__36150),
            .I(N__36143));
    CascadeMux I__7521 (
            .O(N__36149),
            .I(N__36140));
    LocalMux I__7520 (
            .O(N__36146),
            .I(N__36136));
    LocalMux I__7519 (
            .O(N__36143),
            .I(N__36133));
    InMux I__7518 (
            .O(N__36140),
            .I(N__36130));
    CascadeMux I__7517 (
            .O(N__36139),
            .I(N__36126));
    Span4Mux_h I__7516 (
            .O(N__36136),
            .I(N__36123));
    Span4Mux_v I__7515 (
            .O(N__36133),
            .I(N__36120));
    LocalMux I__7514 (
            .O(N__36130),
            .I(N__36117));
    InMux I__7513 (
            .O(N__36129),
            .I(N__36114));
    InMux I__7512 (
            .O(N__36126),
            .I(N__36111));
    Span4Mux_h I__7511 (
            .O(N__36123),
            .I(N__36108));
    Span4Mux_h I__7510 (
            .O(N__36120),
            .I(N__36101));
    Span4Mux_v I__7509 (
            .O(N__36117),
            .I(N__36101));
    LocalMux I__7508 (
            .O(N__36114),
            .I(N__36101));
    LocalMux I__7507 (
            .O(N__36111),
            .I(measured_delay_hc_5));
    Odrv4 I__7506 (
            .O(N__36108),
            .I(measured_delay_hc_5));
    Odrv4 I__7505 (
            .O(N__36101),
            .I(measured_delay_hc_5));
    CascadeMux I__7504 (
            .O(N__36094),
            .I(N__36091));
    InMux I__7503 (
            .O(N__36091),
            .I(N__36088));
    LocalMux I__7502 (
            .O(N__36088),
            .I(N__36082));
    InMux I__7501 (
            .O(N__36087),
            .I(N__36079));
    CascadeMux I__7500 (
            .O(N__36086),
            .I(N__36076));
    InMux I__7499 (
            .O(N__36085),
            .I(N__36073));
    Span4Mux_h I__7498 (
            .O(N__36082),
            .I(N__36070));
    LocalMux I__7497 (
            .O(N__36079),
            .I(N__36067));
    InMux I__7496 (
            .O(N__36076),
            .I(N__36064));
    LocalMux I__7495 (
            .O(N__36073),
            .I(N__36060));
    Span4Mux_h I__7494 (
            .O(N__36070),
            .I(N__36055));
    Span4Mux_h I__7493 (
            .O(N__36067),
            .I(N__36055));
    LocalMux I__7492 (
            .O(N__36064),
            .I(N__36052));
    InMux I__7491 (
            .O(N__36063),
            .I(N__36049));
    Span4Mux_h I__7490 (
            .O(N__36060),
            .I(N__36046));
    Span4Mux_v I__7489 (
            .O(N__36055),
            .I(N__36043));
    Span4Mux_v I__7488 (
            .O(N__36052),
            .I(N__36040));
    LocalMux I__7487 (
            .O(N__36049),
            .I(measured_delay_hc_3));
    Odrv4 I__7486 (
            .O(N__36046),
            .I(measured_delay_hc_3));
    Odrv4 I__7485 (
            .O(N__36043),
            .I(measured_delay_hc_3));
    Odrv4 I__7484 (
            .O(N__36040),
            .I(measured_delay_hc_3));
    InMux I__7483 (
            .O(N__36031),
            .I(N__36028));
    LocalMux I__7482 (
            .O(N__36028),
            .I(N__36024));
    InMux I__7481 (
            .O(N__36027),
            .I(N__36021));
    Span4Mux_h I__7480 (
            .O(N__36024),
            .I(N__36015));
    LocalMux I__7479 (
            .O(N__36021),
            .I(N__36012));
    InMux I__7478 (
            .O(N__36020),
            .I(N__36009));
    CascadeMux I__7477 (
            .O(N__36019),
            .I(N__36006));
    InMux I__7476 (
            .O(N__36018),
            .I(N__36003));
    Span4Mux_h I__7475 (
            .O(N__36015),
            .I(N__35996));
    Span4Mux_h I__7474 (
            .O(N__36012),
            .I(N__35996));
    LocalMux I__7473 (
            .O(N__36009),
            .I(N__35996));
    InMux I__7472 (
            .O(N__36006),
            .I(N__35993));
    LocalMux I__7471 (
            .O(N__36003),
            .I(measured_delay_hc_13));
    Odrv4 I__7470 (
            .O(N__35996),
            .I(measured_delay_hc_13));
    LocalMux I__7469 (
            .O(N__35993),
            .I(measured_delay_hc_13));
    InMux I__7468 (
            .O(N__35986),
            .I(N__35980));
    InMux I__7467 (
            .O(N__35985),
            .I(N__35977));
    CascadeMux I__7466 (
            .O(N__35984),
            .I(N__35974));
    InMux I__7465 (
            .O(N__35983),
            .I(N__35971));
    LocalMux I__7464 (
            .O(N__35980),
            .I(N__35968));
    LocalMux I__7463 (
            .O(N__35977),
            .I(N__35963));
    InMux I__7462 (
            .O(N__35974),
            .I(N__35960));
    LocalMux I__7461 (
            .O(N__35971),
            .I(N__35957));
    Span4Mux_v I__7460 (
            .O(N__35968),
            .I(N__35954));
    InMux I__7459 (
            .O(N__35967),
            .I(N__35951));
    InMux I__7458 (
            .O(N__35966),
            .I(N__35948));
    Span4Mux_h I__7457 (
            .O(N__35963),
            .I(N__35945));
    LocalMux I__7456 (
            .O(N__35960),
            .I(measured_delay_hc_9));
    Odrv12 I__7455 (
            .O(N__35957),
            .I(measured_delay_hc_9));
    Odrv4 I__7454 (
            .O(N__35954),
            .I(measured_delay_hc_9));
    LocalMux I__7453 (
            .O(N__35951),
            .I(measured_delay_hc_9));
    LocalMux I__7452 (
            .O(N__35948),
            .I(measured_delay_hc_9));
    Odrv4 I__7451 (
            .O(N__35945),
            .I(measured_delay_hc_9));
    InMux I__7450 (
            .O(N__35932),
            .I(N__35927));
    InMux I__7449 (
            .O(N__35931),
            .I(N__35924));
    InMux I__7448 (
            .O(N__35930),
            .I(N__35920));
    LocalMux I__7447 (
            .O(N__35927),
            .I(N__35917));
    LocalMux I__7446 (
            .O(N__35924),
            .I(N__35914));
    InMux I__7445 (
            .O(N__35923),
            .I(N__35911));
    LocalMux I__7444 (
            .O(N__35920),
            .I(N__35905));
    Span4Mux_h I__7443 (
            .O(N__35917),
            .I(N__35905));
    Span4Mux_h I__7442 (
            .O(N__35914),
            .I(N__35900));
    LocalMux I__7441 (
            .O(N__35911),
            .I(N__35900));
    InMux I__7440 (
            .O(N__35910),
            .I(N__35897));
    Odrv4 I__7439 (
            .O(N__35905),
            .I(measured_delay_hc_10));
    Odrv4 I__7438 (
            .O(N__35900),
            .I(measured_delay_hc_10));
    LocalMux I__7437 (
            .O(N__35897),
            .I(measured_delay_hc_10));
    InMux I__7436 (
            .O(N__35890),
            .I(N__35885));
    InMux I__7435 (
            .O(N__35889),
            .I(N__35882));
    InMux I__7434 (
            .O(N__35888),
            .I(N__35878));
    LocalMux I__7433 (
            .O(N__35885),
            .I(N__35875));
    LocalMux I__7432 (
            .O(N__35882),
            .I(N__35872));
    InMux I__7431 (
            .O(N__35881),
            .I(N__35869));
    LocalMux I__7430 (
            .O(N__35878),
            .I(N__35863));
    Span4Mux_h I__7429 (
            .O(N__35875),
            .I(N__35863));
    Span4Mux_h I__7428 (
            .O(N__35872),
            .I(N__35858));
    LocalMux I__7427 (
            .O(N__35869),
            .I(N__35858));
    InMux I__7426 (
            .O(N__35868),
            .I(N__35855));
    Odrv4 I__7425 (
            .O(N__35863),
            .I(measured_delay_hc_11));
    Odrv4 I__7424 (
            .O(N__35858),
            .I(measured_delay_hc_11));
    LocalMux I__7423 (
            .O(N__35855),
            .I(measured_delay_hc_11));
    CascadeMux I__7422 (
            .O(N__35848),
            .I(N__35845));
    InMux I__7421 (
            .O(N__35845),
            .I(N__35842));
    LocalMux I__7420 (
            .O(N__35842),
            .I(N__35838));
    InMux I__7419 (
            .O(N__35841),
            .I(N__35834));
    Span4Mux_v I__7418 (
            .O(N__35838),
            .I(N__35831));
    InMux I__7417 (
            .O(N__35837),
            .I(N__35828));
    LocalMux I__7416 (
            .O(N__35834),
            .I(N__35824));
    Span4Mux_h I__7415 (
            .O(N__35831),
            .I(N__35819));
    LocalMux I__7414 (
            .O(N__35828),
            .I(N__35819));
    InMux I__7413 (
            .O(N__35827),
            .I(N__35816));
    Span4Mux_h I__7412 (
            .O(N__35824),
            .I(N__35813));
    Span4Mux_h I__7411 (
            .O(N__35819),
            .I(N__35810));
    LocalMux I__7410 (
            .O(N__35816),
            .I(measured_delay_hc_0));
    Odrv4 I__7409 (
            .O(N__35813),
            .I(measured_delay_hc_0));
    Odrv4 I__7408 (
            .O(N__35810),
            .I(measured_delay_hc_0));
    CascadeMux I__7407 (
            .O(N__35803),
            .I(N__35798));
    CascadeMux I__7406 (
            .O(N__35802),
            .I(N__35795));
    CascadeMux I__7405 (
            .O(N__35801),
            .I(N__35792));
    InMux I__7404 (
            .O(N__35798),
            .I(N__35781));
    InMux I__7403 (
            .O(N__35795),
            .I(N__35781));
    InMux I__7402 (
            .O(N__35792),
            .I(N__35781));
    InMux I__7401 (
            .O(N__35791),
            .I(N__35781));
    InMux I__7400 (
            .O(N__35790),
            .I(N__35770));
    LocalMux I__7399 (
            .O(N__35781),
            .I(N__35766));
    InMux I__7398 (
            .O(N__35780),
            .I(N__35759));
    InMux I__7397 (
            .O(N__35779),
            .I(N__35759));
    InMux I__7396 (
            .O(N__35778),
            .I(N__35759));
    InMux I__7395 (
            .O(N__35777),
            .I(N__35748));
    InMux I__7394 (
            .O(N__35776),
            .I(N__35748));
    InMux I__7393 (
            .O(N__35775),
            .I(N__35748));
    InMux I__7392 (
            .O(N__35774),
            .I(N__35748));
    InMux I__7391 (
            .O(N__35773),
            .I(N__35748));
    LocalMux I__7390 (
            .O(N__35770),
            .I(N__35745));
    InMux I__7389 (
            .O(N__35769),
            .I(N__35742));
    Span4Mux_v I__7388 (
            .O(N__35766),
            .I(N__35737));
    LocalMux I__7387 (
            .O(N__35759),
            .I(N__35737));
    LocalMux I__7386 (
            .O(N__35748),
            .I(N__35734));
    Span4Mux_v I__7385 (
            .O(N__35745),
            .I(N__35729));
    LocalMux I__7384 (
            .O(N__35742),
            .I(N__35729));
    Span4Mux_h I__7383 (
            .O(N__35737),
            .I(N__35726));
    Span4Mux_h I__7382 (
            .O(N__35734),
            .I(N__35723));
    Span4Mux_h I__7381 (
            .O(N__35729),
            .I(N__35720));
    Odrv4 I__7380 (
            .O(N__35726),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    Odrv4 I__7379 (
            .O(N__35723),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    Odrv4 I__7378 (
            .O(N__35720),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    InMux I__7377 (
            .O(N__35713),
            .I(N__35710));
    LocalMux I__7376 (
            .O(N__35710),
            .I(N__35705));
    CascadeMux I__7375 (
            .O(N__35709),
            .I(N__35701));
    InMux I__7374 (
            .O(N__35708),
            .I(N__35698));
    Span4Mux_h I__7373 (
            .O(N__35705),
            .I(N__35695));
    InMux I__7372 (
            .O(N__35704),
            .I(N__35692));
    InMux I__7371 (
            .O(N__35701),
            .I(N__35688));
    LocalMux I__7370 (
            .O(N__35698),
            .I(N__35685));
    Span4Mux_h I__7369 (
            .O(N__35695),
            .I(N__35680));
    LocalMux I__7368 (
            .O(N__35692),
            .I(N__35680));
    InMux I__7367 (
            .O(N__35691),
            .I(N__35677));
    LocalMux I__7366 (
            .O(N__35688),
            .I(measured_delay_hc_1));
    Odrv12 I__7365 (
            .O(N__35685),
            .I(measured_delay_hc_1));
    Odrv4 I__7364 (
            .O(N__35680),
            .I(measured_delay_hc_1));
    LocalMux I__7363 (
            .O(N__35677),
            .I(measured_delay_hc_1));
    InMux I__7362 (
            .O(N__35668),
            .I(N__35665));
    LocalMux I__7361 (
            .O(N__35665),
            .I(N__35659));
    InMux I__7360 (
            .O(N__35664),
            .I(N__35655));
    CascadeMux I__7359 (
            .O(N__35663),
            .I(N__35652));
    InMux I__7358 (
            .O(N__35662),
            .I(N__35649));
    Span4Mux_h I__7357 (
            .O(N__35659),
            .I(N__35646));
    InMux I__7356 (
            .O(N__35658),
            .I(N__35643));
    LocalMux I__7355 (
            .O(N__35655),
            .I(N__35640));
    InMux I__7354 (
            .O(N__35652),
            .I(N__35637));
    LocalMux I__7353 (
            .O(N__35649),
            .I(N__35634));
    Span4Mux_h I__7352 (
            .O(N__35646),
            .I(N__35631));
    LocalMux I__7351 (
            .O(N__35643),
            .I(N__35628));
    Span4Mux_v I__7350 (
            .O(N__35640),
            .I(N__35625));
    LocalMux I__7349 (
            .O(N__35637),
            .I(measured_delay_hc_15));
    Odrv12 I__7348 (
            .O(N__35634),
            .I(measured_delay_hc_15));
    Odrv4 I__7347 (
            .O(N__35631),
            .I(measured_delay_hc_15));
    Odrv4 I__7346 (
            .O(N__35628),
            .I(measured_delay_hc_15));
    Odrv4 I__7345 (
            .O(N__35625),
            .I(measured_delay_hc_15));
    InMux I__7344 (
            .O(N__35614),
            .I(\current_shift_inst.timer_phase.counter_cry_26 ));
    InMux I__7343 (
            .O(N__35611),
            .I(\current_shift_inst.timer_phase.counter_cry_27 ));
    InMux I__7342 (
            .O(N__35608),
            .I(N__35570));
    InMux I__7341 (
            .O(N__35607),
            .I(N__35570));
    InMux I__7340 (
            .O(N__35606),
            .I(N__35570));
    InMux I__7339 (
            .O(N__35605),
            .I(N__35570));
    InMux I__7338 (
            .O(N__35604),
            .I(N__35561));
    InMux I__7337 (
            .O(N__35603),
            .I(N__35561));
    InMux I__7336 (
            .O(N__35602),
            .I(N__35561));
    InMux I__7335 (
            .O(N__35601),
            .I(N__35561));
    InMux I__7334 (
            .O(N__35600),
            .I(N__35556));
    InMux I__7333 (
            .O(N__35599),
            .I(N__35556));
    InMux I__7332 (
            .O(N__35598),
            .I(N__35547));
    InMux I__7331 (
            .O(N__35597),
            .I(N__35547));
    InMux I__7330 (
            .O(N__35596),
            .I(N__35547));
    InMux I__7329 (
            .O(N__35595),
            .I(N__35547));
    InMux I__7328 (
            .O(N__35594),
            .I(N__35538));
    InMux I__7327 (
            .O(N__35593),
            .I(N__35538));
    InMux I__7326 (
            .O(N__35592),
            .I(N__35538));
    InMux I__7325 (
            .O(N__35591),
            .I(N__35538));
    InMux I__7324 (
            .O(N__35590),
            .I(N__35529));
    InMux I__7323 (
            .O(N__35589),
            .I(N__35529));
    InMux I__7322 (
            .O(N__35588),
            .I(N__35529));
    InMux I__7321 (
            .O(N__35587),
            .I(N__35529));
    InMux I__7320 (
            .O(N__35586),
            .I(N__35520));
    InMux I__7319 (
            .O(N__35585),
            .I(N__35520));
    InMux I__7318 (
            .O(N__35584),
            .I(N__35520));
    InMux I__7317 (
            .O(N__35583),
            .I(N__35520));
    InMux I__7316 (
            .O(N__35582),
            .I(N__35511));
    InMux I__7315 (
            .O(N__35581),
            .I(N__35511));
    InMux I__7314 (
            .O(N__35580),
            .I(N__35511));
    InMux I__7313 (
            .O(N__35579),
            .I(N__35511));
    LocalMux I__7312 (
            .O(N__35570),
            .I(N__35506));
    LocalMux I__7311 (
            .O(N__35561),
            .I(N__35506));
    LocalMux I__7310 (
            .O(N__35556),
            .I(N__35497));
    LocalMux I__7309 (
            .O(N__35547),
            .I(N__35497));
    LocalMux I__7308 (
            .O(N__35538),
            .I(N__35497));
    LocalMux I__7307 (
            .O(N__35529),
            .I(N__35497));
    LocalMux I__7306 (
            .O(N__35520),
            .I(N__35488));
    LocalMux I__7305 (
            .O(N__35511),
            .I(N__35488));
    Span4Mux_v I__7304 (
            .O(N__35506),
            .I(N__35488));
    Span4Mux_v I__7303 (
            .O(N__35497),
            .I(N__35488));
    Odrv4 I__7302 (
            .O(N__35488),
            .I(\current_shift_inst.timer_phase.running_i ));
    InMux I__7301 (
            .O(N__35485),
            .I(\current_shift_inst.timer_phase.counter_cry_28 ));
    CEMux I__7300 (
            .O(N__35482),
            .I(N__35477));
    CEMux I__7299 (
            .O(N__35481),
            .I(N__35473));
    CEMux I__7298 (
            .O(N__35480),
            .I(N__35470));
    LocalMux I__7297 (
            .O(N__35477),
            .I(N__35467));
    CEMux I__7296 (
            .O(N__35476),
            .I(N__35464));
    LocalMux I__7295 (
            .O(N__35473),
            .I(N__35459));
    LocalMux I__7294 (
            .O(N__35470),
            .I(N__35459));
    Span4Mux_v I__7293 (
            .O(N__35467),
            .I(N__35454));
    LocalMux I__7292 (
            .O(N__35464),
            .I(N__35454));
    Span4Mux_v I__7291 (
            .O(N__35459),
            .I(N__35451));
    Span4Mux_v I__7290 (
            .O(N__35454),
            .I(N__35446));
    Span4Mux_h I__7289 (
            .O(N__35451),
            .I(N__35446));
    Odrv4 I__7288 (
            .O(N__35446),
            .I(\current_shift_inst.timer_phase.N_192_i ));
    InMux I__7287 (
            .O(N__35443),
            .I(N__35440));
    LocalMux I__7286 (
            .O(N__35440),
            .I(N__35437));
    Odrv12 I__7285 (
            .O(N__35437),
            .I(delay_tr_input_c));
    InMux I__7284 (
            .O(N__35434),
            .I(N__35431));
    LocalMux I__7283 (
            .O(N__35431),
            .I(delay_tr_d1));
    InMux I__7282 (
            .O(N__35428),
            .I(N__35425));
    LocalMux I__7281 (
            .O(N__35425),
            .I(N__35420));
    InMux I__7280 (
            .O(N__35424),
            .I(N__35417));
    CascadeMux I__7279 (
            .O(N__35423),
            .I(N__35413));
    Span4Mux_h I__7278 (
            .O(N__35420),
            .I(N__35410));
    LocalMux I__7277 (
            .O(N__35417),
            .I(N__35407));
    InMux I__7276 (
            .O(N__35416),
            .I(N__35404));
    InMux I__7275 (
            .O(N__35413),
            .I(N__35400));
    Span4Mux_h I__7274 (
            .O(N__35410),
            .I(N__35397));
    Span4Mux_v I__7273 (
            .O(N__35407),
            .I(N__35392));
    LocalMux I__7272 (
            .O(N__35404),
            .I(N__35392));
    InMux I__7271 (
            .O(N__35403),
            .I(N__35389));
    LocalMux I__7270 (
            .O(N__35400),
            .I(measured_delay_hc_7));
    Odrv4 I__7269 (
            .O(N__35397),
            .I(measured_delay_hc_7));
    Odrv4 I__7268 (
            .O(N__35392),
            .I(measured_delay_hc_7));
    LocalMux I__7267 (
            .O(N__35389),
            .I(measured_delay_hc_7));
    CascadeMux I__7266 (
            .O(N__35380),
            .I(N__35375));
    InMux I__7265 (
            .O(N__35379),
            .I(N__35371));
    CascadeMux I__7264 (
            .O(N__35378),
            .I(N__35367));
    InMux I__7263 (
            .O(N__35375),
            .I(N__35364));
    InMux I__7262 (
            .O(N__35374),
            .I(N__35361));
    LocalMux I__7261 (
            .O(N__35371),
            .I(N__35358));
    InMux I__7260 (
            .O(N__35370),
            .I(N__35355));
    InMux I__7259 (
            .O(N__35367),
            .I(N__35352));
    LocalMux I__7258 (
            .O(N__35364),
            .I(N__35349));
    LocalMux I__7257 (
            .O(N__35361),
            .I(N__35346));
    Span4Mux_v I__7256 (
            .O(N__35358),
            .I(N__35341));
    LocalMux I__7255 (
            .O(N__35355),
            .I(N__35341));
    LocalMux I__7254 (
            .O(N__35352),
            .I(N__35336));
    Span4Mux_v I__7253 (
            .O(N__35349),
            .I(N__35336));
    Span12Mux_h I__7252 (
            .O(N__35346),
            .I(N__35333));
    Span4Mux_h I__7251 (
            .O(N__35341),
            .I(N__35330));
    Odrv4 I__7250 (
            .O(N__35336),
            .I(measured_delay_hc_2));
    Odrv12 I__7249 (
            .O(N__35333),
            .I(measured_delay_hc_2));
    Odrv4 I__7248 (
            .O(N__35330),
            .I(measured_delay_hc_2));
    InMux I__7247 (
            .O(N__35323),
            .I(N__35320));
    LocalMux I__7246 (
            .O(N__35320),
            .I(N__35316));
    InMux I__7245 (
            .O(N__35319),
            .I(N__35310));
    Span4Mux_v I__7244 (
            .O(N__35316),
            .I(N__35307));
    InMux I__7243 (
            .O(N__35315),
            .I(N__35304));
    InMux I__7242 (
            .O(N__35314),
            .I(N__35301));
    CascadeMux I__7241 (
            .O(N__35313),
            .I(N__35298));
    LocalMux I__7240 (
            .O(N__35310),
            .I(N__35295));
    Sp12to4 I__7239 (
            .O(N__35307),
            .I(N__35290));
    LocalMux I__7238 (
            .O(N__35304),
            .I(N__35290));
    LocalMux I__7237 (
            .O(N__35301),
            .I(N__35287));
    InMux I__7236 (
            .O(N__35298),
            .I(N__35284));
    Span12Mux_h I__7235 (
            .O(N__35295),
            .I(N__35281));
    Span12Mux_h I__7234 (
            .O(N__35290),
            .I(N__35278));
    Span4Mux_h I__7233 (
            .O(N__35287),
            .I(N__35275));
    LocalMux I__7232 (
            .O(N__35284),
            .I(measured_delay_hc_6));
    Odrv12 I__7231 (
            .O(N__35281),
            .I(measured_delay_hc_6));
    Odrv12 I__7230 (
            .O(N__35278),
            .I(measured_delay_hc_6));
    Odrv4 I__7229 (
            .O(N__35275),
            .I(measured_delay_hc_6));
    CascadeMux I__7228 (
            .O(N__35266),
            .I(N__35262));
    InMux I__7227 (
            .O(N__35265),
            .I(N__35259));
    InMux I__7226 (
            .O(N__35262),
            .I(N__35256));
    LocalMux I__7225 (
            .O(N__35259),
            .I(N__35251));
    LocalMux I__7224 (
            .O(N__35256),
            .I(N__35248));
    InMux I__7223 (
            .O(N__35255),
            .I(N__35245));
    InMux I__7222 (
            .O(N__35254),
            .I(N__35241));
    Span4Mux_v I__7221 (
            .O(N__35251),
            .I(N__35238));
    Span4Mux_h I__7220 (
            .O(N__35248),
            .I(N__35235));
    LocalMux I__7219 (
            .O(N__35245),
            .I(N__35232));
    InMux I__7218 (
            .O(N__35244),
            .I(N__35229));
    LocalMux I__7217 (
            .O(N__35241),
            .I(N__35226));
    Span4Mux_h I__7216 (
            .O(N__35238),
            .I(N__35219));
    Span4Mux_v I__7215 (
            .O(N__35235),
            .I(N__35219));
    Span4Mux_v I__7214 (
            .O(N__35232),
            .I(N__35219));
    LocalMux I__7213 (
            .O(N__35229),
            .I(measured_delay_hc_4));
    Odrv4 I__7212 (
            .O(N__35226),
            .I(measured_delay_hc_4));
    Odrv4 I__7211 (
            .O(N__35219),
            .I(measured_delay_hc_4));
    InMux I__7210 (
            .O(N__35212),
            .I(\current_shift_inst.timer_phase.counter_cry_17 ));
    InMux I__7209 (
            .O(N__35209),
            .I(\current_shift_inst.timer_phase.counter_cry_18 ));
    InMux I__7208 (
            .O(N__35206),
            .I(\current_shift_inst.timer_phase.counter_cry_19 ));
    InMux I__7207 (
            .O(N__35203),
            .I(\current_shift_inst.timer_phase.counter_cry_20 ));
    InMux I__7206 (
            .O(N__35200),
            .I(\current_shift_inst.timer_phase.counter_cry_21 ));
    InMux I__7205 (
            .O(N__35197),
            .I(\current_shift_inst.timer_phase.counter_cry_22 ));
    InMux I__7204 (
            .O(N__35194),
            .I(bfn_14_25_0_));
    InMux I__7203 (
            .O(N__35191),
            .I(\current_shift_inst.timer_phase.counter_cry_24 ));
    InMux I__7202 (
            .O(N__35188),
            .I(\current_shift_inst.timer_phase.counter_cry_25 ));
    InMux I__7201 (
            .O(N__35185),
            .I(\current_shift_inst.timer_phase.counter_cry_8 ));
    InMux I__7200 (
            .O(N__35182),
            .I(\current_shift_inst.timer_phase.counter_cry_9 ));
    InMux I__7199 (
            .O(N__35179),
            .I(\current_shift_inst.timer_phase.counter_cry_10 ));
    InMux I__7198 (
            .O(N__35176),
            .I(\current_shift_inst.timer_phase.counter_cry_11 ));
    InMux I__7197 (
            .O(N__35173),
            .I(\current_shift_inst.timer_phase.counter_cry_12 ));
    InMux I__7196 (
            .O(N__35170),
            .I(\current_shift_inst.timer_phase.counter_cry_13 ));
    InMux I__7195 (
            .O(N__35167),
            .I(\current_shift_inst.timer_phase.counter_cry_14 ));
    InMux I__7194 (
            .O(N__35164),
            .I(bfn_14_24_0_));
    InMux I__7193 (
            .O(N__35161),
            .I(\current_shift_inst.timer_phase.counter_cry_16 ));
    InMux I__7192 (
            .O(N__35158),
            .I(bfn_14_22_0_));
    InMux I__7191 (
            .O(N__35155),
            .I(\current_shift_inst.timer_phase.counter_cry_0 ));
    InMux I__7190 (
            .O(N__35152),
            .I(\current_shift_inst.timer_phase.counter_cry_1 ));
    InMux I__7189 (
            .O(N__35149),
            .I(\current_shift_inst.timer_phase.counter_cry_2 ));
    InMux I__7188 (
            .O(N__35146),
            .I(\current_shift_inst.timer_phase.counter_cry_3 ));
    InMux I__7187 (
            .O(N__35143),
            .I(\current_shift_inst.timer_phase.counter_cry_4 ));
    InMux I__7186 (
            .O(N__35140),
            .I(\current_shift_inst.timer_phase.counter_cry_5 ));
    InMux I__7185 (
            .O(N__35137),
            .I(\current_shift_inst.timer_phase.counter_cry_6 ));
    InMux I__7184 (
            .O(N__35134),
            .I(bfn_14_23_0_));
    CascadeMux I__7183 (
            .O(N__35131),
            .I(N__35127));
    InMux I__7182 (
            .O(N__35130),
            .I(N__35122));
    InMux I__7181 (
            .O(N__35127),
            .I(N__35122));
    LocalMux I__7180 (
            .O(N__35122),
            .I(N__35119));
    Span4Mux_v I__7179 (
            .O(N__35119),
            .I(N__35114));
    InMux I__7178 (
            .O(N__35118),
            .I(N__35111));
    InMux I__7177 (
            .O(N__35117),
            .I(N__35108));
    Span4Mux_v I__7176 (
            .O(N__35114),
            .I(N__35105));
    LocalMux I__7175 (
            .O(N__35111),
            .I(N__35102));
    LocalMux I__7174 (
            .O(N__35108),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    Odrv4 I__7173 (
            .O(N__35105),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    Odrv12 I__7172 (
            .O(N__35102),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    InMux I__7171 (
            .O(N__35095),
            .I(N__35092));
    LocalMux I__7170 (
            .O(N__35092),
            .I(N__35087));
    CascadeMux I__7169 (
            .O(N__35091),
            .I(N__35084));
    CascadeMux I__7168 (
            .O(N__35090),
            .I(N__35081));
    Span4Mux_v I__7167 (
            .O(N__35087),
            .I(N__35077));
    InMux I__7166 (
            .O(N__35084),
            .I(N__35074));
    InMux I__7165 (
            .O(N__35081),
            .I(N__35069));
    InMux I__7164 (
            .O(N__35080),
            .I(N__35069));
    Span4Mux_v I__7163 (
            .O(N__35077),
            .I(N__35066));
    LocalMux I__7162 (
            .O(N__35074),
            .I(N__35063));
    LocalMux I__7161 (
            .O(N__35069),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    Odrv4 I__7160 (
            .O(N__35066),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    Odrv12 I__7159 (
            .O(N__35063),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    CascadeMux I__7158 (
            .O(N__35056),
            .I(N__35051));
    InMux I__7157 (
            .O(N__35055),
            .I(N__35047));
    InMux I__7156 (
            .O(N__35054),
            .I(N__35044));
    InMux I__7155 (
            .O(N__35051),
            .I(N__35039));
    InMux I__7154 (
            .O(N__35050),
            .I(N__35039));
    LocalMux I__7153 (
            .O(N__35047),
            .I(N__35036));
    LocalMux I__7152 (
            .O(N__35044),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    LocalMux I__7151 (
            .O(N__35039),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    Odrv12 I__7150 (
            .O(N__35036),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    CascadeMux I__7149 (
            .O(N__35029),
            .I(N__35025));
    InMux I__7148 (
            .O(N__35028),
            .I(N__35020));
    InMux I__7147 (
            .O(N__35025),
            .I(N__35017));
    InMux I__7146 (
            .O(N__35024),
            .I(N__35012));
    InMux I__7145 (
            .O(N__35023),
            .I(N__35012));
    LocalMux I__7144 (
            .O(N__35020),
            .I(N__35009));
    LocalMux I__7143 (
            .O(N__35017),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    LocalMux I__7142 (
            .O(N__35012),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    Odrv12 I__7141 (
            .O(N__35009),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    CascadeMux I__7140 (
            .O(N__35002),
            .I(N__34998));
    CascadeMux I__7139 (
            .O(N__35001),
            .I(N__34995));
    InMux I__7138 (
            .O(N__34998),
            .I(N__34992));
    InMux I__7137 (
            .O(N__34995),
            .I(N__34989));
    LocalMux I__7136 (
            .O(N__34992),
            .I(N__34986));
    LocalMux I__7135 (
            .O(N__34989),
            .I(N__34981));
    Span4Mux_h I__7134 (
            .O(N__34986),
            .I(N__34978));
    InMux I__7133 (
            .O(N__34985),
            .I(N__34975));
    InMux I__7132 (
            .O(N__34984),
            .I(N__34972));
    Span4Mux_v I__7131 (
            .O(N__34981),
            .I(N__34969));
    Odrv4 I__7130 (
            .O(N__34978),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    LocalMux I__7129 (
            .O(N__34975),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    LocalMux I__7128 (
            .O(N__34972),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    Odrv4 I__7127 (
            .O(N__34969),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    InMux I__7126 (
            .O(N__34960),
            .I(N__34955));
    InMux I__7125 (
            .O(N__34959),
            .I(N__34952));
    InMux I__7124 (
            .O(N__34958),
            .I(N__34949));
    LocalMux I__7123 (
            .O(N__34955),
            .I(N__34946));
    LocalMux I__7122 (
            .O(N__34952),
            .I(N__34943));
    LocalMux I__7121 (
            .O(N__34949),
            .I(N__34940));
    Span4Mux_h I__7120 (
            .O(N__34946),
            .I(N__34937));
    Span4Mux_h I__7119 (
            .O(N__34943),
            .I(N__34932));
    Span4Mux_v I__7118 (
            .O(N__34940),
            .I(N__34932));
    Odrv4 I__7117 (
            .O(N__34937),
            .I(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ));
    Odrv4 I__7116 (
            .O(N__34932),
            .I(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ));
    InMux I__7115 (
            .O(N__34927),
            .I(N__34923));
    CascadeMux I__7114 (
            .O(N__34926),
            .I(N__34920));
    LocalMux I__7113 (
            .O(N__34923),
            .I(N__34917));
    InMux I__7112 (
            .O(N__34920),
            .I(N__34914));
    Span4Mux_h I__7111 (
            .O(N__34917),
            .I(N__34908));
    LocalMux I__7110 (
            .O(N__34914),
            .I(N__34908));
    InMux I__7109 (
            .O(N__34913),
            .I(N__34905));
    Span4Mux_v I__7108 (
            .O(N__34908),
            .I(N__34902));
    LocalMux I__7107 (
            .O(N__34905),
            .I(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ));
    Odrv4 I__7106 (
            .O(N__34902),
            .I(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ));
    InMux I__7105 (
            .O(N__34897),
            .I(\current_shift_inst.z_cry_30 ));
    InMux I__7104 (
            .O(N__34894),
            .I(N__34890));
    InMux I__7103 (
            .O(N__34893),
            .I(N__34887));
    LocalMux I__7102 (
            .O(N__34890),
            .I(N__34884));
    LocalMux I__7101 (
            .O(N__34887),
            .I(N__34881));
    Span4Mux_h I__7100 (
            .O(N__34884),
            .I(N__34876));
    Span4Mux_h I__7099 (
            .O(N__34881),
            .I(N__34876));
    Odrv4 I__7098 (
            .O(N__34876),
            .I(\current_shift_inst.z_31 ));
    CascadeMux I__7097 (
            .O(N__34873),
            .I(N__34870));
    InMux I__7096 (
            .O(N__34870),
            .I(N__34867));
    LocalMux I__7095 (
            .O(N__34867),
            .I(N__34862));
    InMux I__7094 (
            .O(N__34866),
            .I(N__34858));
    InMux I__7093 (
            .O(N__34865),
            .I(N__34855));
    Span4Mux_h I__7092 (
            .O(N__34862),
            .I(N__34852));
    InMux I__7091 (
            .O(N__34861),
            .I(N__34849));
    LocalMux I__7090 (
            .O(N__34858),
            .I(N__34846));
    LocalMux I__7089 (
            .O(N__34855),
            .I(N__34843));
    Odrv4 I__7088 (
            .O(N__34852),
            .I(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ));
    LocalMux I__7087 (
            .O(N__34849),
            .I(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ));
    Odrv12 I__7086 (
            .O(N__34846),
            .I(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ));
    Odrv12 I__7085 (
            .O(N__34843),
            .I(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ));
    InMux I__7084 (
            .O(N__34834),
            .I(N__34830));
    InMux I__7083 (
            .O(N__34833),
            .I(N__34826));
    LocalMux I__7082 (
            .O(N__34830),
            .I(N__34823));
    InMux I__7081 (
            .O(N__34829),
            .I(N__34820));
    LocalMux I__7080 (
            .O(N__34826),
            .I(N__34812));
    Span4Mux_h I__7079 (
            .O(N__34823),
            .I(N__34812));
    LocalMux I__7078 (
            .O(N__34820),
            .I(N__34812));
    InMux I__7077 (
            .O(N__34819),
            .I(N__34809));
    Span4Mux_v I__7076 (
            .O(N__34812),
            .I(N__34806));
    LocalMux I__7075 (
            .O(N__34809),
            .I(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ));
    Odrv4 I__7074 (
            .O(N__34806),
            .I(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ));
    CascadeMux I__7073 (
            .O(N__34801),
            .I(N__34798));
    InMux I__7072 (
            .O(N__34798),
            .I(N__34795));
    LocalMux I__7071 (
            .O(N__34795),
            .I(N__34791));
    CascadeMux I__7070 (
            .O(N__34794),
            .I(N__34788));
    Span4Mux_h I__7069 (
            .O(N__34791),
            .I(N__34785));
    InMux I__7068 (
            .O(N__34788),
            .I(N__34780));
    Span4Mux_v I__7067 (
            .O(N__34785),
            .I(N__34777));
    InMux I__7066 (
            .O(N__34784),
            .I(N__34774));
    InMux I__7065 (
            .O(N__34783),
            .I(N__34771));
    LocalMux I__7064 (
            .O(N__34780),
            .I(N__34768));
    Odrv4 I__7063 (
            .O(N__34777),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    LocalMux I__7062 (
            .O(N__34774),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    LocalMux I__7061 (
            .O(N__34771),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    Odrv12 I__7060 (
            .O(N__34768),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    CascadeMux I__7059 (
            .O(N__34759),
            .I(N__34756));
    InMux I__7058 (
            .O(N__34756),
            .I(N__34750));
    InMux I__7057 (
            .O(N__34755),
            .I(N__34750));
    LocalMux I__7056 (
            .O(N__34750),
            .I(N__34745));
    InMux I__7055 (
            .O(N__34749),
            .I(N__34742));
    InMux I__7054 (
            .O(N__34748),
            .I(N__34739));
    Span4Mux_h I__7053 (
            .O(N__34745),
            .I(N__34736));
    LocalMux I__7052 (
            .O(N__34742),
            .I(N__34733));
    LocalMux I__7051 (
            .O(N__34739),
            .I(N__34730));
    Odrv4 I__7050 (
            .O(N__34736),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    Odrv12 I__7049 (
            .O(N__34733),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    Odrv12 I__7048 (
            .O(N__34730),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    InMux I__7047 (
            .O(N__34723),
            .I(N__34719));
    CascadeMux I__7046 (
            .O(N__34722),
            .I(N__34715));
    LocalMux I__7045 (
            .O(N__34719),
            .I(N__34712));
    CascadeMux I__7044 (
            .O(N__34718),
            .I(N__34709));
    InMux I__7043 (
            .O(N__34715),
            .I(N__34705));
    Span4Mux_h I__7042 (
            .O(N__34712),
            .I(N__34702));
    InMux I__7041 (
            .O(N__34709),
            .I(N__34697));
    InMux I__7040 (
            .O(N__34708),
            .I(N__34697));
    LocalMux I__7039 (
            .O(N__34705),
            .I(N__34694));
    Odrv4 I__7038 (
            .O(N__34702),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    LocalMux I__7037 (
            .O(N__34697),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    Odrv12 I__7036 (
            .O(N__34694),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    CascadeMux I__7035 (
            .O(N__34687),
            .I(N__34682));
    CascadeMux I__7034 (
            .O(N__34686),
            .I(N__34679));
    InMux I__7033 (
            .O(N__34685),
            .I(N__34676));
    InMux I__7032 (
            .O(N__34682),
            .I(N__34673));
    InMux I__7031 (
            .O(N__34679),
            .I(N__34670));
    LocalMux I__7030 (
            .O(N__34676),
            .I(N__34666));
    LocalMux I__7029 (
            .O(N__34673),
            .I(N__34663));
    LocalMux I__7028 (
            .O(N__34670),
            .I(N__34660));
    InMux I__7027 (
            .O(N__34669),
            .I(N__34657));
    Span4Mux_h I__7026 (
            .O(N__34666),
            .I(N__34654));
    Span4Mux_v I__7025 (
            .O(N__34663),
            .I(N__34651));
    Odrv12 I__7024 (
            .O(N__34660),
            .I(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ));
    LocalMux I__7023 (
            .O(N__34657),
            .I(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ));
    Odrv4 I__7022 (
            .O(N__34654),
            .I(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ));
    Odrv4 I__7021 (
            .O(N__34651),
            .I(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ));
    CascadeMux I__7020 (
            .O(N__34642),
            .I(N__34639));
    InMux I__7019 (
            .O(N__34639),
            .I(N__34636));
    LocalMux I__7018 (
            .O(N__34636),
            .I(N__34632));
    CascadeMux I__7017 (
            .O(N__34635),
            .I(N__34629));
    Span4Mux_v I__7016 (
            .O(N__34632),
            .I(N__34624));
    InMux I__7015 (
            .O(N__34629),
            .I(N__34621));
    InMux I__7014 (
            .O(N__34628),
            .I(N__34616));
    InMux I__7013 (
            .O(N__34627),
            .I(N__34616));
    Span4Mux_h I__7012 (
            .O(N__34624),
            .I(N__34611));
    LocalMux I__7011 (
            .O(N__34621),
            .I(N__34611));
    LocalMux I__7010 (
            .O(N__34616),
            .I(N__34608));
    Span4Mux_v I__7009 (
            .O(N__34611),
            .I(N__34605));
    Odrv12 I__7008 (
            .O(N__34608),
            .I(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ));
    Odrv4 I__7007 (
            .O(N__34605),
            .I(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ));
    InMux I__7006 (
            .O(N__34600),
            .I(N__34597));
    LocalMux I__7005 (
            .O(N__34597),
            .I(N__34591));
    InMux I__7004 (
            .O(N__34596),
            .I(N__34586));
    InMux I__7003 (
            .O(N__34595),
            .I(N__34586));
    CascadeMux I__7002 (
            .O(N__34594),
            .I(N__34583));
    Span4Mux_v I__7001 (
            .O(N__34591),
            .I(N__34580));
    LocalMux I__7000 (
            .O(N__34586),
            .I(N__34577));
    InMux I__6999 (
            .O(N__34583),
            .I(N__34574));
    Span4Mux_h I__6998 (
            .O(N__34580),
            .I(N__34571));
    Span4Mux_h I__6997 (
            .O(N__34577),
            .I(N__34568));
    LocalMux I__6996 (
            .O(N__34574),
            .I(N__34565));
    Odrv4 I__6995 (
            .O(N__34571),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    Odrv4 I__6994 (
            .O(N__34568),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    Odrv12 I__6993 (
            .O(N__34565),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    InMux I__6992 (
            .O(N__34558),
            .I(N__34555));
    LocalMux I__6991 (
            .O(N__34555),
            .I(N__34551));
    InMux I__6990 (
            .O(N__34554),
            .I(N__34546));
    Span4Mux_h I__6989 (
            .O(N__34551),
            .I(N__34543));
    InMux I__6988 (
            .O(N__34550),
            .I(N__34540));
    InMux I__6987 (
            .O(N__34549),
            .I(N__34537));
    LocalMux I__6986 (
            .O(N__34546),
            .I(N__34534));
    Sp12to4 I__6985 (
            .O(N__34543),
            .I(N__34529));
    LocalMux I__6984 (
            .O(N__34540),
            .I(N__34529));
    LocalMux I__6983 (
            .O(N__34537),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    Odrv12 I__6982 (
            .O(N__34534),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    Odrv12 I__6981 (
            .O(N__34529),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    InMux I__6980 (
            .O(N__34522),
            .I(N__34516));
    InMux I__6979 (
            .O(N__34521),
            .I(N__34516));
    LocalMux I__6978 (
            .O(N__34516),
            .I(N__34512));
    InMux I__6977 (
            .O(N__34515),
            .I(N__34509));
    Span4Mux_h I__6976 (
            .O(N__34512),
            .I(N__34506));
    LocalMux I__6975 (
            .O(N__34509),
            .I(N__34500));
    Span4Mux_v I__6974 (
            .O(N__34506),
            .I(N__34500));
    InMux I__6973 (
            .O(N__34505),
            .I(N__34497));
    Span4Mux_v I__6972 (
            .O(N__34500),
            .I(N__34494));
    LocalMux I__6971 (
            .O(N__34497),
            .I(N__34491));
    Odrv4 I__6970 (
            .O(N__34494),
            .I(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ));
    Odrv12 I__6969 (
            .O(N__34491),
            .I(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ));
    InMux I__6968 (
            .O(N__34486),
            .I(N__34483));
    LocalMux I__6967 (
            .O(N__34483),
            .I(N__34480));
    Span4Mux_v I__6966 (
            .O(N__34480),
            .I(N__34475));
    InMux I__6965 (
            .O(N__34479),
            .I(N__34472));
    CascadeMux I__6964 (
            .O(N__34478),
            .I(N__34469));
    Span4Mux_h I__6963 (
            .O(N__34475),
            .I(N__34463));
    LocalMux I__6962 (
            .O(N__34472),
            .I(N__34463));
    InMux I__6961 (
            .O(N__34469),
            .I(N__34460));
    InMux I__6960 (
            .O(N__34468),
            .I(N__34457));
    Span4Mux_v I__6959 (
            .O(N__34463),
            .I(N__34454));
    LocalMux I__6958 (
            .O(N__34460),
            .I(N__34451));
    LocalMux I__6957 (
            .O(N__34457),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    Odrv4 I__6956 (
            .O(N__34454),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    Odrv12 I__6955 (
            .O(N__34451),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    CascadeMux I__6954 (
            .O(N__34444),
            .I(N__34441));
    InMux I__6953 (
            .O(N__34441),
            .I(N__34434));
    InMux I__6952 (
            .O(N__34440),
            .I(N__34434));
    InMux I__6951 (
            .O(N__34439),
            .I(N__34431));
    LocalMux I__6950 (
            .O(N__34434),
            .I(N__34428));
    LocalMux I__6949 (
            .O(N__34431),
            .I(N__34425));
    Span4Mux_h I__6948 (
            .O(N__34428),
            .I(N__34422));
    Span4Mux_h I__6947 (
            .O(N__34425),
            .I(N__34418));
    Span4Mux_h I__6946 (
            .O(N__34422),
            .I(N__34415));
    InMux I__6945 (
            .O(N__34421),
            .I(N__34412));
    Sp12to4 I__6944 (
            .O(N__34418),
            .I(N__34405));
    Sp12to4 I__6943 (
            .O(N__34415),
            .I(N__34405));
    LocalMux I__6942 (
            .O(N__34412),
            .I(N__34405));
    Odrv12 I__6941 (
            .O(N__34405),
            .I(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ));
    CascadeMux I__6940 (
            .O(N__34402),
            .I(N__34397));
    InMux I__6939 (
            .O(N__34401),
            .I(N__34394));
    InMux I__6938 (
            .O(N__34400),
            .I(N__34390));
    InMux I__6937 (
            .O(N__34397),
            .I(N__34387));
    LocalMux I__6936 (
            .O(N__34394),
            .I(N__34384));
    CascadeMux I__6935 (
            .O(N__34393),
            .I(N__34381));
    LocalMux I__6934 (
            .O(N__34390),
            .I(N__34378));
    LocalMux I__6933 (
            .O(N__34387),
            .I(N__34373));
    Span4Mux_v I__6932 (
            .O(N__34384),
            .I(N__34373));
    InMux I__6931 (
            .O(N__34381),
            .I(N__34370));
    Span4Mux_h I__6930 (
            .O(N__34378),
            .I(N__34363));
    Span4Mux_h I__6929 (
            .O(N__34373),
            .I(N__34363));
    LocalMux I__6928 (
            .O(N__34370),
            .I(N__34363));
    Span4Mux_v I__6927 (
            .O(N__34363),
            .I(N__34360));
    Odrv4 I__6926 (
            .O(N__34360),
            .I(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ));
    InMux I__6925 (
            .O(N__34357),
            .I(N__34352));
    CascadeMux I__6924 (
            .O(N__34356),
            .I(N__34349));
    InMux I__6923 (
            .O(N__34355),
            .I(N__34346));
    LocalMux I__6922 (
            .O(N__34352),
            .I(N__34343));
    InMux I__6921 (
            .O(N__34349),
            .I(N__34340));
    LocalMux I__6920 (
            .O(N__34346),
            .I(N__34336));
    Span4Mux_v I__6919 (
            .O(N__34343),
            .I(N__34333));
    LocalMux I__6918 (
            .O(N__34340),
            .I(N__34330));
    InMux I__6917 (
            .O(N__34339),
            .I(N__34327));
    Span4Mux_v I__6916 (
            .O(N__34336),
            .I(N__34324));
    Span4Mux_h I__6915 (
            .O(N__34333),
            .I(N__34319));
    Span4Mux_v I__6914 (
            .O(N__34330),
            .I(N__34319));
    LocalMux I__6913 (
            .O(N__34327),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    Odrv4 I__6912 (
            .O(N__34324),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    Odrv4 I__6911 (
            .O(N__34319),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    InMux I__6910 (
            .O(N__34312),
            .I(N__34308));
    CascadeMux I__6909 (
            .O(N__34311),
            .I(N__34304));
    LocalMux I__6908 (
            .O(N__34308),
            .I(N__34300));
    InMux I__6907 (
            .O(N__34307),
            .I(N__34297));
    InMux I__6906 (
            .O(N__34304),
            .I(N__34294));
    InMux I__6905 (
            .O(N__34303),
            .I(N__34291));
    Span4Mux_v I__6904 (
            .O(N__34300),
            .I(N__34288));
    LocalMux I__6903 (
            .O(N__34297),
            .I(N__34285));
    LocalMux I__6902 (
            .O(N__34294),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    LocalMux I__6901 (
            .O(N__34291),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    Odrv4 I__6900 (
            .O(N__34288),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    Odrv12 I__6899 (
            .O(N__34285),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    InMux I__6898 (
            .O(N__34276),
            .I(N__34272));
    InMux I__6897 (
            .O(N__34275),
            .I(N__34269));
    LocalMux I__6896 (
            .O(N__34272),
            .I(N__34265));
    LocalMux I__6895 (
            .O(N__34269),
            .I(N__34262));
    CascadeMux I__6894 (
            .O(N__34268),
            .I(N__34259));
    Span4Mux_v I__6893 (
            .O(N__34265),
            .I(N__34253));
    Span4Mux_v I__6892 (
            .O(N__34262),
            .I(N__34253));
    InMux I__6891 (
            .O(N__34259),
            .I(N__34250));
    InMux I__6890 (
            .O(N__34258),
            .I(N__34247));
    Span4Mux_h I__6889 (
            .O(N__34253),
            .I(N__34244));
    LocalMux I__6888 (
            .O(N__34250),
            .I(N__34241));
    LocalMux I__6887 (
            .O(N__34247),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    Odrv4 I__6886 (
            .O(N__34244),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    Odrv12 I__6885 (
            .O(N__34241),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    InMux I__6884 (
            .O(N__34234),
            .I(N__34229));
    CascadeMux I__6883 (
            .O(N__34233),
            .I(N__34226));
    InMux I__6882 (
            .O(N__34232),
            .I(N__34223));
    LocalMux I__6881 (
            .O(N__34229),
            .I(N__34220));
    InMux I__6880 (
            .O(N__34226),
            .I(N__34216));
    LocalMux I__6879 (
            .O(N__34223),
            .I(N__34211));
    Span4Mux_v I__6878 (
            .O(N__34220),
            .I(N__34211));
    InMux I__6877 (
            .O(N__34219),
            .I(N__34208));
    LocalMux I__6876 (
            .O(N__34216),
            .I(N__34205));
    Span4Mux_h I__6875 (
            .O(N__34211),
            .I(N__34202));
    LocalMux I__6874 (
            .O(N__34208),
            .I(N__34199));
    Odrv4 I__6873 (
            .O(N__34205),
            .I(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ));
    Odrv4 I__6872 (
            .O(N__34202),
            .I(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ));
    Odrv12 I__6871 (
            .O(N__34199),
            .I(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ));
    InMux I__6870 (
            .O(N__34192),
            .I(\current_shift_inst.un4_control_input_cry_30 ));
    CascadeMux I__6869 (
            .O(N__34189),
            .I(N__34186));
    InMux I__6868 (
            .O(N__34186),
            .I(N__34183));
    LocalMux I__6867 (
            .O(N__34183),
            .I(N__34180));
    Span4Mux_v I__6866 (
            .O(N__34180),
            .I(N__34177));
    Span4Mux_h I__6865 (
            .O(N__34177),
            .I(N__34174));
    Odrv4 I__6864 (
            .O(N__34174),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ));
    CascadeMux I__6863 (
            .O(N__34171),
            .I(N__34168));
    InMux I__6862 (
            .O(N__34168),
            .I(N__34165));
    LocalMux I__6861 (
            .O(N__34165),
            .I(N__34162));
    Span4Mux_v I__6860 (
            .O(N__34162),
            .I(N__34158));
    InMux I__6859 (
            .O(N__34161),
            .I(N__34155));
    Span4Mux_h I__6858 (
            .O(N__34158),
            .I(N__34150));
    LocalMux I__6857 (
            .O(N__34155),
            .I(N__34150));
    Span4Mux_v I__6856 (
            .O(N__34150),
            .I(N__34147));
    Odrv4 I__6855 (
            .O(N__34147),
            .I(\current_shift_inst.un38_control_input_0 ));
    InMux I__6854 (
            .O(N__34144),
            .I(N__34140));
    CascadeMux I__6853 (
            .O(N__34143),
            .I(N__34137));
    LocalMux I__6852 (
            .O(N__34140),
            .I(N__34133));
    InMux I__6851 (
            .O(N__34137),
            .I(N__34130));
    InMux I__6850 (
            .O(N__34136),
            .I(N__34127));
    Span4Mux_v I__6849 (
            .O(N__34133),
            .I(N__34122));
    LocalMux I__6848 (
            .O(N__34130),
            .I(N__34122));
    LocalMux I__6847 (
            .O(N__34127),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    Odrv4 I__6846 (
            .O(N__34122),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    CascadeMux I__6845 (
            .O(N__34117),
            .I(N__34114));
    InMux I__6844 (
            .O(N__34114),
            .I(N__34111));
    LocalMux I__6843 (
            .O(N__34111),
            .I(G_407));
    InMux I__6842 (
            .O(N__34108),
            .I(N__34104));
    InMux I__6841 (
            .O(N__34107),
            .I(N__34101));
    LocalMux I__6840 (
            .O(N__34104),
            .I(N__34096));
    LocalMux I__6839 (
            .O(N__34101),
            .I(N__34096));
    Span4Mux_v I__6838 (
            .O(N__34096),
            .I(N__34092));
    InMux I__6837 (
            .O(N__34095),
            .I(N__34089));
    Span4Mux_h I__6836 (
            .O(N__34092),
            .I(N__34084));
    LocalMux I__6835 (
            .O(N__34089),
            .I(N__34084));
    Span4Mux_v I__6834 (
            .O(N__34084),
            .I(N__34081));
    Odrv4 I__6833 (
            .O(N__34081),
            .I(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ));
    CascadeMux I__6832 (
            .O(N__34078),
            .I(N__34075));
    InMux I__6831 (
            .O(N__34075),
            .I(N__34072));
    LocalMux I__6830 (
            .O(N__34072),
            .I(G_406));
    InMux I__6829 (
            .O(N__34069),
            .I(N__34066));
    LocalMux I__6828 (
            .O(N__34066),
            .I(N__34062));
    InMux I__6827 (
            .O(N__34065),
            .I(N__34059));
    Span4Mux_v I__6826 (
            .O(N__34062),
            .I(N__34053));
    LocalMux I__6825 (
            .O(N__34059),
            .I(N__34053));
    CascadeMux I__6824 (
            .O(N__34058),
            .I(N__34050));
    Span4Mux_h I__6823 (
            .O(N__34053),
            .I(N__34047));
    InMux I__6822 (
            .O(N__34050),
            .I(N__34044));
    Span4Mux_v I__6821 (
            .O(N__34047),
            .I(N__34041));
    LocalMux I__6820 (
            .O(N__34044),
            .I(N__34038));
    Odrv4 I__6819 (
            .O(N__34041),
            .I(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ));
    Odrv12 I__6818 (
            .O(N__34038),
            .I(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ));
    InMux I__6817 (
            .O(N__34033),
            .I(N__34029));
    CascadeMux I__6816 (
            .O(N__34032),
            .I(N__34026));
    LocalMux I__6815 (
            .O(N__34029),
            .I(N__34023));
    InMux I__6814 (
            .O(N__34026),
            .I(N__34020));
    Span4Mux_h I__6813 (
            .O(N__34023),
            .I(N__34017));
    LocalMux I__6812 (
            .O(N__34020),
            .I(N__34014));
    Span4Mux_v I__6811 (
            .O(N__34017),
            .I(N__34009));
    Span4Mux_v I__6810 (
            .O(N__34014),
            .I(N__34009));
    Odrv4 I__6809 (
            .O(N__34009),
            .I(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ));
    CascadeMux I__6808 (
            .O(N__34006),
            .I(N__34003));
    InMux I__6807 (
            .O(N__34003),
            .I(N__33996));
    InMux I__6806 (
            .O(N__34002),
            .I(N__33996));
    InMux I__6805 (
            .O(N__34001),
            .I(N__33993));
    LocalMux I__6804 (
            .O(N__33996),
            .I(N__33990));
    LocalMux I__6803 (
            .O(N__33993),
            .I(N__33986));
    Span4Mux_v I__6802 (
            .O(N__33990),
            .I(N__33983));
    InMux I__6801 (
            .O(N__33989),
            .I(N__33980));
    Span4Mux_v I__6800 (
            .O(N__33986),
            .I(N__33977));
    Span4Mux_h I__6799 (
            .O(N__33983),
            .I(N__33974));
    LocalMux I__6798 (
            .O(N__33980),
            .I(N__33971));
    Odrv4 I__6797 (
            .O(N__33977),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    Odrv4 I__6796 (
            .O(N__33974),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    Odrv12 I__6795 (
            .O(N__33971),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    CascadeMux I__6794 (
            .O(N__33964),
            .I(N__33961));
    InMux I__6793 (
            .O(N__33961),
            .I(N__33957));
    InMux I__6792 (
            .O(N__33960),
            .I(N__33954));
    LocalMux I__6791 (
            .O(N__33957),
            .I(N__33950));
    LocalMux I__6790 (
            .O(N__33954),
            .I(N__33947));
    InMux I__6789 (
            .O(N__33953),
            .I(N__33944));
    Span4Mux_h I__6788 (
            .O(N__33950),
            .I(N__33936));
    Span4Mux_v I__6787 (
            .O(N__33947),
            .I(N__33936));
    LocalMux I__6786 (
            .O(N__33944),
            .I(N__33936));
    CascadeMux I__6785 (
            .O(N__33943),
            .I(N__33933));
    Span4Mux_v I__6784 (
            .O(N__33936),
            .I(N__33930));
    InMux I__6783 (
            .O(N__33933),
            .I(N__33927));
    Span4Mux_h I__6782 (
            .O(N__33930),
            .I(N__33924));
    LocalMux I__6781 (
            .O(N__33927),
            .I(N__33921));
    Odrv4 I__6780 (
            .O(N__33924),
            .I(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ));
    Odrv12 I__6779 (
            .O(N__33921),
            .I(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ));
    InMux I__6778 (
            .O(N__33916),
            .I(N__33909));
    InMux I__6777 (
            .O(N__33915),
            .I(N__33909));
    InMux I__6776 (
            .O(N__33914),
            .I(N__33906));
    LocalMux I__6775 (
            .O(N__33909),
            .I(N__33903));
    LocalMux I__6774 (
            .O(N__33906),
            .I(N__33898));
    Span4Mux_h I__6773 (
            .O(N__33903),
            .I(N__33898));
    Span4Mux_v I__6772 (
            .O(N__33898),
            .I(N__33894));
    InMux I__6771 (
            .O(N__33897),
            .I(N__33891));
    Span4Mux_v I__6770 (
            .O(N__33894),
            .I(N__33888));
    LocalMux I__6769 (
            .O(N__33891),
            .I(N__33885));
    Odrv4 I__6768 (
            .O(N__33888),
            .I(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ));
    Odrv12 I__6767 (
            .O(N__33885),
            .I(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ));
    InMux I__6766 (
            .O(N__33880),
            .I(\current_shift_inst.un4_control_input_cry_21 ));
    InMux I__6765 (
            .O(N__33877),
            .I(\current_shift_inst.un4_control_input_cry_22 ));
    InMux I__6764 (
            .O(N__33874),
            .I(\current_shift_inst.un4_control_input_cry_23 ));
    InMux I__6763 (
            .O(N__33871),
            .I(bfn_14_17_0_));
    InMux I__6762 (
            .O(N__33868),
            .I(\current_shift_inst.un4_control_input_cry_25 ));
    InMux I__6761 (
            .O(N__33865),
            .I(\current_shift_inst.un4_control_input_cry_26 ));
    InMux I__6760 (
            .O(N__33862),
            .I(\current_shift_inst.un4_control_input_cry_27 ));
    InMux I__6759 (
            .O(N__33859),
            .I(\current_shift_inst.un4_control_input_cry_28 ));
    InMux I__6758 (
            .O(N__33856),
            .I(\current_shift_inst.un4_control_input_cry_29 ));
    InMux I__6757 (
            .O(N__33853),
            .I(\current_shift_inst.un4_control_input_cry_12 ));
    InMux I__6756 (
            .O(N__33850),
            .I(\current_shift_inst.un4_control_input_cry_13 ));
    InMux I__6755 (
            .O(N__33847),
            .I(\current_shift_inst.un4_control_input_cry_14 ));
    InMux I__6754 (
            .O(N__33844),
            .I(\current_shift_inst.un4_control_input_cry_15 ));
    InMux I__6753 (
            .O(N__33841),
            .I(bfn_14_16_0_));
    InMux I__6752 (
            .O(N__33838),
            .I(\current_shift_inst.un4_control_input_cry_17 ));
    InMux I__6751 (
            .O(N__33835),
            .I(\current_shift_inst.un4_control_input_cry_18 ));
    InMux I__6750 (
            .O(N__33832),
            .I(\current_shift_inst.un4_control_input_cry_19 ));
    InMux I__6749 (
            .O(N__33829),
            .I(\current_shift_inst.un4_control_input_cry_20 ));
    InMux I__6748 (
            .O(N__33826),
            .I(\current_shift_inst.un4_control_input_cry_3 ));
    InMux I__6747 (
            .O(N__33823),
            .I(\current_shift_inst.un4_control_input_cry_4 ));
    InMux I__6746 (
            .O(N__33820),
            .I(\current_shift_inst.un4_control_input_cry_5 ));
    InMux I__6745 (
            .O(N__33817),
            .I(\current_shift_inst.un4_control_input_cry_6 ));
    InMux I__6744 (
            .O(N__33814),
            .I(\current_shift_inst.un4_control_input_cry_7 ));
    InMux I__6743 (
            .O(N__33811),
            .I(bfn_14_15_0_));
    InMux I__6742 (
            .O(N__33808),
            .I(\current_shift_inst.un4_control_input_cry_9 ));
    InMux I__6741 (
            .O(N__33805),
            .I(\current_shift_inst.un4_control_input_cry_10 ));
    InMux I__6740 (
            .O(N__33802),
            .I(\current_shift_inst.un4_control_input_cry_11 ));
    InMux I__6739 (
            .O(N__33799),
            .I(bfn_14_13_0_));
    InMux I__6738 (
            .O(N__33796),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__6737 (
            .O(N__33793),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__6736 (
            .O(N__33790),
            .I(N__33787));
    LocalMux I__6735 (
            .O(N__33787),
            .I(N__33784));
    Odrv4 I__6734 (
            .O(N__33784),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ));
    InMux I__6733 (
            .O(N__33781),
            .I(N__33776));
    InMux I__6732 (
            .O(N__33780),
            .I(N__33773));
    InMux I__6731 (
            .O(N__33779),
            .I(N__33770));
    LocalMux I__6730 (
            .O(N__33776),
            .I(N__33767));
    LocalMux I__6729 (
            .O(N__33773),
            .I(N__33761));
    LocalMux I__6728 (
            .O(N__33770),
            .I(N__33761));
    Span4Mux_v I__6727 (
            .O(N__33767),
            .I(N__33758));
    InMux I__6726 (
            .O(N__33766),
            .I(N__33755));
    Span4Mux_h I__6725 (
            .O(N__33761),
            .I(N__33752));
    Span4Mux_h I__6724 (
            .O(N__33758),
            .I(N__33749));
    LocalMux I__6723 (
            .O(N__33755),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv4 I__6722 (
            .O(N__33752),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv4 I__6721 (
            .O(N__33749),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__6720 (
            .O(N__33742),
            .I(N__33739));
    LocalMux I__6719 (
            .O(N__33739),
            .I(\current_shift_inst.un4_control_input_axb_1 ));
    InMux I__6718 (
            .O(N__33736),
            .I(N__33733));
    LocalMux I__6717 (
            .O(N__33733),
            .I(\current_shift_inst.un4_control_input_axb_2 ));
    InMux I__6716 (
            .O(N__33730),
            .I(\current_shift_inst.un4_control_input_cry_1 ));
    InMux I__6715 (
            .O(N__33727),
            .I(N__33724));
    LocalMux I__6714 (
            .O(N__33724),
            .I(\current_shift_inst.un4_control_input_axb_3 ));
    InMux I__6713 (
            .O(N__33721),
            .I(\current_shift_inst.un4_control_input_cry_2 ));
    InMux I__6712 (
            .O(N__33718),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__6711 (
            .O(N__33715),
            .I(bfn_14_12_0_));
    InMux I__6710 (
            .O(N__33712),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__6709 (
            .O(N__33709),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__6708 (
            .O(N__33706),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__6707 (
            .O(N__33703),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__6706 (
            .O(N__33700),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__6705 (
            .O(N__33697),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__6704 (
            .O(N__33694),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ));
    CascadeMux I__6703 (
            .O(N__33691),
            .I(\phase_controller_slave.stoper_tr.time_passed11_cascade_ ));
    InMux I__6702 (
            .O(N__33688),
            .I(N__33685));
    LocalMux I__6701 (
            .O(N__33685),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    InMux I__6700 (
            .O(N__33682),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__6699 (
            .O(N__33679),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__6698 (
            .O(N__33676),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__6697 (
            .O(N__33673),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__6696 (
            .O(N__33670),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__6695 (
            .O(N__33667),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ));
    IoInMux I__6694 (
            .O(N__33664),
            .I(N__33661));
    LocalMux I__6693 (
            .O(N__33661),
            .I(N__33658));
    Odrv12 I__6692 (
            .O(N__33658),
            .I(s2_phy_c));
    CascadeMux I__6691 (
            .O(N__33655),
            .I(N__33652));
    InMux I__6690 (
            .O(N__33652),
            .I(N__33640));
    InMux I__6689 (
            .O(N__33651),
            .I(N__33640));
    InMux I__6688 (
            .O(N__33650),
            .I(N__33635));
    InMux I__6687 (
            .O(N__33649),
            .I(N__33635));
    CascadeMux I__6686 (
            .O(N__33648),
            .I(N__33629));
    CascadeMux I__6685 (
            .O(N__33647),
            .I(N__33623));
    CascadeMux I__6684 (
            .O(N__33646),
            .I(N__33617));
    CascadeMux I__6683 (
            .O(N__33645),
            .I(N__33614));
    LocalMux I__6682 (
            .O(N__33640),
            .I(N__33608));
    LocalMux I__6681 (
            .O(N__33635),
            .I(N__33608));
    InMux I__6680 (
            .O(N__33634),
            .I(N__33605));
    InMux I__6679 (
            .O(N__33633),
            .I(N__33599));
    InMux I__6678 (
            .O(N__33632),
            .I(N__33596));
    InMux I__6677 (
            .O(N__33629),
            .I(N__33593));
    InMux I__6676 (
            .O(N__33628),
            .I(N__33590));
    CascadeMux I__6675 (
            .O(N__33627),
            .I(N__33587));
    InMux I__6674 (
            .O(N__33626),
            .I(N__33575));
    InMux I__6673 (
            .O(N__33623),
            .I(N__33575));
    InMux I__6672 (
            .O(N__33622),
            .I(N__33575));
    InMux I__6671 (
            .O(N__33621),
            .I(N__33575));
    InMux I__6670 (
            .O(N__33620),
            .I(N__33575));
    InMux I__6669 (
            .O(N__33617),
            .I(N__33567));
    InMux I__6668 (
            .O(N__33614),
            .I(N__33567));
    InMux I__6667 (
            .O(N__33613),
            .I(N__33567));
    Span4Mux_v I__6666 (
            .O(N__33608),
            .I(N__33562));
    LocalMux I__6665 (
            .O(N__33605),
            .I(N__33562));
    CascadeMux I__6664 (
            .O(N__33604),
            .I(N__33552));
    CascadeMux I__6663 (
            .O(N__33603),
            .I(N__33549));
    CascadeMux I__6662 (
            .O(N__33602),
            .I(N__33546));
    LocalMux I__6661 (
            .O(N__33599),
            .I(N__33541));
    LocalMux I__6660 (
            .O(N__33596),
            .I(N__33534));
    LocalMux I__6659 (
            .O(N__33593),
            .I(N__33534));
    LocalMux I__6658 (
            .O(N__33590),
            .I(N__33534));
    InMux I__6657 (
            .O(N__33587),
            .I(N__33529));
    InMux I__6656 (
            .O(N__33586),
            .I(N__33529));
    LocalMux I__6655 (
            .O(N__33575),
            .I(N__33526));
    InMux I__6654 (
            .O(N__33574),
            .I(N__33523));
    LocalMux I__6653 (
            .O(N__33567),
            .I(N__33520));
    Span4Mux_v I__6652 (
            .O(N__33562),
            .I(N__33517));
    InMux I__6651 (
            .O(N__33561),
            .I(N__33510));
    InMux I__6650 (
            .O(N__33560),
            .I(N__33510));
    InMux I__6649 (
            .O(N__33559),
            .I(N__33510));
    InMux I__6648 (
            .O(N__33558),
            .I(N__33501));
    InMux I__6647 (
            .O(N__33557),
            .I(N__33501));
    InMux I__6646 (
            .O(N__33556),
            .I(N__33501));
    InMux I__6645 (
            .O(N__33555),
            .I(N__33501));
    InMux I__6644 (
            .O(N__33552),
            .I(N__33490));
    InMux I__6643 (
            .O(N__33549),
            .I(N__33490));
    InMux I__6642 (
            .O(N__33546),
            .I(N__33490));
    InMux I__6641 (
            .O(N__33545),
            .I(N__33490));
    InMux I__6640 (
            .O(N__33544),
            .I(N__33490));
    Span4Mux_h I__6639 (
            .O(N__33541),
            .I(N__33485));
    Span4Mux_v I__6638 (
            .O(N__33534),
            .I(N__33485));
    LocalMux I__6637 (
            .O(N__33529),
            .I(N__33480));
    Span4Mux_h I__6636 (
            .O(N__33526),
            .I(N__33480));
    LocalMux I__6635 (
            .O(N__33523),
            .I(N__33473));
    Span4Mux_h I__6634 (
            .O(N__33520),
            .I(N__33473));
    Span4Mux_h I__6633 (
            .O(N__33517),
            .I(N__33473));
    LocalMux I__6632 (
            .O(N__33510),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__6631 (
            .O(N__33501),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__6630 (
            .O(N__33490),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__6629 (
            .O(N__33485),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__6628 (
            .O(N__33480),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__6627 (
            .O(N__33473),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    InMux I__6626 (
            .O(N__33460),
            .I(N__33457));
    LocalMux I__6625 (
            .O(N__33457),
            .I(N__33452));
    InMux I__6624 (
            .O(N__33456),
            .I(N__33449));
    InMux I__6623 (
            .O(N__33455),
            .I(N__33446));
    Span4Mux_h I__6622 (
            .O(N__33452),
            .I(N__33438));
    LocalMux I__6621 (
            .O(N__33449),
            .I(N__33433));
    LocalMux I__6620 (
            .O(N__33446),
            .I(N__33433));
    InMux I__6619 (
            .O(N__33445),
            .I(N__33424));
    InMux I__6618 (
            .O(N__33444),
            .I(N__33424));
    InMux I__6617 (
            .O(N__33443),
            .I(N__33424));
    InMux I__6616 (
            .O(N__33442),
            .I(N__33424));
    InMux I__6615 (
            .O(N__33441),
            .I(N__33421));
    Odrv4 I__6614 (
            .O(N__33438),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    Odrv12 I__6613 (
            .O(N__33433),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    LocalMux I__6612 (
            .O(N__33424),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    LocalMux I__6611 (
            .O(N__33421),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    InMux I__6610 (
            .O(N__33412),
            .I(N__33408));
    InMux I__6609 (
            .O(N__33411),
            .I(N__33403));
    LocalMux I__6608 (
            .O(N__33408),
            .I(N__33400));
    InMux I__6607 (
            .O(N__33407),
            .I(N__33397));
    InMux I__6606 (
            .O(N__33406),
            .I(N__33394));
    LocalMux I__6605 (
            .O(N__33403),
            .I(N__33388));
    Span4Mux_h I__6604 (
            .O(N__33400),
            .I(N__33388));
    LocalMux I__6603 (
            .O(N__33397),
            .I(N__33385));
    LocalMux I__6602 (
            .O(N__33394),
            .I(N__33382));
    InMux I__6601 (
            .O(N__33393),
            .I(N__33379));
    Odrv4 I__6600 (
            .O(N__33388),
            .I(measured_delay_hc_12));
    Odrv12 I__6599 (
            .O(N__33385),
            .I(measured_delay_hc_12));
    Odrv4 I__6598 (
            .O(N__33382),
            .I(measured_delay_hc_12));
    LocalMux I__6597 (
            .O(N__33379),
            .I(measured_delay_hc_12));
    InMux I__6596 (
            .O(N__33370),
            .I(N__33366));
    InMux I__6595 (
            .O(N__33369),
            .I(N__33361));
    LocalMux I__6594 (
            .O(N__33366),
            .I(N__33357));
    InMux I__6593 (
            .O(N__33365),
            .I(N__33354));
    InMux I__6592 (
            .O(N__33364),
            .I(N__33351));
    LocalMux I__6591 (
            .O(N__33361),
            .I(N__33348));
    CascadeMux I__6590 (
            .O(N__33360),
            .I(N__33345));
    Span4Mux_v I__6589 (
            .O(N__33357),
            .I(N__33342));
    LocalMux I__6588 (
            .O(N__33354),
            .I(N__33339));
    LocalMux I__6587 (
            .O(N__33351),
            .I(N__33336));
    Span4Mux_v I__6586 (
            .O(N__33348),
            .I(N__33333));
    InMux I__6585 (
            .O(N__33345),
            .I(N__33330));
    Span4Mux_h I__6584 (
            .O(N__33342),
            .I(N__33327));
    Span4Mux_v I__6583 (
            .O(N__33339),
            .I(N__33324));
    Span4Mux_v I__6582 (
            .O(N__33336),
            .I(N__33319));
    Span4Mux_h I__6581 (
            .O(N__33333),
            .I(N__33319));
    LocalMux I__6580 (
            .O(N__33330),
            .I(measured_delay_hc_14));
    Odrv4 I__6579 (
            .O(N__33327),
            .I(measured_delay_hc_14));
    Odrv4 I__6578 (
            .O(N__33324),
            .I(measured_delay_hc_14));
    Odrv4 I__6577 (
            .O(N__33319),
            .I(measured_delay_hc_14));
    InMux I__6576 (
            .O(N__33310),
            .I(N__33303));
    InMux I__6575 (
            .O(N__33309),
            .I(N__33300));
    CascadeMux I__6574 (
            .O(N__33308),
            .I(N__33297));
    InMux I__6573 (
            .O(N__33307),
            .I(N__33294));
    CascadeMux I__6572 (
            .O(N__33306),
            .I(N__33291));
    LocalMux I__6571 (
            .O(N__33303),
            .I(N__33288));
    LocalMux I__6570 (
            .O(N__33300),
            .I(N__33285));
    InMux I__6569 (
            .O(N__33297),
            .I(N__33282));
    LocalMux I__6568 (
            .O(N__33294),
            .I(N__33279));
    InMux I__6567 (
            .O(N__33291),
            .I(N__33276));
    Span4Mux_h I__6566 (
            .O(N__33288),
            .I(N__33273));
    Span4Mux_v I__6565 (
            .O(N__33285),
            .I(N__33266));
    LocalMux I__6564 (
            .O(N__33282),
            .I(N__33266));
    Span4Mux_v I__6563 (
            .O(N__33279),
            .I(N__33266));
    LocalMux I__6562 (
            .O(N__33276),
            .I(measured_delay_hc_16));
    Odrv4 I__6561 (
            .O(N__33273),
            .I(measured_delay_hc_16));
    Odrv4 I__6560 (
            .O(N__33266),
            .I(measured_delay_hc_16));
    InMux I__6559 (
            .O(N__33259),
            .I(N__33255));
    InMux I__6558 (
            .O(N__33258),
            .I(N__33250));
    LocalMux I__6557 (
            .O(N__33255),
            .I(N__33246));
    InMux I__6556 (
            .O(N__33254),
            .I(N__33243));
    InMux I__6555 (
            .O(N__33253),
            .I(N__33240));
    LocalMux I__6554 (
            .O(N__33250),
            .I(N__33237));
    InMux I__6553 (
            .O(N__33249),
            .I(N__33234));
    Span4Mux_v I__6552 (
            .O(N__33246),
            .I(N__33231));
    LocalMux I__6551 (
            .O(N__33243),
            .I(N__33226));
    LocalMux I__6550 (
            .O(N__33240),
            .I(N__33226));
    Span4Mux_v I__6549 (
            .O(N__33237),
            .I(N__33223));
    LocalMux I__6548 (
            .O(N__33234),
            .I(N__33216));
    Span4Mux_h I__6547 (
            .O(N__33231),
            .I(N__33216));
    Span4Mux_v I__6546 (
            .O(N__33226),
            .I(N__33216));
    Odrv4 I__6545 (
            .O(N__33223),
            .I(measured_delay_hc_17));
    Odrv4 I__6544 (
            .O(N__33216),
            .I(measured_delay_hc_17));
    InMux I__6543 (
            .O(N__33211),
            .I(N__33205));
    InMux I__6542 (
            .O(N__33210),
            .I(N__33201));
    CascadeMux I__6541 (
            .O(N__33209),
            .I(N__33198));
    InMux I__6540 (
            .O(N__33208),
            .I(N__33195));
    LocalMux I__6539 (
            .O(N__33205),
            .I(N__33192));
    CascadeMux I__6538 (
            .O(N__33204),
            .I(N__33189));
    LocalMux I__6537 (
            .O(N__33201),
            .I(N__33186));
    InMux I__6536 (
            .O(N__33198),
            .I(N__33183));
    LocalMux I__6535 (
            .O(N__33195),
            .I(N__33178));
    Span4Mux_v I__6534 (
            .O(N__33192),
            .I(N__33178));
    InMux I__6533 (
            .O(N__33189),
            .I(N__33175));
    Span4Mux_h I__6532 (
            .O(N__33186),
            .I(N__33170));
    LocalMux I__6531 (
            .O(N__33183),
            .I(N__33170));
    Odrv4 I__6530 (
            .O(N__33178),
            .I(measured_delay_hc_18));
    LocalMux I__6529 (
            .O(N__33175),
            .I(measured_delay_hc_18));
    Odrv4 I__6528 (
            .O(N__33170),
            .I(measured_delay_hc_18));
    InMux I__6527 (
            .O(N__33163),
            .I(N__33160));
    LocalMux I__6526 (
            .O(N__33160),
            .I(N__33156));
    InMux I__6525 (
            .O(N__33159),
            .I(N__33152));
    Span4Mux_v I__6524 (
            .O(N__33156),
            .I(N__33149));
    InMux I__6523 (
            .O(N__33155),
            .I(N__33146));
    LocalMux I__6522 (
            .O(N__33152),
            .I(N__33143));
    Span4Mux_h I__6521 (
            .O(N__33149),
            .I(N__33140));
    LocalMux I__6520 (
            .O(N__33146),
            .I(N__33135));
    Span4Mux_h I__6519 (
            .O(N__33143),
            .I(N__33135));
    Odrv4 I__6518 (
            .O(N__33140),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    Odrv4 I__6517 (
            .O(N__33135),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    InMux I__6516 (
            .O(N__33130),
            .I(N__33126));
    InMux I__6515 (
            .O(N__33129),
            .I(N__33122));
    LocalMux I__6514 (
            .O(N__33126),
            .I(N__33119));
    InMux I__6513 (
            .O(N__33125),
            .I(N__33116));
    LocalMux I__6512 (
            .O(N__33122),
            .I(N__33112));
    Span4Mux_h I__6511 (
            .O(N__33119),
            .I(N__33109));
    LocalMux I__6510 (
            .O(N__33116),
            .I(N__33106));
    InMux I__6509 (
            .O(N__33115),
            .I(N__33103));
    Span4Mux_v I__6508 (
            .O(N__33112),
            .I(N__33100));
    Span4Mux_v I__6507 (
            .O(N__33109),
            .I(N__33097));
    Span4Mux_v I__6506 (
            .O(N__33106),
            .I(N__33094));
    LocalMux I__6505 (
            .O(N__33103),
            .I(N__33091));
    Odrv4 I__6504 (
            .O(N__33100),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ));
    Odrv4 I__6503 (
            .O(N__33097),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ));
    Odrv4 I__6502 (
            .O(N__33094),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ));
    Odrv4 I__6501 (
            .O(N__33091),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ));
    InMux I__6500 (
            .O(N__33082),
            .I(N__33079));
    LocalMux I__6499 (
            .O(N__33079),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ));
    InMux I__6498 (
            .O(N__33076),
            .I(N__33072));
    InMux I__6497 (
            .O(N__33075),
            .I(N__33069));
    LocalMux I__6496 (
            .O(N__33072),
            .I(N__33066));
    LocalMux I__6495 (
            .O(N__33069),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__6494 (
            .O(N__33066),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__6493 (
            .O(N__33061),
            .I(N__33058));
    LocalMux I__6492 (
            .O(N__33058),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ));
    CascadeMux I__6491 (
            .O(N__33055),
            .I(N__33051));
    InMux I__6490 (
            .O(N__33054),
            .I(N__33048));
    InMux I__6489 (
            .O(N__33051),
            .I(N__33045));
    LocalMux I__6488 (
            .O(N__33048),
            .I(N__33042));
    LocalMux I__6487 (
            .O(N__33045),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv12 I__6486 (
            .O(N__33042),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__6485 (
            .O(N__33037),
            .I(N__33034));
    LocalMux I__6484 (
            .O(N__33034),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ));
    CascadeMux I__6483 (
            .O(N__33031),
            .I(N__33027));
    InMux I__6482 (
            .O(N__33030),
            .I(N__33024));
    InMux I__6481 (
            .O(N__33027),
            .I(N__33021));
    LocalMux I__6480 (
            .O(N__33024),
            .I(N__33018));
    LocalMux I__6479 (
            .O(N__33021),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv12 I__6478 (
            .O(N__33018),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__6477 (
            .O(N__33013),
            .I(N__33010));
    LocalMux I__6476 (
            .O(N__33010),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ));
    InMux I__6475 (
            .O(N__33007),
            .I(N__33003));
    InMux I__6474 (
            .O(N__33006),
            .I(N__33000));
    LocalMux I__6473 (
            .O(N__33003),
            .I(N__32997));
    LocalMux I__6472 (
            .O(N__33000),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv12 I__6471 (
            .O(N__32997),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__6470 (
            .O(N__32992),
            .I(N__32989));
    LocalMux I__6469 (
            .O(N__32989),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ));
    InMux I__6468 (
            .O(N__32986),
            .I(N__32982));
    InMux I__6467 (
            .O(N__32985),
            .I(N__32979));
    LocalMux I__6466 (
            .O(N__32982),
            .I(N__32976));
    LocalMux I__6465 (
            .O(N__32979),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv12 I__6464 (
            .O(N__32976),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__6463 (
            .O(N__32971),
            .I(N__32968));
    LocalMux I__6462 (
            .O(N__32968),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ));
    InMux I__6461 (
            .O(N__32965),
            .I(N__32962));
    LocalMux I__6460 (
            .O(N__32962),
            .I(N__32958));
    InMux I__6459 (
            .O(N__32961),
            .I(N__32955));
    Span4Mux_v I__6458 (
            .O(N__32958),
            .I(N__32952));
    LocalMux I__6457 (
            .O(N__32955),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__6456 (
            .O(N__32952),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__6455 (
            .O(N__32947),
            .I(N__32944));
    LocalMux I__6454 (
            .O(N__32944),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ));
    InMux I__6453 (
            .O(N__32941),
            .I(N__32937));
    InMux I__6452 (
            .O(N__32940),
            .I(N__32934));
    LocalMux I__6451 (
            .O(N__32937),
            .I(N__32931));
    LocalMux I__6450 (
            .O(N__32934),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv12 I__6449 (
            .O(N__32931),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__6448 (
            .O(N__32926),
            .I(N__32920));
    CascadeMux I__6447 (
            .O(N__32925),
            .I(N__32917));
    InMux I__6446 (
            .O(N__32924),
            .I(N__32914));
    CascadeMux I__6445 (
            .O(N__32923),
            .I(N__32910));
    InMux I__6444 (
            .O(N__32920),
            .I(N__32889));
    InMux I__6443 (
            .O(N__32917),
            .I(N__32889));
    LocalMux I__6442 (
            .O(N__32914),
            .I(N__32886));
    InMux I__6441 (
            .O(N__32913),
            .I(N__32869));
    InMux I__6440 (
            .O(N__32910),
            .I(N__32869));
    InMux I__6439 (
            .O(N__32909),
            .I(N__32869));
    InMux I__6438 (
            .O(N__32908),
            .I(N__32869));
    InMux I__6437 (
            .O(N__32907),
            .I(N__32869));
    InMux I__6436 (
            .O(N__32906),
            .I(N__32869));
    InMux I__6435 (
            .O(N__32905),
            .I(N__32869));
    InMux I__6434 (
            .O(N__32904),
            .I(N__32869));
    InMux I__6433 (
            .O(N__32903),
            .I(N__32858));
    InMux I__6432 (
            .O(N__32902),
            .I(N__32858));
    InMux I__6431 (
            .O(N__32901),
            .I(N__32858));
    InMux I__6430 (
            .O(N__32900),
            .I(N__32858));
    InMux I__6429 (
            .O(N__32899),
            .I(N__32858));
    InMux I__6428 (
            .O(N__32898),
            .I(N__32853));
    InMux I__6427 (
            .O(N__32897),
            .I(N__32853));
    InMux I__6426 (
            .O(N__32896),
            .I(N__32848));
    InMux I__6425 (
            .O(N__32895),
            .I(N__32843));
    InMux I__6424 (
            .O(N__32894),
            .I(N__32843));
    LocalMux I__6423 (
            .O(N__32889),
            .I(N__32834));
    Span4Mux_v I__6422 (
            .O(N__32886),
            .I(N__32834));
    LocalMux I__6421 (
            .O(N__32869),
            .I(N__32834));
    LocalMux I__6420 (
            .O(N__32858),
            .I(N__32834));
    LocalMux I__6419 (
            .O(N__32853),
            .I(N__32831));
    InMux I__6418 (
            .O(N__32852),
            .I(N__32828));
    InMux I__6417 (
            .O(N__32851),
            .I(N__32825));
    LocalMux I__6416 (
            .O(N__32848),
            .I(N__32822));
    LocalMux I__6415 (
            .O(N__32843),
            .I(N__32819));
    Span4Mux_v I__6414 (
            .O(N__32834),
            .I(N__32814));
    Span4Mux_v I__6413 (
            .O(N__32831),
            .I(N__32814));
    LocalMux I__6412 (
            .O(N__32828),
            .I(N__32811));
    LocalMux I__6411 (
            .O(N__32825),
            .I(N__32805));
    Span12Mux_v I__6410 (
            .O(N__32822),
            .I(N__32805));
    Span4Mux_h I__6409 (
            .O(N__32819),
            .I(N__32800));
    Span4Mux_h I__6408 (
            .O(N__32814),
            .I(N__32800));
    Span4Mux_v I__6407 (
            .O(N__32811),
            .I(N__32797));
    InMux I__6406 (
            .O(N__32810),
            .I(N__32794));
    Odrv12 I__6405 (
            .O(N__32805),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__6404 (
            .O(N__32800),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__6403 (
            .O(N__32797),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__6402 (
            .O(N__32794),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__6401 (
            .O(N__32785),
            .I(N__32782));
    LocalMux I__6400 (
            .O(N__32782),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ));
    CascadeMux I__6399 (
            .O(N__32779),
            .I(N__32767));
    CascadeMux I__6398 (
            .O(N__32778),
            .I(N__32764));
    CascadeMux I__6397 (
            .O(N__32777),
            .I(N__32761));
    CascadeMux I__6396 (
            .O(N__32776),
            .I(N__32754));
    CascadeMux I__6395 (
            .O(N__32775),
            .I(N__32751));
    CascadeMux I__6394 (
            .O(N__32774),
            .I(N__32748));
    CascadeMux I__6393 (
            .O(N__32773),
            .I(N__32745));
    CascadeMux I__6392 (
            .O(N__32772),
            .I(N__32741));
    CascadeMux I__6391 (
            .O(N__32771),
            .I(N__32738));
    CascadeMux I__6390 (
            .O(N__32770),
            .I(N__32734));
    InMux I__6389 (
            .O(N__32767),
            .I(N__32718));
    InMux I__6388 (
            .O(N__32764),
            .I(N__32718));
    InMux I__6387 (
            .O(N__32761),
            .I(N__32718));
    InMux I__6386 (
            .O(N__32760),
            .I(N__32718));
    InMux I__6385 (
            .O(N__32759),
            .I(N__32718));
    InMux I__6384 (
            .O(N__32758),
            .I(N__32718));
    InMux I__6383 (
            .O(N__32757),
            .I(N__32715));
    InMux I__6382 (
            .O(N__32754),
            .I(N__32712));
    InMux I__6381 (
            .O(N__32751),
            .I(N__32703));
    InMux I__6380 (
            .O(N__32748),
            .I(N__32703));
    InMux I__6379 (
            .O(N__32745),
            .I(N__32703));
    InMux I__6378 (
            .O(N__32744),
            .I(N__32703));
    InMux I__6377 (
            .O(N__32741),
            .I(N__32694));
    InMux I__6376 (
            .O(N__32738),
            .I(N__32694));
    InMux I__6375 (
            .O(N__32737),
            .I(N__32694));
    InMux I__6374 (
            .O(N__32734),
            .I(N__32694));
    CascadeMux I__6373 (
            .O(N__32733),
            .I(N__32691));
    CascadeMux I__6372 (
            .O(N__32732),
            .I(N__32687));
    InMux I__6371 (
            .O(N__32731),
            .I(N__32681));
    LocalMux I__6370 (
            .O(N__32718),
            .I(N__32678));
    LocalMux I__6369 (
            .O(N__32715),
            .I(N__32669));
    LocalMux I__6368 (
            .O(N__32712),
            .I(N__32669));
    LocalMux I__6367 (
            .O(N__32703),
            .I(N__32669));
    LocalMux I__6366 (
            .O(N__32694),
            .I(N__32669));
    InMux I__6365 (
            .O(N__32691),
            .I(N__32666));
    InMux I__6364 (
            .O(N__32690),
            .I(N__32661));
    InMux I__6363 (
            .O(N__32687),
            .I(N__32661));
    InMux I__6362 (
            .O(N__32686),
            .I(N__32656));
    InMux I__6361 (
            .O(N__32685),
            .I(N__32656));
    CascadeMux I__6360 (
            .O(N__32684),
            .I(N__32653));
    LocalMux I__6359 (
            .O(N__32681),
            .I(N__32650));
    Span4Mux_v I__6358 (
            .O(N__32678),
            .I(N__32645));
    Span4Mux_v I__6357 (
            .O(N__32669),
            .I(N__32645));
    LocalMux I__6356 (
            .O(N__32666),
            .I(N__32642));
    LocalMux I__6355 (
            .O(N__32661),
            .I(N__32639));
    LocalMux I__6354 (
            .O(N__32656),
            .I(N__32636));
    InMux I__6353 (
            .O(N__32653),
            .I(N__32633));
    Span4Mux_v I__6352 (
            .O(N__32650),
            .I(N__32630));
    Span4Mux_v I__6351 (
            .O(N__32645),
            .I(N__32627));
    Span4Mux_h I__6350 (
            .O(N__32642),
            .I(N__32623));
    Span4Mux_v I__6349 (
            .O(N__32639),
            .I(N__32620));
    Span12Mux_v I__6348 (
            .O(N__32636),
            .I(N__32617));
    LocalMux I__6347 (
            .O(N__32633),
            .I(N__32610));
    Span4Mux_v I__6346 (
            .O(N__32630),
            .I(N__32610));
    Span4Mux_v I__6345 (
            .O(N__32627),
            .I(N__32610));
    InMux I__6344 (
            .O(N__32626),
            .I(N__32607));
    Odrv4 I__6343 (
            .O(N__32623),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__6342 (
            .O(N__32620),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv12 I__6341 (
            .O(N__32617),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__6340 (
            .O(N__32610),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__6339 (
            .O(N__32607),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__6338 (
            .O(N__32596),
            .I(N__32591));
    CascadeMux I__6337 (
            .O(N__32595),
            .I(N__32587));
    CascadeMux I__6336 (
            .O(N__32594),
            .I(N__32577));
    InMux I__6335 (
            .O(N__32591),
            .I(N__32565));
    InMux I__6334 (
            .O(N__32590),
            .I(N__32548));
    InMux I__6333 (
            .O(N__32587),
            .I(N__32548));
    InMux I__6332 (
            .O(N__32586),
            .I(N__32548));
    InMux I__6331 (
            .O(N__32585),
            .I(N__32548));
    InMux I__6330 (
            .O(N__32584),
            .I(N__32548));
    InMux I__6329 (
            .O(N__32583),
            .I(N__32548));
    InMux I__6328 (
            .O(N__32582),
            .I(N__32548));
    InMux I__6327 (
            .O(N__32581),
            .I(N__32548));
    InMux I__6326 (
            .O(N__32580),
            .I(N__32545));
    InMux I__6325 (
            .O(N__32577),
            .I(N__32530));
    InMux I__6324 (
            .O(N__32576),
            .I(N__32530));
    InMux I__6323 (
            .O(N__32575),
            .I(N__32530));
    InMux I__6322 (
            .O(N__32574),
            .I(N__32530));
    InMux I__6321 (
            .O(N__32573),
            .I(N__32530));
    InMux I__6320 (
            .O(N__32572),
            .I(N__32530));
    InMux I__6319 (
            .O(N__32571),
            .I(N__32530));
    CascadeMux I__6318 (
            .O(N__32570),
            .I(N__32527));
    InMux I__6317 (
            .O(N__32569),
            .I(N__32521));
    InMux I__6316 (
            .O(N__32568),
            .I(N__32521));
    LocalMux I__6315 (
            .O(N__32565),
            .I(N__32518));
    LocalMux I__6314 (
            .O(N__32548),
            .I(N__32515));
    LocalMux I__6313 (
            .O(N__32545),
            .I(N__32510));
    LocalMux I__6312 (
            .O(N__32530),
            .I(N__32510));
    InMux I__6311 (
            .O(N__32527),
            .I(N__32506));
    InMux I__6310 (
            .O(N__32526),
            .I(N__32503));
    LocalMux I__6309 (
            .O(N__32521),
            .I(N__32500));
    Span4Mux_v I__6308 (
            .O(N__32518),
            .I(N__32492));
    Span4Mux_v I__6307 (
            .O(N__32515),
            .I(N__32492));
    Span4Mux_v I__6306 (
            .O(N__32510),
            .I(N__32492));
    InMux I__6305 (
            .O(N__32509),
            .I(N__32489));
    LocalMux I__6304 (
            .O(N__32506),
            .I(N__32484));
    LocalMux I__6303 (
            .O(N__32503),
            .I(N__32484));
    Span4Mux_h I__6302 (
            .O(N__32500),
            .I(N__32481));
    InMux I__6301 (
            .O(N__32499),
            .I(N__32478));
    Span4Mux_h I__6300 (
            .O(N__32492),
            .I(N__32473));
    LocalMux I__6299 (
            .O(N__32489),
            .I(N__32473));
    Span4Mux_v I__6298 (
            .O(N__32484),
            .I(N__32469));
    Span4Mux_v I__6297 (
            .O(N__32481),
            .I(N__32466));
    LocalMux I__6296 (
            .O(N__32478),
            .I(N__32461));
    Span4Mux_v I__6295 (
            .O(N__32473),
            .I(N__32461));
    InMux I__6294 (
            .O(N__32472),
            .I(N__32458));
    Span4Mux_h I__6293 (
            .O(N__32469),
            .I(N__32453));
    Span4Mux_v I__6292 (
            .O(N__32466),
            .I(N__32453));
    Span4Mux_v I__6291 (
            .O(N__32461),
            .I(N__32450));
    LocalMux I__6290 (
            .O(N__32458),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__6289 (
            .O(N__32453),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__6288 (
            .O(N__32450),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    InMux I__6287 (
            .O(N__32443),
            .I(N__32439));
    InMux I__6286 (
            .O(N__32442),
            .I(N__32436));
    LocalMux I__6285 (
            .O(N__32439),
            .I(N__32433));
    LocalMux I__6284 (
            .O(N__32436),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__6283 (
            .O(N__32433),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__6282 (
            .O(N__32428),
            .I(N__32425));
    LocalMux I__6281 (
            .O(N__32425),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ));
    InMux I__6280 (
            .O(N__32422),
            .I(N__32418));
    InMux I__6279 (
            .O(N__32421),
            .I(N__32415));
    LocalMux I__6278 (
            .O(N__32418),
            .I(N__32412));
    LocalMux I__6277 (
            .O(N__32415),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__6276 (
            .O(N__32412),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__6275 (
            .O(N__32407),
            .I(N__32403));
    InMux I__6274 (
            .O(N__32406),
            .I(N__32398));
    LocalMux I__6273 (
            .O(N__32403),
            .I(N__32395));
    InMux I__6272 (
            .O(N__32402),
            .I(N__32392));
    InMux I__6271 (
            .O(N__32401),
            .I(N__32389));
    LocalMux I__6270 (
            .O(N__32398),
            .I(N__32386));
    Span4Mux_v I__6269 (
            .O(N__32395),
            .I(N__32379));
    LocalMux I__6268 (
            .O(N__32392),
            .I(N__32379));
    LocalMux I__6267 (
            .O(N__32389),
            .I(N__32379));
    Span4Mux_h I__6266 (
            .O(N__32386),
            .I(N__32376));
    Span4Mux_h I__6265 (
            .O(N__32379),
            .I(N__32373));
    Odrv4 I__6264 (
            .O(N__32376),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    Odrv4 I__6263 (
            .O(N__32373),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    InMux I__6262 (
            .O(N__32368),
            .I(N__32364));
    InMux I__6261 (
            .O(N__32367),
            .I(N__32361));
    LocalMux I__6260 (
            .O(N__32364),
            .I(N__32357));
    LocalMux I__6259 (
            .O(N__32361),
            .I(N__32354));
    InMux I__6258 (
            .O(N__32360),
            .I(N__32351));
    Span4Mux_v I__6257 (
            .O(N__32357),
            .I(N__32345));
    Span12Mux_h I__6256 (
            .O(N__32354),
            .I(N__32342));
    LocalMux I__6255 (
            .O(N__32351),
            .I(N__32339));
    InMux I__6254 (
            .O(N__32350),
            .I(N__32336));
    InMux I__6253 (
            .O(N__32349),
            .I(N__32331));
    InMux I__6252 (
            .O(N__32348),
            .I(N__32331));
    Odrv4 I__6251 (
            .O(N__32345),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__6250 (
            .O(N__32342),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__6249 (
            .O(N__32339),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__6248 (
            .O(N__32336),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__6247 (
            .O(N__32331),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__6246 (
            .O(N__32320),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    CascadeMux I__6245 (
            .O(N__32317),
            .I(N__32312));
    InMux I__6244 (
            .O(N__32316),
            .I(N__32309));
    InMux I__6243 (
            .O(N__32315),
            .I(N__32306));
    InMux I__6242 (
            .O(N__32312),
            .I(N__32303));
    LocalMux I__6241 (
            .O(N__32309),
            .I(N__32300));
    LocalMux I__6240 (
            .O(N__32306),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__6239 (
            .O(N__32303),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__6238 (
            .O(N__32300),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__6237 (
            .O(N__32293),
            .I(N__32290));
    LocalMux I__6236 (
            .O(N__32290),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ));
    InMux I__6235 (
            .O(N__32287),
            .I(N__32283));
    InMux I__6234 (
            .O(N__32286),
            .I(N__32280));
    LocalMux I__6233 (
            .O(N__32283),
            .I(N__32277));
    LocalMux I__6232 (
            .O(N__32280),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__6231 (
            .O(N__32277),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__6230 (
            .O(N__32272),
            .I(N__32269));
    LocalMux I__6229 (
            .O(N__32269),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ));
    InMux I__6228 (
            .O(N__32266),
            .I(N__32262));
    InMux I__6227 (
            .O(N__32265),
            .I(N__32259));
    LocalMux I__6226 (
            .O(N__32262),
            .I(N__32256));
    LocalMux I__6225 (
            .O(N__32259),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__6224 (
            .O(N__32256),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__6223 (
            .O(N__32251),
            .I(N__32248));
    LocalMux I__6222 (
            .O(N__32248),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ));
    InMux I__6221 (
            .O(N__32245),
            .I(N__32241));
    InMux I__6220 (
            .O(N__32244),
            .I(N__32238));
    LocalMux I__6219 (
            .O(N__32241),
            .I(N__32235));
    LocalMux I__6218 (
            .O(N__32238),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__6217 (
            .O(N__32235),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__6216 (
            .O(N__32230),
            .I(N__32227));
    LocalMux I__6215 (
            .O(N__32227),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ));
    InMux I__6214 (
            .O(N__32224),
            .I(N__32220));
    InMux I__6213 (
            .O(N__32223),
            .I(N__32217));
    LocalMux I__6212 (
            .O(N__32220),
            .I(N__32214));
    LocalMux I__6211 (
            .O(N__32217),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__6210 (
            .O(N__32214),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__6209 (
            .O(N__32209),
            .I(N__32206));
    LocalMux I__6208 (
            .O(N__32206),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ));
    InMux I__6207 (
            .O(N__32203),
            .I(N__32199));
    InMux I__6206 (
            .O(N__32202),
            .I(N__32196));
    LocalMux I__6205 (
            .O(N__32199),
            .I(N__32193));
    LocalMux I__6204 (
            .O(N__32196),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__6203 (
            .O(N__32193),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__6202 (
            .O(N__32188),
            .I(N__32185));
    LocalMux I__6201 (
            .O(N__32185),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ));
    InMux I__6200 (
            .O(N__32182),
            .I(N__32178));
    InMux I__6199 (
            .O(N__32181),
            .I(N__32175));
    LocalMux I__6198 (
            .O(N__32178),
            .I(N__32172));
    LocalMux I__6197 (
            .O(N__32175),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__6196 (
            .O(N__32172),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    CascadeMux I__6195 (
            .O(N__32167),
            .I(N__32164));
    InMux I__6194 (
            .O(N__32164),
            .I(N__32161));
    LocalMux I__6193 (
            .O(N__32161),
            .I(N__32158));
    Span4Mux_h I__6192 (
            .O(N__32158),
            .I(N__32155));
    Odrv4 I__6191 (
            .O(N__32155),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__6190 (
            .O(N__32152),
            .I(N__32149));
    LocalMux I__6189 (
            .O(N__32149),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__6188 (
            .O(N__32146),
            .I(N__32142));
    CascadeMux I__6187 (
            .O(N__32145),
            .I(N__32139));
    LocalMux I__6186 (
            .O(N__32142),
            .I(N__32136));
    InMux I__6185 (
            .O(N__32139),
            .I(N__32133));
    Span4Mux_h I__6184 (
            .O(N__32136),
            .I(N__32130));
    LocalMux I__6183 (
            .O(N__32133),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__6182 (
            .O(N__32130),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__6181 (
            .O(N__32125),
            .I(N__32122));
    LocalMux I__6180 (
            .O(N__32122),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    InMux I__6179 (
            .O(N__32119),
            .I(N__32116));
    LocalMux I__6178 (
            .O(N__32116),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    CascadeMux I__6177 (
            .O(N__32113),
            .I(N__32110));
    InMux I__6176 (
            .O(N__32110),
            .I(N__32107));
    LocalMux I__6175 (
            .O(N__32107),
            .I(N__32104));
    Odrv12 I__6174 (
            .O(N__32104),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__6173 (
            .O(N__32101),
            .I(N__32098));
    LocalMux I__6172 (
            .O(N__32098),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    InMux I__6171 (
            .O(N__32095),
            .I(N__32092));
    LocalMux I__6170 (
            .O(N__32092),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__6169 (
            .O(N__32089),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__6168 (
            .O(N__32086),
            .I(N__32083));
    InMux I__6167 (
            .O(N__32083),
            .I(N__32080));
    LocalMux I__6166 (
            .O(N__32080),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__6165 (
            .O(N__32077),
            .I(N__32074));
    InMux I__6164 (
            .O(N__32074),
            .I(N__32071));
    LocalMux I__6163 (
            .O(N__32071),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__6162 (
            .O(N__32068),
            .I(N__32065));
    InMux I__6161 (
            .O(N__32065),
            .I(N__32062));
    LocalMux I__6160 (
            .O(N__32062),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__6159 (
            .O(N__32059),
            .I(N__32056));
    LocalMux I__6158 (
            .O(N__32056),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__6157 (
            .O(N__32053),
            .I(N__32050));
    InMux I__6156 (
            .O(N__32050),
            .I(N__32047));
    LocalMux I__6155 (
            .O(N__32047),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    InMux I__6154 (
            .O(N__32044),
            .I(N__32040));
    InMux I__6153 (
            .O(N__32043),
            .I(N__32037));
    LocalMux I__6152 (
            .O(N__32040),
            .I(N__32034));
    LocalMux I__6151 (
            .O(N__32037),
            .I(N__32031));
    Odrv12 I__6150 (
            .O(N__32034),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__6149 (
            .O(N__32031),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__6148 (
            .O(N__32026),
            .I(N__32023));
    LocalMux I__6147 (
            .O(N__32023),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__6146 (
            .O(N__32020),
            .I(N__32017));
    InMux I__6145 (
            .O(N__32017),
            .I(N__32014));
    LocalMux I__6144 (
            .O(N__32014),
            .I(N__32011));
    Odrv4 I__6143 (
            .O(N__32011),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__6142 (
            .O(N__32008),
            .I(N__32004));
    InMux I__6141 (
            .O(N__32007),
            .I(N__32001));
    LocalMux I__6140 (
            .O(N__32004),
            .I(N__31998));
    LocalMux I__6139 (
            .O(N__32001),
            .I(N__31995));
    Odrv12 I__6138 (
            .O(N__31998),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__6137 (
            .O(N__31995),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__6136 (
            .O(N__31990),
            .I(N__31987));
    LocalMux I__6135 (
            .O(N__31987),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__6134 (
            .O(N__31984),
            .I(N__31981));
    LocalMux I__6133 (
            .O(N__31981),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__6132 (
            .O(N__31978),
            .I(N__31975));
    LocalMux I__6131 (
            .O(N__31975),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__6130 (
            .O(N__31972),
            .I(N__31969));
    LocalMux I__6129 (
            .O(N__31969),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__6128 (
            .O(N__31966),
            .I(N__31963));
    LocalMux I__6127 (
            .O(N__31963),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__6126 (
            .O(N__31960),
            .I(N__31957));
    InMux I__6125 (
            .O(N__31957),
            .I(N__31954));
    LocalMux I__6124 (
            .O(N__31954),
            .I(N__31951));
    Odrv4 I__6123 (
            .O(N__31951),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__6122 (
            .O(N__31948),
            .I(N__31945));
    LocalMux I__6121 (
            .O(N__31945),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__6120 (
            .O(N__31942),
            .I(N__31939));
    InMux I__6119 (
            .O(N__31939),
            .I(N__31936));
    LocalMux I__6118 (
            .O(N__31936),
            .I(N__31933));
    Span4Mux_v I__6117 (
            .O(N__31933),
            .I(N__31930));
    Odrv4 I__6116 (
            .O(N__31930),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__6115 (
            .O(N__31927),
            .I(N__31924));
    LocalMux I__6114 (
            .O(N__31924),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__6113 (
            .O(N__31921),
            .I(N__31918));
    InMux I__6112 (
            .O(N__31918),
            .I(N__31915));
    LocalMux I__6111 (
            .O(N__31915),
            .I(N__31912));
    Odrv4 I__6110 (
            .O(N__31912),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    InMux I__6109 (
            .O(N__31909),
            .I(N__31906));
    LocalMux I__6108 (
            .O(N__31906),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__6107 (
            .O(N__31903),
            .I(N__31900));
    InMux I__6106 (
            .O(N__31900),
            .I(N__31897));
    LocalMux I__6105 (
            .O(N__31897),
            .I(N__31894));
    Odrv12 I__6104 (
            .O(N__31894),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    InMux I__6103 (
            .O(N__31891),
            .I(N__31888));
    LocalMux I__6102 (
            .O(N__31888),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__6101 (
            .O(N__31885),
            .I(N__31882));
    LocalMux I__6100 (
            .O(N__31882),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__6099 (
            .O(N__31879),
            .I(N__31876));
    InMux I__6098 (
            .O(N__31876),
            .I(N__31873));
    LocalMux I__6097 (
            .O(N__31873),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__6096 (
            .O(N__31870),
            .I(N__31867));
    LocalMux I__6095 (
            .O(N__31867),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__6094 (
            .O(N__31864),
            .I(N__31861));
    InMux I__6093 (
            .O(N__31861),
            .I(N__31858));
    LocalMux I__6092 (
            .O(N__31858),
            .I(N__31855));
    Odrv4 I__6091 (
            .O(N__31855),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    InMux I__6090 (
            .O(N__31852),
            .I(N__31849));
    LocalMux I__6089 (
            .O(N__31849),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__6088 (
            .O(N__31846),
            .I(N__31841));
    InMux I__6087 (
            .O(N__31845),
            .I(N__31838));
    InMux I__6086 (
            .O(N__31844),
            .I(N__31835));
    LocalMux I__6085 (
            .O(N__31841),
            .I(N__31832));
    LocalMux I__6084 (
            .O(N__31838),
            .I(N__31826));
    LocalMux I__6083 (
            .O(N__31835),
            .I(N__31826));
    Span4Mux_h I__6082 (
            .O(N__31832),
            .I(N__31823));
    InMux I__6081 (
            .O(N__31831),
            .I(N__31820));
    Span4Mux_v I__6080 (
            .O(N__31826),
            .I(N__31817));
    Span4Mux_v I__6079 (
            .O(N__31823),
            .I(N__31814));
    LocalMux I__6078 (
            .O(N__31820),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    Odrv4 I__6077 (
            .O(N__31817),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    Odrv4 I__6076 (
            .O(N__31814),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    InMux I__6075 (
            .O(N__31807),
            .I(N__31804));
    LocalMux I__6074 (
            .O(N__31804),
            .I(N__31801));
    Span4Mux_h I__6073 (
            .O(N__31801),
            .I(N__31798));
    Span4Mux_v I__6072 (
            .O(N__31798),
            .I(N__31795));
    Odrv4 I__6071 (
            .O(N__31795),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ));
    InMux I__6070 (
            .O(N__31792),
            .I(N__31788));
    InMux I__6069 (
            .O(N__31791),
            .I(N__31785));
    LocalMux I__6068 (
            .O(N__31788),
            .I(N__31781));
    LocalMux I__6067 (
            .O(N__31785),
            .I(N__31778));
    InMux I__6066 (
            .O(N__31784),
            .I(N__31775));
    Span4Mux_v I__6065 (
            .O(N__31781),
            .I(N__31772));
    Span4Mux_v I__6064 (
            .O(N__31778),
            .I(N__31769));
    LocalMux I__6063 (
            .O(N__31775),
            .I(\current_shift_inst.start_timer_phaseZ0 ));
    Odrv4 I__6062 (
            .O(N__31772),
            .I(\current_shift_inst.start_timer_phaseZ0 ));
    Odrv4 I__6061 (
            .O(N__31769),
            .I(\current_shift_inst.start_timer_phaseZ0 ));
    InMux I__6060 (
            .O(N__31762),
            .I(N__31757));
    InMux I__6059 (
            .O(N__31761),
            .I(N__31754));
    InMux I__6058 (
            .O(N__31760),
            .I(N__31751));
    LocalMux I__6057 (
            .O(N__31757),
            .I(N__31747));
    LocalMux I__6056 (
            .O(N__31754),
            .I(N__31744));
    LocalMux I__6055 (
            .O(N__31751),
            .I(N__31741));
    InMux I__6054 (
            .O(N__31750),
            .I(N__31738));
    Span12Mux_h I__6053 (
            .O(N__31747),
            .I(N__31735));
    Span12Mux_v I__6052 (
            .O(N__31744),
            .I(N__31732));
    Span4Mux_h I__6051 (
            .O(N__31741),
            .I(N__31729));
    LocalMux I__6050 (
            .O(N__31738),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    Odrv12 I__6049 (
            .O(N__31735),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    Odrv12 I__6048 (
            .O(N__31732),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    Odrv4 I__6047 (
            .O(N__31729),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    CascadeMux I__6046 (
            .O(N__31720),
            .I(N__31717));
    InMux I__6045 (
            .O(N__31717),
            .I(N__31714));
    LocalMux I__6044 (
            .O(N__31714),
            .I(N__31711));
    Span4Mux_v I__6043 (
            .O(N__31711),
            .I(N__31708));
    Span4Mux_h I__6042 (
            .O(N__31708),
            .I(N__31705));
    Span4Mux_v I__6041 (
            .O(N__31705),
            .I(N__31702));
    Odrv4 I__6040 (
            .O(N__31702),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ));
    CascadeMux I__6039 (
            .O(N__31699),
            .I(N__31696));
    InMux I__6038 (
            .O(N__31696),
            .I(N__31693));
    LocalMux I__6037 (
            .O(N__31693),
            .I(N__31690));
    Span4Mux_v I__6036 (
            .O(N__31690),
            .I(N__31687));
    Span4Mux_v I__6035 (
            .O(N__31687),
            .I(N__31684));
    Odrv4 I__6034 (
            .O(N__31684),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ));
    InMux I__6033 (
            .O(N__31681),
            .I(N__31678));
    LocalMux I__6032 (
            .O(N__31678),
            .I(N__31675));
    Span4Mux_h I__6031 (
            .O(N__31675),
            .I(N__31672));
    Span4Mux_v I__6030 (
            .O(N__31672),
            .I(N__31669));
    Odrv4 I__6029 (
            .O(N__31669),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ));
    InMux I__6028 (
            .O(N__31666),
            .I(N__31663));
    LocalMux I__6027 (
            .O(N__31663),
            .I(N__31660));
    Span4Mux_h I__6026 (
            .O(N__31660),
            .I(N__31657));
    Span4Mux_v I__6025 (
            .O(N__31657),
            .I(N__31654));
    Odrv4 I__6024 (
            .O(N__31654),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ));
    InMux I__6023 (
            .O(N__31651),
            .I(N__31648));
    LocalMux I__6022 (
            .O(N__31648),
            .I(N__31645));
    Span4Mux_v I__6021 (
            .O(N__31645),
            .I(N__31642));
    Span4Mux_h I__6020 (
            .O(N__31642),
            .I(N__31639));
    Odrv4 I__6019 (
            .O(N__31639),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ));
    InMux I__6018 (
            .O(N__31636),
            .I(N__31633));
    LocalMux I__6017 (
            .O(N__31633),
            .I(N__31630));
    Span4Mux_h I__6016 (
            .O(N__31630),
            .I(N__31627));
    Span4Mux_v I__6015 (
            .O(N__31627),
            .I(N__31624));
    Odrv4 I__6014 (
            .O(N__31624),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ));
    InMux I__6013 (
            .O(N__31621),
            .I(N__31618));
    LocalMux I__6012 (
            .O(N__31618),
            .I(N__31615));
    Span4Mux_v I__6011 (
            .O(N__31615),
            .I(N__31612));
    Odrv4 I__6010 (
            .O(N__31612),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ));
    CascadeMux I__6009 (
            .O(N__31609),
            .I(N__31606));
    InMux I__6008 (
            .O(N__31606),
            .I(N__31603));
    LocalMux I__6007 (
            .O(N__31603),
            .I(N__31600));
    Span4Mux_v I__6006 (
            .O(N__31600),
            .I(N__31597));
    Span4Mux_h I__6005 (
            .O(N__31597),
            .I(N__31594));
    Span4Mux_v I__6004 (
            .O(N__31594),
            .I(N__31591));
    Odrv4 I__6003 (
            .O(N__31591),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ));
    InMux I__6002 (
            .O(N__31588),
            .I(N__31585));
    LocalMux I__6001 (
            .O(N__31585),
            .I(N__31582));
    Span4Mux_v I__6000 (
            .O(N__31582),
            .I(N__31579));
    Span4Mux_v I__5999 (
            .O(N__31579),
            .I(N__31576));
    Odrv4 I__5998 (
            .O(N__31576),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ));
    CascadeMux I__5997 (
            .O(N__31573),
            .I(N__31570));
    InMux I__5996 (
            .O(N__31570),
            .I(N__31567));
    LocalMux I__5995 (
            .O(N__31567),
            .I(N__31564));
    Span4Mux_v I__5994 (
            .O(N__31564),
            .I(N__31561));
    Span4Mux_v I__5993 (
            .O(N__31561),
            .I(N__31558));
    Odrv4 I__5992 (
            .O(N__31558),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ));
    InMux I__5991 (
            .O(N__31555),
            .I(N__31552));
    LocalMux I__5990 (
            .O(N__31552),
            .I(N__31549));
    Span4Mux_h I__5989 (
            .O(N__31549),
            .I(N__31546));
    Span4Mux_v I__5988 (
            .O(N__31546),
            .I(N__31543));
    Odrv4 I__5987 (
            .O(N__31543),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ));
    InMux I__5986 (
            .O(N__31540),
            .I(N__31537));
    LocalMux I__5985 (
            .O(N__31537),
            .I(N__31534));
    Span4Mux_h I__5984 (
            .O(N__31534),
            .I(N__31531));
    Span4Mux_v I__5983 (
            .O(N__31531),
            .I(N__31528));
    Odrv4 I__5982 (
            .O(N__31528),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ));
    InMux I__5981 (
            .O(N__31525),
            .I(N__31522));
    LocalMux I__5980 (
            .O(N__31522),
            .I(N__31519));
    Span4Mux_h I__5979 (
            .O(N__31519),
            .I(N__31516));
    Span4Mux_v I__5978 (
            .O(N__31516),
            .I(N__31513));
    Odrv4 I__5977 (
            .O(N__31513),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ));
    InMux I__5976 (
            .O(N__31510),
            .I(N__31507));
    LocalMux I__5975 (
            .O(N__31507),
            .I(N__31504));
    Span4Mux_h I__5974 (
            .O(N__31504),
            .I(N__31501));
    Span4Mux_v I__5973 (
            .O(N__31501),
            .I(N__31498));
    Odrv4 I__5972 (
            .O(N__31498),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ));
    InMux I__5971 (
            .O(N__31495),
            .I(N__31492));
    LocalMux I__5970 (
            .O(N__31492),
            .I(N__31489));
    Span12Mux_h I__5969 (
            .O(N__31489),
            .I(N__31486));
    Odrv12 I__5968 (
            .O(N__31486),
            .I(\current_shift_inst.un38_control_input_0_axb_31 ));
    CascadeMux I__5967 (
            .O(N__31483),
            .I(N__31480));
    InMux I__5966 (
            .O(N__31480),
            .I(N__31477));
    LocalMux I__5965 (
            .O(N__31477),
            .I(N__31474));
    Span4Mux_h I__5964 (
            .O(N__31474),
            .I(N__31471));
    Span4Mux_v I__5963 (
            .O(N__31471),
            .I(N__31468));
    Odrv4 I__5962 (
            .O(N__31468),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ));
    CEMux I__5961 (
            .O(N__31465),
            .I(N__31461));
    CEMux I__5960 (
            .O(N__31464),
            .I(N__31458));
    LocalMux I__5959 (
            .O(N__31461),
            .I(N__31455));
    LocalMux I__5958 (
            .O(N__31458),
            .I(N__31451));
    Span4Mux_v I__5957 (
            .O(N__31455),
            .I(N__31448));
    CEMux I__5956 (
            .O(N__31454),
            .I(N__31445));
    Span4Mux_v I__5955 (
            .O(N__31451),
            .I(N__31441));
    Span4Mux_v I__5954 (
            .O(N__31448),
            .I(N__31436));
    LocalMux I__5953 (
            .O(N__31445),
            .I(N__31436));
    CEMux I__5952 (
            .O(N__31444),
            .I(N__31433));
    Span4Mux_h I__5951 (
            .O(N__31441),
            .I(N__31424));
    Span4Mux_v I__5950 (
            .O(N__31436),
            .I(N__31424));
    LocalMux I__5949 (
            .O(N__31433),
            .I(N__31424));
    CEMux I__5948 (
            .O(N__31432),
            .I(N__31421));
    IoInMux I__5947 (
            .O(N__31431),
            .I(N__31418));
    Span4Mux_v I__5946 (
            .O(N__31424),
            .I(N__31413));
    LocalMux I__5945 (
            .O(N__31421),
            .I(N__31413));
    LocalMux I__5944 (
            .O(N__31418),
            .I(N__31409));
    Span4Mux_v I__5943 (
            .O(N__31413),
            .I(N__31406));
    CEMux I__5942 (
            .O(N__31412),
            .I(N__31403));
    Span4Mux_s1_v I__5941 (
            .O(N__31409),
            .I(N__31400));
    Sp12to4 I__5940 (
            .O(N__31406),
            .I(N__31395));
    LocalMux I__5939 (
            .O(N__31403),
            .I(N__31395));
    Span4Mux_h I__5938 (
            .O(N__31400),
            .I(N__31392));
    Odrv12 I__5937 (
            .O(N__31395),
            .I(red_c_i));
    Odrv4 I__5936 (
            .O(N__31392),
            .I(red_c_i));
    InMux I__5935 (
            .O(N__31387),
            .I(N__31384));
    LocalMux I__5934 (
            .O(N__31384),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ));
    InMux I__5933 (
            .O(N__31381),
            .I(N__31378));
    LocalMux I__5932 (
            .O(N__31378),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ));
    CascadeMux I__5931 (
            .O(N__31375),
            .I(N__31372));
    InMux I__5930 (
            .O(N__31372),
            .I(N__31369));
    LocalMux I__5929 (
            .O(N__31369),
            .I(N__31366));
    Span4Mux_h I__5928 (
            .O(N__31366),
            .I(N__31363));
    Span4Mux_v I__5927 (
            .O(N__31363),
            .I(N__31360));
    Odrv4 I__5926 (
            .O(N__31360),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ));
    CascadeMux I__5925 (
            .O(N__31357),
            .I(N__31352));
    CascadeMux I__5924 (
            .O(N__31356),
            .I(N__31349));
    InMux I__5923 (
            .O(N__31355),
            .I(N__31346));
    InMux I__5922 (
            .O(N__31352),
            .I(N__31341));
    InMux I__5921 (
            .O(N__31349),
            .I(N__31341));
    LocalMux I__5920 (
            .O(N__31346),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__5919 (
            .O(N__31341),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__5918 (
            .O(N__31336),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__5917 (
            .O(N__31333),
            .I(N__31328));
    InMux I__5916 (
            .O(N__31332),
            .I(N__31325));
    InMux I__5915 (
            .O(N__31331),
            .I(N__31322));
    LocalMux I__5914 (
            .O(N__31328),
            .I(N__31319));
    LocalMux I__5913 (
            .O(N__31325),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__5912 (
            .O(N__31322),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__5911 (
            .O(N__31319),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__5910 (
            .O(N__31312),
            .I(bfn_13_10_0_));
    InMux I__5909 (
            .O(N__31309),
            .I(N__31304));
    InMux I__5908 (
            .O(N__31308),
            .I(N__31301));
    InMux I__5907 (
            .O(N__31307),
            .I(N__31298));
    LocalMux I__5906 (
            .O(N__31304),
            .I(N__31295));
    LocalMux I__5905 (
            .O(N__31301),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__5904 (
            .O(N__31298),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__5903 (
            .O(N__31295),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__5902 (
            .O(N__31288),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__5901 (
            .O(N__31285),
            .I(N__31280));
    CascadeMux I__5900 (
            .O(N__31284),
            .I(N__31277));
    InMux I__5899 (
            .O(N__31283),
            .I(N__31274));
    InMux I__5898 (
            .O(N__31280),
            .I(N__31269));
    InMux I__5897 (
            .O(N__31277),
            .I(N__31269));
    LocalMux I__5896 (
            .O(N__31274),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__5895 (
            .O(N__31269),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__5894 (
            .O(N__31264),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__5893 (
            .O(N__31261),
            .I(N__31256));
    CascadeMux I__5892 (
            .O(N__31260),
            .I(N__31253));
    InMux I__5891 (
            .O(N__31259),
            .I(N__31250));
    InMux I__5890 (
            .O(N__31256),
            .I(N__31245));
    InMux I__5889 (
            .O(N__31253),
            .I(N__31245));
    LocalMux I__5888 (
            .O(N__31250),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__5887 (
            .O(N__31245),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__5886 (
            .O(N__31240),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__5885 (
            .O(N__31237),
            .I(N__31233));
    InMux I__5884 (
            .O(N__31236),
            .I(N__31230));
    LocalMux I__5883 (
            .O(N__31233),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__5882 (
            .O(N__31230),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__5881 (
            .O(N__31225),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__5880 (
            .O(N__31222),
            .I(N__31188));
    InMux I__5879 (
            .O(N__31221),
            .I(N__31188));
    InMux I__5878 (
            .O(N__31220),
            .I(N__31179));
    InMux I__5877 (
            .O(N__31219),
            .I(N__31179));
    InMux I__5876 (
            .O(N__31218),
            .I(N__31179));
    InMux I__5875 (
            .O(N__31217),
            .I(N__31179));
    InMux I__5874 (
            .O(N__31216),
            .I(N__31170));
    InMux I__5873 (
            .O(N__31215),
            .I(N__31170));
    InMux I__5872 (
            .O(N__31214),
            .I(N__31170));
    InMux I__5871 (
            .O(N__31213),
            .I(N__31170));
    InMux I__5870 (
            .O(N__31212),
            .I(N__31161));
    InMux I__5869 (
            .O(N__31211),
            .I(N__31161));
    InMux I__5868 (
            .O(N__31210),
            .I(N__31161));
    InMux I__5867 (
            .O(N__31209),
            .I(N__31161));
    InMux I__5866 (
            .O(N__31208),
            .I(N__31152));
    InMux I__5865 (
            .O(N__31207),
            .I(N__31152));
    InMux I__5864 (
            .O(N__31206),
            .I(N__31152));
    InMux I__5863 (
            .O(N__31205),
            .I(N__31152));
    InMux I__5862 (
            .O(N__31204),
            .I(N__31143));
    InMux I__5861 (
            .O(N__31203),
            .I(N__31143));
    InMux I__5860 (
            .O(N__31202),
            .I(N__31143));
    InMux I__5859 (
            .O(N__31201),
            .I(N__31143));
    InMux I__5858 (
            .O(N__31200),
            .I(N__31134));
    InMux I__5857 (
            .O(N__31199),
            .I(N__31134));
    InMux I__5856 (
            .O(N__31198),
            .I(N__31134));
    InMux I__5855 (
            .O(N__31197),
            .I(N__31134));
    InMux I__5854 (
            .O(N__31196),
            .I(N__31125));
    InMux I__5853 (
            .O(N__31195),
            .I(N__31125));
    InMux I__5852 (
            .O(N__31194),
            .I(N__31125));
    InMux I__5851 (
            .O(N__31193),
            .I(N__31125));
    LocalMux I__5850 (
            .O(N__31188),
            .I(N__31116));
    LocalMux I__5849 (
            .O(N__31179),
            .I(N__31116));
    LocalMux I__5848 (
            .O(N__31170),
            .I(N__31116));
    LocalMux I__5847 (
            .O(N__31161),
            .I(N__31116));
    LocalMux I__5846 (
            .O(N__31152),
            .I(N__31109));
    LocalMux I__5845 (
            .O(N__31143),
            .I(N__31109));
    LocalMux I__5844 (
            .O(N__31134),
            .I(N__31109));
    LocalMux I__5843 (
            .O(N__31125),
            .I(N__31104));
    Span4Mux_v I__5842 (
            .O(N__31116),
            .I(N__31104));
    Odrv12 I__5841 (
            .O(N__31109),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__5840 (
            .O(N__31104),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__5839 (
            .O(N__31099),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__5838 (
            .O(N__31096),
            .I(N__31092));
    InMux I__5837 (
            .O(N__31095),
            .I(N__31089));
    LocalMux I__5836 (
            .O(N__31092),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__5835 (
            .O(N__31089),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CEMux I__5834 (
            .O(N__31084),
            .I(N__31079));
    CEMux I__5833 (
            .O(N__31083),
            .I(N__31076));
    CEMux I__5832 (
            .O(N__31082),
            .I(N__31073));
    LocalMux I__5831 (
            .O(N__31079),
            .I(N__31069));
    LocalMux I__5830 (
            .O(N__31076),
            .I(N__31066));
    LocalMux I__5829 (
            .O(N__31073),
            .I(N__31063));
    CEMux I__5828 (
            .O(N__31072),
            .I(N__31060));
    Span4Mux_v I__5827 (
            .O(N__31069),
            .I(N__31055));
    Span4Mux_h I__5826 (
            .O(N__31066),
            .I(N__31055));
    Span4Mux_h I__5825 (
            .O(N__31063),
            .I(N__31052));
    LocalMux I__5824 (
            .O(N__31060),
            .I(N__31049));
    Span4Mux_h I__5823 (
            .O(N__31055),
            .I(N__31046));
    Span4Mux_h I__5822 (
            .O(N__31052),
            .I(N__31043));
    Span4Mux_h I__5821 (
            .O(N__31049),
            .I(N__31040));
    Odrv4 I__5820 (
            .O(N__31046),
            .I(\delay_measurement_inst.delay_hc_timer.N_337_i ));
    Odrv4 I__5819 (
            .O(N__31043),
            .I(\delay_measurement_inst.delay_hc_timer.N_337_i ));
    Odrv4 I__5818 (
            .O(N__31040),
            .I(\delay_measurement_inst.delay_hc_timer.N_337_i ));
    CascadeMux I__5817 (
            .O(N__31033),
            .I(N__31029));
    InMux I__5816 (
            .O(N__31032),
            .I(N__31025));
    InMux I__5815 (
            .O(N__31029),
            .I(N__31022));
    InMux I__5814 (
            .O(N__31028),
            .I(N__31018));
    LocalMux I__5813 (
            .O(N__31025),
            .I(N__31015));
    LocalMux I__5812 (
            .O(N__31022),
            .I(N__31012));
    InMux I__5811 (
            .O(N__31021),
            .I(N__31009));
    LocalMux I__5810 (
            .O(N__31018),
            .I(N__31005));
    Span4Mux_v I__5809 (
            .O(N__31015),
            .I(N__31002));
    Span4Mux_h I__5808 (
            .O(N__31012),
            .I(N__30999));
    LocalMux I__5807 (
            .O(N__31009),
            .I(N__30996));
    InMux I__5806 (
            .O(N__31008),
            .I(N__30993));
    Span4Mux_s3_v I__5805 (
            .O(N__31005),
            .I(N__30989));
    Span4Mux_h I__5804 (
            .O(N__31002),
            .I(N__30985));
    Span4Mux_h I__5803 (
            .O(N__30999),
            .I(N__30977));
    Span4Mux_v I__5802 (
            .O(N__30996),
            .I(N__30977));
    LocalMux I__5801 (
            .O(N__30993),
            .I(N__30977));
    InMux I__5800 (
            .O(N__30992),
            .I(N__30974));
    Span4Mux_v I__5799 (
            .O(N__30989),
            .I(N__30971));
    InMux I__5798 (
            .O(N__30988),
            .I(N__30968));
    Sp12to4 I__5797 (
            .O(N__30985),
            .I(N__30965));
    InMux I__5796 (
            .O(N__30984),
            .I(N__30962));
    Span4Mux_h I__5795 (
            .O(N__30977),
            .I(N__30957));
    LocalMux I__5794 (
            .O(N__30974),
            .I(N__30957));
    Sp12to4 I__5793 (
            .O(N__30971),
            .I(N__30954));
    LocalMux I__5792 (
            .O(N__30968),
            .I(N__30951));
    Span12Mux_v I__5791 (
            .O(N__30965),
            .I(N__30948));
    LocalMux I__5790 (
            .O(N__30962),
            .I(N__30945));
    Span4Mux_v I__5789 (
            .O(N__30957),
            .I(N__30942));
    Span12Mux_h I__5788 (
            .O(N__30954),
            .I(N__30939));
    Span12Mux_s6_h I__5787 (
            .O(N__30951),
            .I(N__30936));
    Span12Mux_v I__5786 (
            .O(N__30948),
            .I(N__30933));
    Span12Mux_h I__5785 (
            .O(N__30945),
            .I(N__30930));
    Span4Mux_h I__5784 (
            .O(N__30942),
            .I(N__30927));
    Span12Mux_v I__5783 (
            .O(N__30939),
            .I(N__30922));
    Span12Mux_h I__5782 (
            .O(N__30936),
            .I(N__30922));
    Span12Mux_h I__5781 (
            .O(N__30933),
            .I(N__30917));
    Span12Mux_v I__5780 (
            .O(N__30930),
            .I(N__30917));
    Span4Mux_v I__5779 (
            .O(N__30927),
            .I(N__30914));
    Odrv12 I__5778 (
            .O(N__30922),
            .I(start_stop_c));
    Odrv12 I__5777 (
            .O(N__30917),
            .I(start_stop_c));
    Odrv4 I__5776 (
            .O(N__30914),
            .I(start_stop_c));
    CascadeMux I__5775 (
            .O(N__30907),
            .I(N__30902));
    CascadeMux I__5774 (
            .O(N__30906),
            .I(N__30899));
    InMux I__5773 (
            .O(N__30905),
            .I(N__30896));
    InMux I__5772 (
            .O(N__30902),
            .I(N__30891));
    InMux I__5771 (
            .O(N__30899),
            .I(N__30891));
    LocalMux I__5770 (
            .O(N__30896),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__5769 (
            .O(N__30891),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__5768 (
            .O(N__30886),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__5767 (
            .O(N__30883),
            .I(N__30878));
    InMux I__5766 (
            .O(N__30882),
            .I(N__30875));
    InMux I__5765 (
            .O(N__30881),
            .I(N__30872));
    LocalMux I__5764 (
            .O(N__30878),
            .I(N__30869));
    LocalMux I__5763 (
            .O(N__30875),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__5762 (
            .O(N__30872),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__5761 (
            .O(N__30869),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__5760 (
            .O(N__30862),
            .I(bfn_13_9_0_));
    InMux I__5759 (
            .O(N__30859),
            .I(N__30854));
    InMux I__5758 (
            .O(N__30858),
            .I(N__30851));
    InMux I__5757 (
            .O(N__30857),
            .I(N__30848));
    LocalMux I__5756 (
            .O(N__30854),
            .I(N__30845));
    LocalMux I__5755 (
            .O(N__30851),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__5754 (
            .O(N__30848),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__5753 (
            .O(N__30845),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__5752 (
            .O(N__30838),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    CascadeMux I__5751 (
            .O(N__30835),
            .I(N__30830));
    CascadeMux I__5750 (
            .O(N__30834),
            .I(N__30827));
    InMux I__5749 (
            .O(N__30833),
            .I(N__30824));
    InMux I__5748 (
            .O(N__30830),
            .I(N__30819));
    InMux I__5747 (
            .O(N__30827),
            .I(N__30819));
    LocalMux I__5746 (
            .O(N__30824),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__5745 (
            .O(N__30819),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__5744 (
            .O(N__30814),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    CascadeMux I__5743 (
            .O(N__30811),
            .I(N__30806));
    CascadeMux I__5742 (
            .O(N__30810),
            .I(N__30803));
    InMux I__5741 (
            .O(N__30809),
            .I(N__30800));
    InMux I__5740 (
            .O(N__30806),
            .I(N__30795));
    InMux I__5739 (
            .O(N__30803),
            .I(N__30795));
    LocalMux I__5738 (
            .O(N__30800),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__5737 (
            .O(N__30795),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__5736 (
            .O(N__30790),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__5735 (
            .O(N__30787),
            .I(N__30782));
    InMux I__5734 (
            .O(N__30786),
            .I(N__30777));
    InMux I__5733 (
            .O(N__30785),
            .I(N__30777));
    LocalMux I__5732 (
            .O(N__30782),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__5731 (
            .O(N__30777),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__5730 (
            .O(N__30772),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__5729 (
            .O(N__30769),
            .I(N__30764));
    InMux I__5728 (
            .O(N__30768),
            .I(N__30759));
    InMux I__5727 (
            .O(N__30767),
            .I(N__30759));
    LocalMux I__5726 (
            .O(N__30764),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__5725 (
            .O(N__30759),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__5724 (
            .O(N__30754),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    CascadeMux I__5723 (
            .O(N__30751),
            .I(N__30746));
    CascadeMux I__5722 (
            .O(N__30750),
            .I(N__30743));
    InMux I__5721 (
            .O(N__30749),
            .I(N__30740));
    InMux I__5720 (
            .O(N__30746),
            .I(N__30735));
    InMux I__5719 (
            .O(N__30743),
            .I(N__30735));
    LocalMux I__5718 (
            .O(N__30740),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__5717 (
            .O(N__30735),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__5716 (
            .O(N__30730),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    CascadeMux I__5715 (
            .O(N__30727),
            .I(N__30722));
    CascadeMux I__5714 (
            .O(N__30726),
            .I(N__30719));
    InMux I__5713 (
            .O(N__30725),
            .I(N__30716));
    InMux I__5712 (
            .O(N__30722),
            .I(N__30711));
    InMux I__5711 (
            .O(N__30719),
            .I(N__30711));
    LocalMux I__5710 (
            .O(N__30716),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__5709 (
            .O(N__30711),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__5708 (
            .O(N__30706),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    CascadeMux I__5707 (
            .O(N__30703),
            .I(N__30698));
    CascadeMux I__5706 (
            .O(N__30702),
            .I(N__30695));
    InMux I__5705 (
            .O(N__30701),
            .I(N__30692));
    InMux I__5704 (
            .O(N__30698),
            .I(N__30687));
    InMux I__5703 (
            .O(N__30695),
            .I(N__30687));
    LocalMux I__5702 (
            .O(N__30692),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__5701 (
            .O(N__30687),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__5700 (
            .O(N__30682),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__5699 (
            .O(N__30679),
            .I(N__30674));
    InMux I__5698 (
            .O(N__30678),
            .I(N__30671));
    InMux I__5697 (
            .O(N__30677),
            .I(N__30668));
    LocalMux I__5696 (
            .O(N__30674),
            .I(N__30665));
    LocalMux I__5695 (
            .O(N__30671),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__5694 (
            .O(N__30668),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__5693 (
            .O(N__30665),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__5692 (
            .O(N__30658),
            .I(bfn_13_8_0_));
    InMux I__5691 (
            .O(N__30655),
            .I(N__30650));
    InMux I__5690 (
            .O(N__30654),
            .I(N__30647));
    InMux I__5689 (
            .O(N__30653),
            .I(N__30644));
    LocalMux I__5688 (
            .O(N__30650),
            .I(N__30641));
    LocalMux I__5687 (
            .O(N__30647),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__5686 (
            .O(N__30644),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__5685 (
            .O(N__30641),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__5684 (
            .O(N__30634),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    CascadeMux I__5683 (
            .O(N__30631),
            .I(N__30626));
    CascadeMux I__5682 (
            .O(N__30630),
            .I(N__30623));
    InMux I__5681 (
            .O(N__30629),
            .I(N__30620));
    InMux I__5680 (
            .O(N__30626),
            .I(N__30615));
    InMux I__5679 (
            .O(N__30623),
            .I(N__30615));
    LocalMux I__5678 (
            .O(N__30620),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__5677 (
            .O(N__30615),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__5676 (
            .O(N__30610),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    CascadeMux I__5675 (
            .O(N__30607),
            .I(N__30602));
    CascadeMux I__5674 (
            .O(N__30606),
            .I(N__30599));
    InMux I__5673 (
            .O(N__30605),
            .I(N__30596));
    InMux I__5672 (
            .O(N__30602),
            .I(N__30591));
    InMux I__5671 (
            .O(N__30599),
            .I(N__30591));
    LocalMux I__5670 (
            .O(N__30596),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__5669 (
            .O(N__30591),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__5668 (
            .O(N__30586),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__5667 (
            .O(N__30583),
            .I(N__30578));
    InMux I__5666 (
            .O(N__30582),
            .I(N__30573));
    InMux I__5665 (
            .O(N__30581),
            .I(N__30573));
    LocalMux I__5664 (
            .O(N__30578),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__5663 (
            .O(N__30573),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__5662 (
            .O(N__30568),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__5661 (
            .O(N__30565),
            .I(N__30560));
    InMux I__5660 (
            .O(N__30564),
            .I(N__30555));
    InMux I__5659 (
            .O(N__30563),
            .I(N__30555));
    LocalMux I__5658 (
            .O(N__30560),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__5657 (
            .O(N__30555),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__5656 (
            .O(N__30550),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    CascadeMux I__5655 (
            .O(N__30547),
            .I(N__30542));
    CascadeMux I__5654 (
            .O(N__30546),
            .I(N__30539));
    InMux I__5653 (
            .O(N__30545),
            .I(N__30536));
    InMux I__5652 (
            .O(N__30542),
            .I(N__30531));
    InMux I__5651 (
            .O(N__30539),
            .I(N__30531));
    LocalMux I__5650 (
            .O(N__30536),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__5649 (
            .O(N__30531),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__5648 (
            .O(N__30526),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__5647 (
            .O(N__30523),
            .I(N__30520));
    LocalMux I__5646 (
            .O(N__30520),
            .I(N__30516));
    CascadeMux I__5645 (
            .O(N__30519),
            .I(N__30512));
    Span4Mux_v I__5644 (
            .O(N__30516),
            .I(N__30508));
    InMux I__5643 (
            .O(N__30515),
            .I(N__30505));
    InMux I__5642 (
            .O(N__30512),
            .I(N__30502));
    InMux I__5641 (
            .O(N__30511),
            .I(N__30499));
    Odrv4 I__5640 (
            .O(N__30508),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__5639 (
            .O(N__30505),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__5638 (
            .O(N__30502),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__5637 (
            .O(N__30499),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    InMux I__5636 (
            .O(N__30490),
            .I(N__30487));
    LocalMux I__5635 (
            .O(N__30487),
            .I(N__30477));
    InMux I__5634 (
            .O(N__30486),
            .I(N__30474));
    InMux I__5633 (
            .O(N__30485),
            .I(N__30469));
    InMux I__5632 (
            .O(N__30484),
            .I(N__30469));
    InMux I__5631 (
            .O(N__30483),
            .I(N__30460));
    InMux I__5630 (
            .O(N__30482),
            .I(N__30460));
    InMux I__5629 (
            .O(N__30481),
            .I(N__30460));
    InMux I__5628 (
            .O(N__30480),
            .I(N__30457));
    Span4Mux_v I__5627 (
            .O(N__30477),
            .I(N__30452));
    LocalMux I__5626 (
            .O(N__30474),
            .I(N__30449));
    LocalMux I__5625 (
            .O(N__30469),
            .I(N__30446));
    InMux I__5624 (
            .O(N__30468),
            .I(N__30441));
    InMux I__5623 (
            .O(N__30467),
            .I(N__30441));
    LocalMux I__5622 (
            .O(N__30460),
            .I(N__30438));
    LocalMux I__5621 (
            .O(N__30457),
            .I(N__30434));
    InMux I__5620 (
            .O(N__30456),
            .I(N__30429));
    InMux I__5619 (
            .O(N__30455),
            .I(N__30429));
    Span4Mux_v I__5618 (
            .O(N__30452),
            .I(N__30411));
    Span4Mux_v I__5617 (
            .O(N__30449),
            .I(N__30411));
    Span4Mux_v I__5616 (
            .O(N__30446),
            .I(N__30411));
    LocalMux I__5615 (
            .O(N__30441),
            .I(N__30408));
    Span4Mux_h I__5614 (
            .O(N__30438),
            .I(N__30405));
    InMux I__5613 (
            .O(N__30437),
            .I(N__30402));
    Span4Mux_v I__5612 (
            .O(N__30434),
            .I(N__30397));
    LocalMux I__5611 (
            .O(N__30429),
            .I(N__30397));
    InMux I__5610 (
            .O(N__30428),
            .I(N__30382));
    InMux I__5609 (
            .O(N__30427),
            .I(N__30382));
    InMux I__5608 (
            .O(N__30426),
            .I(N__30382));
    InMux I__5607 (
            .O(N__30425),
            .I(N__30382));
    InMux I__5606 (
            .O(N__30424),
            .I(N__30382));
    InMux I__5605 (
            .O(N__30423),
            .I(N__30382));
    InMux I__5604 (
            .O(N__30422),
            .I(N__30382));
    InMux I__5603 (
            .O(N__30421),
            .I(N__30373));
    InMux I__5602 (
            .O(N__30420),
            .I(N__30373));
    InMux I__5601 (
            .O(N__30419),
            .I(N__30373));
    InMux I__5600 (
            .O(N__30418),
            .I(N__30373));
    Odrv4 I__5599 (
            .O(N__30411),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv4 I__5598 (
            .O(N__30408),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv4 I__5597 (
            .O(N__30405),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__5596 (
            .O(N__30402),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv4 I__5595 (
            .O(N__30397),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__5594 (
            .O(N__30382),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__5593 (
            .O(N__30373),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    InMux I__5592 (
            .O(N__30358),
            .I(N__30353));
    InMux I__5591 (
            .O(N__30357),
            .I(N__30350));
    InMux I__5590 (
            .O(N__30356),
            .I(N__30347));
    LocalMux I__5589 (
            .O(N__30353),
            .I(N__30344));
    LocalMux I__5588 (
            .O(N__30350),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    LocalMux I__5587 (
            .O(N__30347),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    Odrv12 I__5586 (
            .O(N__30344),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    InMux I__5585 (
            .O(N__30337),
            .I(N__30332));
    InMux I__5584 (
            .O(N__30336),
            .I(N__30329));
    InMux I__5583 (
            .O(N__30335),
            .I(N__30326));
    LocalMux I__5582 (
            .O(N__30332),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__5581 (
            .O(N__30329),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__5580 (
            .O(N__30326),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__5579 (
            .O(N__30319),
            .I(bfn_13_7_0_));
    InMux I__5578 (
            .O(N__30316),
            .I(N__30311));
    InMux I__5577 (
            .O(N__30315),
            .I(N__30308));
    InMux I__5576 (
            .O(N__30314),
            .I(N__30305));
    LocalMux I__5575 (
            .O(N__30311),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__5574 (
            .O(N__30308),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__5573 (
            .O(N__30305),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__5572 (
            .O(N__30298),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    CascadeMux I__5571 (
            .O(N__30295),
            .I(N__30290));
    CascadeMux I__5570 (
            .O(N__30294),
            .I(N__30287));
    InMux I__5569 (
            .O(N__30293),
            .I(N__30284));
    InMux I__5568 (
            .O(N__30290),
            .I(N__30279));
    InMux I__5567 (
            .O(N__30287),
            .I(N__30279));
    LocalMux I__5566 (
            .O(N__30284),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__5565 (
            .O(N__30279),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__5564 (
            .O(N__30274),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    CascadeMux I__5563 (
            .O(N__30271),
            .I(N__30266));
    CascadeMux I__5562 (
            .O(N__30270),
            .I(N__30263));
    InMux I__5561 (
            .O(N__30269),
            .I(N__30260));
    InMux I__5560 (
            .O(N__30266),
            .I(N__30255));
    InMux I__5559 (
            .O(N__30263),
            .I(N__30255));
    LocalMux I__5558 (
            .O(N__30260),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__5557 (
            .O(N__30255),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__5556 (
            .O(N__30250),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__5555 (
            .O(N__30247),
            .I(N__30242));
    InMux I__5554 (
            .O(N__30246),
            .I(N__30237));
    InMux I__5553 (
            .O(N__30245),
            .I(N__30237));
    LocalMux I__5552 (
            .O(N__30242),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__5551 (
            .O(N__30237),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__5550 (
            .O(N__30232),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__5549 (
            .O(N__30229),
            .I(N__30224));
    InMux I__5548 (
            .O(N__30228),
            .I(N__30219));
    InMux I__5547 (
            .O(N__30227),
            .I(N__30219));
    LocalMux I__5546 (
            .O(N__30224),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__5545 (
            .O(N__30219),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__5544 (
            .O(N__30214),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__5543 (
            .O(N__30211),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__5542 (
            .O(N__30208),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__5541 (
            .O(N__30205),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__5540 (
            .O(N__30202),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    CascadeMux I__5539 (
            .O(N__30199),
            .I(N__30196));
    InMux I__5538 (
            .O(N__30196),
            .I(N__30193));
    LocalMux I__5537 (
            .O(N__30193),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ));
    InMux I__5536 (
            .O(N__30190),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__5535 (
            .O(N__30187),
            .I(bfn_12_26_0_));
    InMux I__5534 (
            .O(N__30184),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__5533 (
            .O(N__30181),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__5532 (
            .O(N__30178),
            .I(N__30175));
    LocalMux I__5531 (
            .O(N__30175),
            .I(N__30169));
    InMux I__5530 (
            .O(N__30174),
            .I(N__30166));
    InMux I__5529 (
            .O(N__30173),
            .I(N__30163));
    InMux I__5528 (
            .O(N__30172),
            .I(N__30160));
    Span4Mux_h I__5527 (
            .O(N__30169),
            .I(N__30157));
    LocalMux I__5526 (
            .O(N__30166),
            .I(N__30154));
    LocalMux I__5525 (
            .O(N__30163),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__5524 (
            .O(N__30160),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__5523 (
            .O(N__30157),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__5522 (
            .O(N__30154),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__5521 (
            .O(N__30145),
            .I(N__30142));
    LocalMux I__5520 (
            .O(N__30142),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ));
    InMux I__5519 (
            .O(N__30139),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__5518 (
            .O(N__30136),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__5517 (
            .O(N__30133),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__5516 (
            .O(N__30130),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__5515 (
            .O(N__30127),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__5514 (
            .O(N__30124),
            .I(N__30121));
    LocalMux I__5513 (
            .O(N__30121),
            .I(N__30118));
    Odrv12 I__5512 (
            .O(N__30118),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ));
    InMux I__5511 (
            .O(N__30115),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__5510 (
            .O(N__30112),
            .I(N__30109));
    LocalMux I__5509 (
            .O(N__30109),
            .I(N__30106));
    Odrv12 I__5508 (
            .O(N__30106),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ));
    InMux I__5507 (
            .O(N__30103),
            .I(bfn_12_25_0_));
    InMux I__5506 (
            .O(N__30100),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__5505 (
            .O(N__30097),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    CascadeMux I__5504 (
            .O(N__30094),
            .I(N__30090));
    InMux I__5503 (
            .O(N__30093),
            .I(N__30087));
    InMux I__5502 (
            .O(N__30090),
            .I(N__30084));
    LocalMux I__5501 (
            .O(N__30087),
            .I(\current_shift_inst.z_i_31 ));
    LocalMux I__5500 (
            .O(N__30084),
            .I(\current_shift_inst.z_i_31 ));
    InMux I__5499 (
            .O(N__30079),
            .I(N__30076));
    LocalMux I__5498 (
            .O(N__30076),
            .I(N__30073));
    Odrv4 I__5497 (
            .O(N__30073),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ));
    IoInMux I__5496 (
            .O(N__30070),
            .I(N__30067));
    LocalMux I__5495 (
            .O(N__30067),
            .I(N__30064));
    Span4Mux_s2_v I__5494 (
            .O(N__30064),
            .I(N__30061));
    Span4Mux_v I__5493 (
            .O(N__30061),
            .I(N__30058));
    Odrv4 I__5492 (
            .O(N__30058),
            .I(\current_shift_inst.timer_phase.N_188_i ));
    InMux I__5491 (
            .O(N__30055),
            .I(N__30052));
    LocalMux I__5490 (
            .O(N__30052),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    InMux I__5489 (
            .O(N__30049),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    IoInMux I__5488 (
            .O(N__30046),
            .I(N__30043));
    LocalMux I__5487 (
            .O(N__30043),
            .I(N__30040));
    Span4Mux_s3_v I__5486 (
            .O(N__30040),
            .I(N__30037));
    Span4Mux_h I__5485 (
            .O(N__30037),
            .I(N__30034));
    Sp12to4 I__5484 (
            .O(N__30034),
            .I(N__30031));
    Span12Mux_v I__5483 (
            .O(N__30031),
            .I(N__30027));
    InMux I__5482 (
            .O(N__30030),
            .I(N__30024));
    Odrv12 I__5481 (
            .O(N__30027),
            .I(s1_phy_c));
    LocalMux I__5480 (
            .O(N__30024),
            .I(s1_phy_c));
    InMux I__5479 (
            .O(N__30019),
            .I(N__30016));
    LocalMux I__5478 (
            .O(N__30016),
            .I(N__30013));
    Span4Mux_v I__5477 (
            .O(N__30013),
            .I(N__30010));
    Span4Mux_v I__5476 (
            .O(N__30010),
            .I(N__30007));
    Odrv4 I__5475 (
            .O(N__30007),
            .I(\phase_controller_inst1.stoper_tr.N_21 ));
    InMux I__5474 (
            .O(N__30004),
            .I(N__30001));
    LocalMux I__5473 (
            .O(N__30001),
            .I(N__29998));
    Odrv4 I__5472 (
            .O(N__29998),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3 ));
    InMux I__5471 (
            .O(N__29995),
            .I(N__29992));
    LocalMux I__5470 (
            .O(N__29992),
            .I(N__29987));
    InMux I__5469 (
            .O(N__29991),
            .I(N__29982));
    InMux I__5468 (
            .O(N__29990),
            .I(N__29982));
    Odrv4 I__5467 (
            .O(N__29987),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    LocalMux I__5466 (
            .O(N__29982),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    InMux I__5465 (
            .O(N__29977),
            .I(N__29974));
    LocalMux I__5464 (
            .O(N__29974),
            .I(N__29971));
    Span4Mux_h I__5463 (
            .O(N__29971),
            .I(N__29965));
    InMux I__5462 (
            .O(N__29970),
            .I(N__29962));
    InMux I__5461 (
            .O(N__29969),
            .I(N__29959));
    InMux I__5460 (
            .O(N__29968),
            .I(N__29956));
    Odrv4 I__5459 (
            .O(N__29965),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__5458 (
            .O(N__29962),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__5457 (
            .O(N__29959),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__5456 (
            .O(N__29956),
            .I(\phase_controller_inst1.hc_time_passed ));
    CascadeMux I__5455 (
            .O(N__29947),
            .I(N__29943));
    InMux I__5454 (
            .O(N__29946),
            .I(N__29940));
    InMux I__5453 (
            .O(N__29943),
            .I(N__29937));
    LocalMux I__5452 (
            .O(N__29940),
            .I(N__29933));
    LocalMux I__5451 (
            .O(N__29937),
            .I(N__29930));
    CascadeMux I__5450 (
            .O(N__29936),
            .I(N__29927));
    Span4Mux_h I__5449 (
            .O(N__29933),
            .I(N__29923));
    Span4Mux_h I__5448 (
            .O(N__29930),
            .I(N__29920));
    InMux I__5447 (
            .O(N__29927),
            .I(N__29917));
    InMux I__5446 (
            .O(N__29926),
            .I(N__29914));
    Odrv4 I__5445 (
            .O(N__29923),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__5444 (
            .O(N__29920),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__5443 (
            .O(N__29917),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__5442 (
            .O(N__29914),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__5441 (
            .O(N__29905),
            .I(N__29900));
    InMux I__5440 (
            .O(N__29904),
            .I(N__29897));
    InMux I__5439 (
            .O(N__29903),
            .I(N__29894));
    LocalMux I__5438 (
            .O(N__29900),
            .I(N__29891));
    LocalMux I__5437 (
            .O(N__29897),
            .I(N__29886));
    LocalMux I__5436 (
            .O(N__29894),
            .I(N__29886));
    Odrv4 I__5435 (
            .O(N__29891),
            .I(il_min_comp1_D2));
    Odrv4 I__5434 (
            .O(N__29886),
            .I(il_min_comp1_D2));
    InMux I__5433 (
            .O(N__29881),
            .I(N__29874));
    InMux I__5432 (
            .O(N__29880),
            .I(N__29871));
    CascadeMux I__5431 (
            .O(N__29879),
            .I(N__29868));
    CascadeMux I__5430 (
            .O(N__29878),
            .I(N__29865));
    CascadeMux I__5429 (
            .O(N__29877),
            .I(N__29862));
    LocalMux I__5428 (
            .O(N__29874),
            .I(N__29857));
    LocalMux I__5427 (
            .O(N__29871),
            .I(N__29857));
    InMux I__5426 (
            .O(N__29868),
            .I(N__29854));
    InMux I__5425 (
            .O(N__29865),
            .I(N__29851));
    InMux I__5424 (
            .O(N__29862),
            .I(N__29848));
    Span12Mux_v I__5423 (
            .O(N__29857),
            .I(N__29845));
    LocalMux I__5422 (
            .O(N__29854),
            .I(N__29840));
    LocalMux I__5421 (
            .O(N__29851),
            .I(N__29840));
    LocalMux I__5420 (
            .O(N__29848),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv12 I__5419 (
            .O(N__29845),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv4 I__5418 (
            .O(N__29840),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__5417 (
            .O(N__29833),
            .I(N__29829));
    InMux I__5416 (
            .O(N__29832),
            .I(N__29826));
    LocalMux I__5415 (
            .O(N__29829),
            .I(N__29823));
    LocalMux I__5414 (
            .O(N__29826),
            .I(N__29819));
    Span4Mux_h I__5413 (
            .O(N__29823),
            .I(N__29816));
    InMux I__5412 (
            .O(N__29822),
            .I(N__29812));
    Span4Mux_h I__5411 (
            .O(N__29819),
            .I(N__29807));
    Span4Mux_v I__5410 (
            .O(N__29816),
            .I(N__29807));
    InMux I__5409 (
            .O(N__29815),
            .I(N__29804));
    LocalMux I__5408 (
            .O(N__29812),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv4 I__5407 (
            .O(N__29807),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__5406 (
            .O(N__29804),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    InMux I__5405 (
            .O(N__29797),
            .I(N__29794));
    LocalMux I__5404 (
            .O(N__29794),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__5403 (
            .O(N__29791),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__5402 (
            .O(N__29788),
            .I(N__29785));
    LocalMux I__5401 (
            .O(N__29785),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__5400 (
            .O(N__29782),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__5399 (
            .O(N__29779),
            .I(N__29776));
    InMux I__5398 (
            .O(N__29776),
            .I(N__29773));
    LocalMux I__5397 (
            .O(N__29773),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__5396 (
            .O(N__29770),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__5395 (
            .O(N__29767),
            .I(N__29764));
    LocalMux I__5394 (
            .O(N__29764),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__5393 (
            .O(N__29761),
            .I(bfn_12_10_0_));
    InMux I__5392 (
            .O(N__29758),
            .I(N__29755));
    LocalMux I__5391 (
            .O(N__29755),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__5390 (
            .O(N__29752),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__5389 (
            .O(N__29749),
            .I(N__29746));
    LocalMux I__5388 (
            .O(N__29746),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__5387 (
            .O(N__29743),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__5386 (
            .O(N__29740),
            .I(N__29737));
    InMux I__5385 (
            .O(N__29737),
            .I(N__29734));
    LocalMux I__5384 (
            .O(N__29734),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__5383 (
            .O(N__29731),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__5382 (
            .O(N__29728),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__5381 (
            .O(N__29725),
            .I(N__29722));
    InMux I__5380 (
            .O(N__29722),
            .I(N__29715));
    InMux I__5379 (
            .O(N__29721),
            .I(N__29715));
    CascadeMux I__5378 (
            .O(N__29720),
            .I(N__29712));
    LocalMux I__5377 (
            .O(N__29715),
            .I(N__29709));
    InMux I__5376 (
            .O(N__29712),
            .I(N__29706));
    Span4Mux_h I__5375 (
            .O(N__29709),
            .I(N__29703));
    LocalMux I__5374 (
            .O(N__29706),
            .I(N__29700));
    Odrv4 I__5373 (
            .O(N__29703),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__5372 (
            .O(N__29700),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    CEMux I__5371 (
            .O(N__29695),
            .I(N__29680));
    CEMux I__5370 (
            .O(N__29694),
            .I(N__29680));
    CEMux I__5369 (
            .O(N__29693),
            .I(N__29680));
    CEMux I__5368 (
            .O(N__29692),
            .I(N__29680));
    CEMux I__5367 (
            .O(N__29691),
            .I(N__29680));
    GlobalMux I__5366 (
            .O(N__29680),
            .I(N__29677));
    gio2CtrlBuf I__5365 (
            .O(N__29677),
            .I(\delay_measurement_inst.delay_hc_timer.N_336_i_g ));
    InMux I__5364 (
            .O(N__29674),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__5363 (
            .O(N__29671),
            .I(N__29668));
    LocalMux I__5362 (
            .O(N__29668),
            .I(N__29665));
    Span4Mux_h I__5361 (
            .O(N__29665),
            .I(N__29660));
    InMux I__5360 (
            .O(N__29664),
            .I(N__29657));
    InMux I__5359 (
            .O(N__29663),
            .I(N__29654));
    Odrv4 I__5358 (
            .O(N__29660),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    LocalMux I__5357 (
            .O(N__29657),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    LocalMux I__5356 (
            .O(N__29654),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    InMux I__5355 (
            .O(N__29647),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__5354 (
            .O(N__29644),
            .I(N__29641));
    LocalMux I__5353 (
            .O(N__29641),
            .I(N__29638));
    Span4Mux_h I__5352 (
            .O(N__29638),
            .I(N__29633));
    InMux I__5351 (
            .O(N__29637),
            .I(N__29630));
    InMux I__5350 (
            .O(N__29636),
            .I(N__29627));
    Odrv4 I__5349 (
            .O(N__29633),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    LocalMux I__5348 (
            .O(N__29630),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    LocalMux I__5347 (
            .O(N__29627),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    InMux I__5346 (
            .O(N__29620),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__5345 (
            .O(N__29617),
            .I(N__29612));
    InMux I__5344 (
            .O(N__29616),
            .I(N__29609));
    CascadeMux I__5343 (
            .O(N__29615),
            .I(N__29606));
    LocalMux I__5342 (
            .O(N__29612),
            .I(N__29603));
    LocalMux I__5341 (
            .O(N__29609),
            .I(N__29600));
    InMux I__5340 (
            .O(N__29606),
            .I(N__29597));
    Odrv12 I__5339 (
            .O(N__29603),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    Odrv4 I__5338 (
            .O(N__29600),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    LocalMux I__5337 (
            .O(N__29597),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    InMux I__5336 (
            .O(N__29590),
            .I(bfn_12_9_0_));
    InMux I__5335 (
            .O(N__29587),
            .I(N__29583));
    InMux I__5334 (
            .O(N__29586),
            .I(N__29580));
    LocalMux I__5333 (
            .O(N__29583),
            .I(N__29577));
    LocalMux I__5332 (
            .O(N__29580),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    Odrv4 I__5331 (
            .O(N__29577),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__5330 (
            .O(N__29572),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__5329 (
            .O(N__29569),
            .I(N__29563));
    InMux I__5328 (
            .O(N__29568),
            .I(N__29563));
    LocalMux I__5327 (
            .O(N__29563),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__5326 (
            .O(N__29560),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__5325 (
            .O(N__29557),
            .I(N__29554));
    InMux I__5324 (
            .O(N__29554),
            .I(N__29548));
    InMux I__5323 (
            .O(N__29553),
            .I(N__29548));
    LocalMux I__5322 (
            .O(N__29548),
            .I(N__29545));
    Odrv4 I__5321 (
            .O(N__29545),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__5320 (
            .O(N__29542),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__5319 (
            .O(N__29539),
            .I(N__29536));
    LocalMux I__5318 (
            .O(N__29536),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__5317 (
            .O(N__29533),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__5316 (
            .O(N__29530),
            .I(N__29525));
    InMux I__5315 (
            .O(N__29529),
            .I(N__29522));
    InMux I__5314 (
            .O(N__29528),
            .I(N__29519));
    LocalMux I__5313 (
            .O(N__29525),
            .I(N__29512));
    LocalMux I__5312 (
            .O(N__29522),
            .I(N__29512));
    LocalMux I__5311 (
            .O(N__29519),
            .I(N__29512));
    Span4Mux_v I__5310 (
            .O(N__29512),
            .I(N__29508));
    InMux I__5309 (
            .O(N__29511),
            .I(N__29505));
    Odrv4 I__5308 (
            .O(N__29508),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__5307 (
            .O(N__29505),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    InMux I__5306 (
            .O(N__29500),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__5305 (
            .O(N__29497),
            .I(N__29492));
    InMux I__5304 (
            .O(N__29496),
            .I(N__29489));
    InMux I__5303 (
            .O(N__29495),
            .I(N__29486));
    InMux I__5302 (
            .O(N__29492),
            .I(N__29483));
    LocalMux I__5301 (
            .O(N__29489),
            .I(N__29476));
    LocalMux I__5300 (
            .O(N__29486),
            .I(N__29476));
    LocalMux I__5299 (
            .O(N__29483),
            .I(N__29476));
    Span4Mux_v I__5298 (
            .O(N__29476),
            .I(N__29472));
    InMux I__5297 (
            .O(N__29475),
            .I(N__29469));
    Odrv4 I__5296 (
            .O(N__29472),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__5295 (
            .O(N__29469),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    InMux I__5294 (
            .O(N__29464),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__5293 (
            .O(N__29461),
            .I(N__29458));
    LocalMux I__5292 (
            .O(N__29458),
            .I(N__29453));
    InMux I__5291 (
            .O(N__29457),
            .I(N__29450));
    InMux I__5290 (
            .O(N__29456),
            .I(N__29447));
    Span4Mux_v I__5289 (
            .O(N__29453),
            .I(N__29442));
    LocalMux I__5288 (
            .O(N__29450),
            .I(N__29442));
    LocalMux I__5287 (
            .O(N__29447),
            .I(N__29439));
    Span4Mux_h I__5286 (
            .O(N__29442),
            .I(N__29435));
    Span4Mux_h I__5285 (
            .O(N__29439),
            .I(N__29432));
    InMux I__5284 (
            .O(N__29438),
            .I(N__29429));
    Odrv4 I__5283 (
            .O(N__29435),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    Odrv4 I__5282 (
            .O(N__29432),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__5281 (
            .O(N__29429),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    InMux I__5280 (
            .O(N__29422),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__5279 (
            .O(N__29419),
            .I(N__29416));
    InMux I__5278 (
            .O(N__29416),
            .I(N__29412));
    InMux I__5277 (
            .O(N__29415),
            .I(N__29409));
    LocalMux I__5276 (
            .O(N__29412),
            .I(N__29406));
    LocalMux I__5275 (
            .O(N__29409),
            .I(N__29402));
    Span4Mux_h I__5274 (
            .O(N__29406),
            .I(N__29399));
    InMux I__5273 (
            .O(N__29405),
            .I(N__29396));
    Span4Mux_h I__5272 (
            .O(N__29402),
            .I(N__29393));
    Odrv4 I__5271 (
            .O(N__29399),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    LocalMux I__5270 (
            .O(N__29396),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    Odrv4 I__5269 (
            .O(N__29393),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    InMux I__5268 (
            .O(N__29386),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__5267 (
            .O(N__29383),
            .I(N__29380));
    LocalMux I__5266 (
            .O(N__29380),
            .I(N__29376));
    InMux I__5265 (
            .O(N__29379),
            .I(N__29373));
    Span4Mux_h I__5264 (
            .O(N__29376),
            .I(N__29369));
    LocalMux I__5263 (
            .O(N__29373),
            .I(N__29366));
    InMux I__5262 (
            .O(N__29372),
            .I(N__29363));
    Odrv4 I__5261 (
            .O(N__29369),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    Odrv4 I__5260 (
            .O(N__29366),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    LocalMux I__5259 (
            .O(N__29363),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    InMux I__5258 (
            .O(N__29356),
            .I(bfn_12_8_0_));
    CascadeMux I__5257 (
            .O(N__29353),
            .I(N__29349));
    CascadeMux I__5256 (
            .O(N__29352),
            .I(N__29345));
    InMux I__5255 (
            .O(N__29349),
            .I(N__29342));
    InMux I__5254 (
            .O(N__29348),
            .I(N__29339));
    InMux I__5253 (
            .O(N__29345),
            .I(N__29336));
    LocalMux I__5252 (
            .O(N__29342),
            .I(N__29333));
    LocalMux I__5251 (
            .O(N__29339),
            .I(N__29330));
    LocalMux I__5250 (
            .O(N__29336),
            .I(N__29327));
    Span4Mux_h I__5249 (
            .O(N__29333),
            .I(N__29324));
    Span4Mux_v I__5248 (
            .O(N__29330),
            .I(N__29319));
    Span4Mux_h I__5247 (
            .O(N__29327),
            .I(N__29319));
    Odrv4 I__5246 (
            .O(N__29324),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    Odrv4 I__5245 (
            .O(N__29319),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    InMux I__5244 (
            .O(N__29314),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__5243 (
            .O(N__29311),
            .I(N__29308));
    LocalMux I__5242 (
            .O(N__29308),
            .I(N__29303));
    InMux I__5241 (
            .O(N__29307),
            .I(N__29300));
    CascadeMux I__5240 (
            .O(N__29306),
            .I(N__29297));
    Span4Mux_h I__5239 (
            .O(N__29303),
            .I(N__29294));
    LocalMux I__5238 (
            .O(N__29300),
            .I(N__29291));
    InMux I__5237 (
            .O(N__29297),
            .I(N__29288));
    Odrv4 I__5236 (
            .O(N__29294),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    Odrv4 I__5235 (
            .O(N__29291),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    LocalMux I__5234 (
            .O(N__29288),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    InMux I__5233 (
            .O(N__29281),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__5232 (
            .O(N__29278),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__5231 (
            .O(N__29275),
            .I(N__29272));
    LocalMux I__5230 (
            .O(N__29272),
            .I(N__29263));
    InMux I__5229 (
            .O(N__29271),
            .I(N__29260));
    InMux I__5228 (
            .O(N__29270),
            .I(N__29255));
    InMux I__5227 (
            .O(N__29269),
            .I(N__29255));
    InMux I__5226 (
            .O(N__29268),
            .I(N__29252));
    InMux I__5225 (
            .O(N__29267),
            .I(N__29247));
    InMux I__5224 (
            .O(N__29266),
            .I(N__29247));
    Span4Mux_v I__5223 (
            .O(N__29263),
            .I(N__29240));
    LocalMux I__5222 (
            .O(N__29260),
            .I(N__29240));
    LocalMux I__5221 (
            .O(N__29255),
            .I(N__29240));
    LocalMux I__5220 (
            .O(N__29252),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    LocalMux I__5219 (
            .O(N__29247),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    Odrv4 I__5218 (
            .O(N__29240),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    InMux I__5217 (
            .O(N__29233),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__5216 (
            .O(N__29230),
            .I(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_ ));
    InMux I__5215 (
            .O(N__29227),
            .I(N__29223));
    InMux I__5214 (
            .O(N__29226),
            .I(N__29220));
    LocalMux I__5213 (
            .O(N__29223),
            .I(N__29215));
    LocalMux I__5212 (
            .O(N__29220),
            .I(N__29215));
    Span4Mux_v I__5211 (
            .O(N__29215),
            .I(N__29212));
    Odrv4 I__5210 (
            .O(N__29212),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    InMux I__5209 (
            .O(N__29209),
            .I(N__29205));
    CascadeMux I__5208 (
            .O(N__29208),
            .I(N__29201));
    LocalMux I__5207 (
            .O(N__29205),
            .I(N__29198));
    InMux I__5206 (
            .O(N__29204),
            .I(N__29195));
    InMux I__5205 (
            .O(N__29201),
            .I(N__29192));
    Span4Mux_v I__5204 (
            .O(N__29198),
            .I(N__29187));
    LocalMux I__5203 (
            .O(N__29195),
            .I(N__29187));
    LocalMux I__5202 (
            .O(N__29192),
            .I(N__29182));
    Span4Mux_h I__5201 (
            .O(N__29187),
            .I(N__29182));
    Odrv4 I__5200 (
            .O(N__29182),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    InMux I__5199 (
            .O(N__29179),
            .I(N__29175));
    InMux I__5198 (
            .O(N__29178),
            .I(N__29172));
    LocalMux I__5197 (
            .O(N__29175),
            .I(N__29168));
    LocalMux I__5196 (
            .O(N__29172),
            .I(N__29165));
    InMux I__5195 (
            .O(N__29171),
            .I(N__29162));
    Span4Mux_h I__5194 (
            .O(N__29168),
            .I(N__29159));
    Odrv12 I__5193 (
            .O(N__29165),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    LocalMux I__5192 (
            .O(N__29162),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    Odrv4 I__5191 (
            .O(N__29159),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    InMux I__5190 (
            .O(N__29152),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__5189 (
            .O(N__29149),
            .I(N__29145));
    InMux I__5188 (
            .O(N__29148),
            .I(N__29141));
    InMux I__5187 (
            .O(N__29145),
            .I(N__29138));
    InMux I__5186 (
            .O(N__29144),
            .I(N__29135));
    LocalMux I__5185 (
            .O(N__29141),
            .I(N__29130));
    LocalMux I__5184 (
            .O(N__29138),
            .I(N__29130));
    LocalMux I__5183 (
            .O(N__29135),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    Odrv4 I__5182 (
            .O(N__29130),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    InMux I__5181 (
            .O(N__29125),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__5180 (
            .O(N__29122),
            .I(N__29118));
    CascadeMux I__5179 (
            .O(N__29121),
            .I(N__29114));
    LocalMux I__5178 (
            .O(N__29118),
            .I(N__29111));
    InMux I__5177 (
            .O(N__29117),
            .I(N__29106));
    InMux I__5176 (
            .O(N__29114),
            .I(N__29106));
    Span4Mux_h I__5175 (
            .O(N__29111),
            .I(N__29101));
    LocalMux I__5174 (
            .O(N__29106),
            .I(N__29101));
    Span4Mux_h I__5173 (
            .O(N__29101),
            .I(N__29097));
    InMux I__5172 (
            .O(N__29100),
            .I(N__29094));
    Odrv4 I__5171 (
            .O(N__29097),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    LocalMux I__5170 (
            .O(N__29094),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    InMux I__5169 (
            .O(N__29089),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__5168 (
            .O(N__29086),
            .I(N__29083));
    InMux I__5167 (
            .O(N__29083),
            .I(N__29080));
    LocalMux I__5166 (
            .O(N__29080),
            .I(N__29077));
    Odrv4 I__5165 (
            .O(N__29077),
            .I(\current_shift_inst.control_input_1_axb_22 ));
    InMux I__5164 (
            .O(N__29074),
            .I(N__29070));
    CascadeMux I__5163 (
            .O(N__29073),
            .I(N__29067));
    LocalMux I__5162 (
            .O(N__29070),
            .I(N__29064));
    InMux I__5161 (
            .O(N__29067),
            .I(N__29061));
    Span4Mux_h I__5160 (
            .O(N__29064),
            .I(N__29056));
    LocalMux I__5159 (
            .O(N__29061),
            .I(N__29056));
    Span4Mux_h I__5158 (
            .O(N__29056),
            .I(N__29053));
    Span4Mux_h I__5157 (
            .O(N__29053),
            .I(N__29050));
    Odrv4 I__5156 (
            .O(N__29050),
            .I(\current_shift_inst.control_inputZ0Z_22 ));
    InMux I__5155 (
            .O(N__29047),
            .I(\current_shift_inst.control_input_1_cry_21 ));
    CascadeMux I__5154 (
            .O(N__29044),
            .I(N__29041));
    InMux I__5153 (
            .O(N__29041),
            .I(N__29038));
    LocalMux I__5152 (
            .O(N__29038),
            .I(N__29035));
    Odrv4 I__5151 (
            .O(N__29035),
            .I(\current_shift_inst.control_input_1_axb_23 ));
    InMux I__5150 (
            .O(N__29032),
            .I(N__29028));
    CascadeMux I__5149 (
            .O(N__29031),
            .I(N__29025));
    LocalMux I__5148 (
            .O(N__29028),
            .I(N__29022));
    InMux I__5147 (
            .O(N__29025),
            .I(N__29019));
    Span4Mux_v I__5146 (
            .O(N__29022),
            .I(N__29016));
    LocalMux I__5145 (
            .O(N__29019),
            .I(N__29013));
    Span4Mux_h I__5144 (
            .O(N__29016),
            .I(N__29008));
    Span4Mux_v I__5143 (
            .O(N__29013),
            .I(N__29008));
    Odrv4 I__5142 (
            .O(N__29008),
            .I(\current_shift_inst.control_inputZ0Z_23 ));
    InMux I__5141 (
            .O(N__29005),
            .I(\current_shift_inst.control_input_1_cry_22 ));
    InMux I__5140 (
            .O(N__29002),
            .I(N__28999));
    LocalMux I__5139 (
            .O(N__28999),
            .I(\current_shift_inst.control_input_1_axb_24 ));
    InMux I__5138 (
            .O(N__28996),
            .I(N__28992));
    CascadeMux I__5137 (
            .O(N__28995),
            .I(N__28989));
    LocalMux I__5136 (
            .O(N__28992),
            .I(N__28986));
    InMux I__5135 (
            .O(N__28989),
            .I(N__28983));
    Span4Mux_h I__5134 (
            .O(N__28986),
            .I(N__28978));
    LocalMux I__5133 (
            .O(N__28983),
            .I(N__28978));
    Span4Mux_h I__5132 (
            .O(N__28978),
            .I(N__28975));
    Odrv4 I__5131 (
            .O(N__28975),
            .I(\current_shift_inst.control_inputZ0Z_24 ));
    InMux I__5130 (
            .O(N__28972),
            .I(bfn_11_23_0_));
    CEMux I__5129 (
            .O(N__28969),
            .I(N__28966));
    LocalMux I__5128 (
            .O(N__28966),
            .I(N__28960));
    CEMux I__5127 (
            .O(N__28965),
            .I(N__28957));
    CEMux I__5126 (
            .O(N__28964),
            .I(N__28954));
    CEMux I__5125 (
            .O(N__28963),
            .I(N__28951));
    Span4Mux_v I__5124 (
            .O(N__28960),
            .I(N__28945));
    LocalMux I__5123 (
            .O(N__28957),
            .I(N__28945));
    LocalMux I__5122 (
            .O(N__28954),
            .I(N__28942));
    LocalMux I__5121 (
            .O(N__28951),
            .I(N__28939));
    CEMux I__5120 (
            .O(N__28950),
            .I(N__28936));
    Span4Mux_v I__5119 (
            .O(N__28945),
            .I(N__28933));
    Span4Mux_v I__5118 (
            .O(N__28942),
            .I(N__28930));
    Span4Mux_v I__5117 (
            .O(N__28939),
            .I(N__28927));
    LocalMux I__5116 (
            .O(N__28936),
            .I(N__28924));
    Span4Mux_h I__5115 (
            .O(N__28933),
            .I(N__28921));
    Span4Mux_h I__5114 (
            .O(N__28930),
            .I(N__28918));
    Sp12to4 I__5113 (
            .O(N__28927),
            .I(N__28915));
    Span4Mux_v I__5112 (
            .O(N__28924),
            .I(N__28912));
    Span4Mux_h I__5111 (
            .O(N__28921),
            .I(N__28909));
    Span4Mux_h I__5110 (
            .O(N__28918),
            .I(N__28906));
    Span12Mux_h I__5109 (
            .O(N__28915),
            .I(N__28903));
    Span4Mux_v I__5108 (
            .O(N__28912),
            .I(N__28900));
    Span4Mux_v I__5107 (
            .O(N__28909),
            .I(N__28897));
    Span4Mux_v I__5106 (
            .O(N__28906),
            .I(N__28894));
    Span12Mux_v I__5105 (
            .O(N__28903),
            .I(N__28889));
    Sp12to4 I__5104 (
            .O(N__28900),
            .I(N__28889));
    Odrv4 I__5103 (
            .O(N__28897),
            .I(\current_shift_inst.phase_valid_RNISLORZ0Z2 ));
    Odrv4 I__5102 (
            .O(N__28894),
            .I(\current_shift_inst.phase_valid_RNISLORZ0Z2 ));
    Odrv12 I__5101 (
            .O(N__28889),
            .I(\current_shift_inst.phase_valid_RNISLORZ0Z2 ));
    InMux I__5100 (
            .O(N__28882),
            .I(\current_shift_inst.control_input_1_cry_24 ));
    CascadeMux I__5099 (
            .O(N__28879),
            .I(N__28876));
    InMux I__5098 (
            .O(N__28876),
            .I(N__28873));
    LocalMux I__5097 (
            .O(N__28873),
            .I(N__28870));
    Odrv4 I__5096 (
            .O(N__28870),
            .I(\current_shift_inst.control_input_1_cry_24_THRU_CO ));
    InMux I__5095 (
            .O(N__28867),
            .I(N__28863));
    CascadeMux I__5094 (
            .O(N__28866),
            .I(N__28860));
    LocalMux I__5093 (
            .O(N__28863),
            .I(N__28857));
    InMux I__5092 (
            .O(N__28860),
            .I(N__28854));
    Span4Mux_h I__5091 (
            .O(N__28857),
            .I(N__28849));
    LocalMux I__5090 (
            .O(N__28854),
            .I(N__28849));
    Span4Mux_v I__5089 (
            .O(N__28849),
            .I(N__28846));
    Odrv4 I__5088 (
            .O(N__28846),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ));
    InMux I__5087 (
            .O(N__28843),
            .I(N__28840));
    LocalMux I__5086 (
            .O(N__28840),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ));
    InMux I__5085 (
            .O(N__28837),
            .I(N__28834));
    LocalMux I__5084 (
            .O(N__28834),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ));
    CascadeMux I__5083 (
            .O(N__28831),
            .I(N__28828));
    InMux I__5082 (
            .O(N__28828),
            .I(N__28825));
    LocalMux I__5081 (
            .O(N__28825),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ));
    CascadeMux I__5080 (
            .O(N__28822),
            .I(N__28819));
    InMux I__5079 (
            .O(N__28819),
            .I(N__28816));
    LocalMux I__5078 (
            .O(N__28816),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ));
    CascadeMux I__5077 (
            .O(N__28813),
            .I(N__28810));
    InMux I__5076 (
            .O(N__28810),
            .I(N__28807));
    LocalMux I__5075 (
            .O(N__28807),
            .I(N__28804));
    Odrv4 I__5074 (
            .O(N__28804),
            .I(\current_shift_inst.control_input_1_axb_14 ));
    InMux I__5073 (
            .O(N__28801),
            .I(N__28797));
    CascadeMux I__5072 (
            .O(N__28800),
            .I(N__28794));
    LocalMux I__5071 (
            .O(N__28797),
            .I(N__28791));
    InMux I__5070 (
            .O(N__28794),
            .I(N__28788));
    Span4Mux_h I__5069 (
            .O(N__28791),
            .I(N__28783));
    LocalMux I__5068 (
            .O(N__28788),
            .I(N__28783));
    Span4Mux_h I__5067 (
            .O(N__28783),
            .I(N__28780));
    Odrv4 I__5066 (
            .O(N__28780),
            .I(\current_shift_inst.control_inputZ0Z_14 ));
    InMux I__5065 (
            .O(N__28777),
            .I(\current_shift_inst.control_input_1_cry_13 ));
    CascadeMux I__5064 (
            .O(N__28774),
            .I(N__28771));
    InMux I__5063 (
            .O(N__28771),
            .I(N__28768));
    LocalMux I__5062 (
            .O(N__28768),
            .I(N__28765));
    Odrv4 I__5061 (
            .O(N__28765),
            .I(\current_shift_inst.control_input_1_axb_15 ));
    InMux I__5060 (
            .O(N__28762),
            .I(N__28758));
    CascadeMux I__5059 (
            .O(N__28761),
            .I(N__28755));
    LocalMux I__5058 (
            .O(N__28758),
            .I(N__28752));
    InMux I__5057 (
            .O(N__28755),
            .I(N__28749));
    Span4Mux_v I__5056 (
            .O(N__28752),
            .I(N__28746));
    LocalMux I__5055 (
            .O(N__28749),
            .I(N__28743));
    Sp12to4 I__5054 (
            .O(N__28746),
            .I(N__28740));
    Span4Mux_v I__5053 (
            .O(N__28743),
            .I(N__28737));
    Odrv12 I__5052 (
            .O(N__28740),
            .I(\current_shift_inst.control_inputZ0Z_15 ));
    Odrv4 I__5051 (
            .O(N__28737),
            .I(\current_shift_inst.control_inputZ0Z_15 ));
    InMux I__5050 (
            .O(N__28732),
            .I(\current_shift_inst.control_input_1_cry_14 ));
    InMux I__5049 (
            .O(N__28729),
            .I(N__28726));
    LocalMux I__5048 (
            .O(N__28726),
            .I(\current_shift_inst.control_input_1_axb_16 ));
    InMux I__5047 (
            .O(N__28723),
            .I(N__28719));
    CascadeMux I__5046 (
            .O(N__28722),
            .I(N__28716));
    LocalMux I__5045 (
            .O(N__28719),
            .I(N__28713));
    InMux I__5044 (
            .O(N__28716),
            .I(N__28710));
    Span4Mux_v I__5043 (
            .O(N__28713),
            .I(N__28707));
    LocalMux I__5042 (
            .O(N__28710),
            .I(N__28704));
    Span4Mux_h I__5041 (
            .O(N__28707),
            .I(N__28699));
    Span4Mux_v I__5040 (
            .O(N__28704),
            .I(N__28699));
    Odrv4 I__5039 (
            .O(N__28699),
            .I(\current_shift_inst.control_inputZ0Z_16 ));
    InMux I__5038 (
            .O(N__28696),
            .I(bfn_11_22_0_));
    InMux I__5037 (
            .O(N__28693),
            .I(N__28690));
    LocalMux I__5036 (
            .O(N__28690),
            .I(N__28687));
    Odrv4 I__5035 (
            .O(N__28687),
            .I(\current_shift_inst.control_input_1_axb_17 ));
    InMux I__5034 (
            .O(N__28684),
            .I(N__28680));
    InMux I__5033 (
            .O(N__28683),
            .I(N__28677));
    LocalMux I__5032 (
            .O(N__28680),
            .I(N__28674));
    LocalMux I__5031 (
            .O(N__28677),
            .I(N__28671));
    Span12Mux_s11_h I__5030 (
            .O(N__28674),
            .I(N__28668));
    Span4Mux_h I__5029 (
            .O(N__28671),
            .I(N__28665));
    Odrv12 I__5028 (
            .O(N__28668),
            .I(\current_shift_inst.control_inputZ0Z_17 ));
    Odrv4 I__5027 (
            .O(N__28665),
            .I(\current_shift_inst.control_inputZ0Z_17 ));
    InMux I__5026 (
            .O(N__28660),
            .I(\current_shift_inst.control_input_1_cry_16 ));
    InMux I__5025 (
            .O(N__28657),
            .I(N__28654));
    LocalMux I__5024 (
            .O(N__28654),
            .I(N__28651));
    Odrv4 I__5023 (
            .O(N__28651),
            .I(\current_shift_inst.control_input_1_axb_18 ));
    CascadeMux I__5022 (
            .O(N__28648),
            .I(N__28644));
    InMux I__5021 (
            .O(N__28647),
            .I(N__28641));
    InMux I__5020 (
            .O(N__28644),
            .I(N__28638));
    LocalMux I__5019 (
            .O(N__28641),
            .I(N__28635));
    LocalMux I__5018 (
            .O(N__28638),
            .I(N__28632));
    Span4Mux_h I__5017 (
            .O(N__28635),
            .I(N__28627));
    Span4Mux_v I__5016 (
            .O(N__28632),
            .I(N__28627));
    Odrv4 I__5015 (
            .O(N__28627),
            .I(\current_shift_inst.control_inputZ0Z_18 ));
    InMux I__5014 (
            .O(N__28624),
            .I(\current_shift_inst.control_input_1_cry_17 ));
    InMux I__5013 (
            .O(N__28621),
            .I(N__28618));
    LocalMux I__5012 (
            .O(N__28618),
            .I(N__28615));
    Odrv4 I__5011 (
            .O(N__28615),
            .I(\current_shift_inst.control_input_1_axb_19 ));
    InMux I__5010 (
            .O(N__28612),
            .I(N__28608));
    CascadeMux I__5009 (
            .O(N__28611),
            .I(N__28605));
    LocalMux I__5008 (
            .O(N__28608),
            .I(N__28602));
    InMux I__5007 (
            .O(N__28605),
            .I(N__28599));
    Span4Mux_h I__5006 (
            .O(N__28602),
            .I(N__28594));
    LocalMux I__5005 (
            .O(N__28599),
            .I(N__28594));
    Span4Mux_h I__5004 (
            .O(N__28594),
            .I(N__28591));
    Odrv4 I__5003 (
            .O(N__28591),
            .I(\current_shift_inst.control_inputZ0Z_19 ));
    InMux I__5002 (
            .O(N__28588),
            .I(\current_shift_inst.control_input_1_cry_18 ));
    CascadeMux I__5001 (
            .O(N__28585),
            .I(N__28582));
    InMux I__5000 (
            .O(N__28582),
            .I(N__28579));
    LocalMux I__4999 (
            .O(N__28579),
            .I(N__28576));
    Odrv4 I__4998 (
            .O(N__28576),
            .I(\current_shift_inst.control_input_1_axb_20 ));
    CascadeMux I__4997 (
            .O(N__28573),
            .I(N__28569));
    InMux I__4996 (
            .O(N__28572),
            .I(N__28566));
    InMux I__4995 (
            .O(N__28569),
            .I(N__28563));
    LocalMux I__4994 (
            .O(N__28566),
            .I(N__28558));
    LocalMux I__4993 (
            .O(N__28563),
            .I(N__28558));
    Span4Mux_v I__4992 (
            .O(N__28558),
            .I(N__28555));
    Odrv4 I__4991 (
            .O(N__28555),
            .I(\current_shift_inst.control_inputZ0Z_20 ));
    InMux I__4990 (
            .O(N__28552),
            .I(\current_shift_inst.control_input_1_cry_19 ));
    CascadeMux I__4989 (
            .O(N__28549),
            .I(N__28546));
    InMux I__4988 (
            .O(N__28546),
            .I(N__28543));
    LocalMux I__4987 (
            .O(N__28543),
            .I(N__28540));
    Odrv4 I__4986 (
            .O(N__28540),
            .I(\current_shift_inst.control_input_1_axb_21 ));
    InMux I__4985 (
            .O(N__28537),
            .I(N__28533));
    CascadeMux I__4984 (
            .O(N__28536),
            .I(N__28530));
    LocalMux I__4983 (
            .O(N__28533),
            .I(N__28527));
    InMux I__4982 (
            .O(N__28530),
            .I(N__28524));
    Span4Mux_v I__4981 (
            .O(N__28527),
            .I(N__28521));
    LocalMux I__4980 (
            .O(N__28524),
            .I(N__28518));
    Sp12to4 I__4979 (
            .O(N__28521),
            .I(N__28515));
    Span4Mux_v I__4978 (
            .O(N__28518),
            .I(N__28512));
    Odrv12 I__4977 (
            .O(N__28515),
            .I(\current_shift_inst.control_inputZ0Z_21 ));
    Odrv4 I__4976 (
            .O(N__28512),
            .I(\current_shift_inst.control_inputZ0Z_21 ));
    InMux I__4975 (
            .O(N__28507),
            .I(\current_shift_inst.control_input_1_cry_20 ));
    CascadeMux I__4974 (
            .O(N__28504),
            .I(N__28501));
    InMux I__4973 (
            .O(N__28501),
            .I(N__28498));
    LocalMux I__4972 (
            .O(N__28498),
            .I(N__28495));
    Odrv4 I__4971 (
            .O(N__28495),
            .I(\current_shift_inst.control_input_1_axb_6 ));
    CascadeMux I__4970 (
            .O(N__28492),
            .I(N__28489));
    InMux I__4969 (
            .O(N__28489),
            .I(N__28486));
    LocalMux I__4968 (
            .O(N__28486),
            .I(N__28482));
    InMux I__4967 (
            .O(N__28485),
            .I(N__28479));
    Span4Mux_h I__4966 (
            .O(N__28482),
            .I(N__28476));
    LocalMux I__4965 (
            .O(N__28479),
            .I(N__28473));
    Span4Mux_h I__4964 (
            .O(N__28476),
            .I(N__28470));
    Odrv12 I__4963 (
            .O(N__28473),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    Odrv4 I__4962 (
            .O(N__28470),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    InMux I__4961 (
            .O(N__28465),
            .I(\current_shift_inst.control_input_1_cry_5 ));
    CascadeMux I__4960 (
            .O(N__28462),
            .I(N__28459));
    InMux I__4959 (
            .O(N__28459),
            .I(N__28456));
    LocalMux I__4958 (
            .O(N__28456),
            .I(N__28453));
    Odrv4 I__4957 (
            .O(N__28453),
            .I(\current_shift_inst.control_input_1_axb_7 ));
    InMux I__4956 (
            .O(N__28450),
            .I(N__28446));
    CascadeMux I__4955 (
            .O(N__28449),
            .I(N__28443));
    LocalMux I__4954 (
            .O(N__28446),
            .I(N__28440));
    InMux I__4953 (
            .O(N__28443),
            .I(N__28437));
    Span4Mux_h I__4952 (
            .O(N__28440),
            .I(N__28434));
    LocalMux I__4951 (
            .O(N__28437),
            .I(N__28431));
    Span4Mux_h I__4950 (
            .O(N__28434),
            .I(N__28428));
    Span4Mux_v I__4949 (
            .O(N__28431),
            .I(N__28425));
    Odrv4 I__4948 (
            .O(N__28428),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    Odrv4 I__4947 (
            .O(N__28425),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    InMux I__4946 (
            .O(N__28420),
            .I(\current_shift_inst.control_input_1_cry_6 ));
    CascadeMux I__4945 (
            .O(N__28417),
            .I(N__28414));
    InMux I__4944 (
            .O(N__28414),
            .I(N__28411));
    LocalMux I__4943 (
            .O(N__28411),
            .I(\current_shift_inst.control_input_1_axb_8 ));
    CascadeMux I__4942 (
            .O(N__28408),
            .I(N__28404));
    InMux I__4941 (
            .O(N__28407),
            .I(N__28401));
    InMux I__4940 (
            .O(N__28404),
            .I(N__28398));
    LocalMux I__4939 (
            .O(N__28401),
            .I(N__28395));
    LocalMux I__4938 (
            .O(N__28398),
            .I(N__28392));
    Span12Mux_v I__4937 (
            .O(N__28395),
            .I(N__28389));
    Span4Mux_v I__4936 (
            .O(N__28392),
            .I(N__28386));
    Odrv12 I__4935 (
            .O(N__28389),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    Odrv4 I__4934 (
            .O(N__28386),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    InMux I__4933 (
            .O(N__28381),
            .I(bfn_11_21_0_));
    InMux I__4932 (
            .O(N__28378),
            .I(N__28375));
    LocalMux I__4931 (
            .O(N__28375),
            .I(N__28372));
    Odrv4 I__4930 (
            .O(N__28372),
            .I(\current_shift_inst.control_input_1_axb_9 ));
    InMux I__4929 (
            .O(N__28369),
            .I(N__28365));
    CascadeMux I__4928 (
            .O(N__28368),
            .I(N__28362));
    LocalMux I__4927 (
            .O(N__28365),
            .I(N__28359));
    InMux I__4926 (
            .O(N__28362),
            .I(N__28356));
    Span4Mux_h I__4925 (
            .O(N__28359),
            .I(N__28351));
    LocalMux I__4924 (
            .O(N__28356),
            .I(N__28351));
    Span4Mux_h I__4923 (
            .O(N__28351),
            .I(N__28348));
    Odrv4 I__4922 (
            .O(N__28348),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    InMux I__4921 (
            .O(N__28345),
            .I(\current_shift_inst.control_input_1_cry_8 ));
    InMux I__4920 (
            .O(N__28342),
            .I(N__28339));
    LocalMux I__4919 (
            .O(N__28339),
            .I(N__28336));
    Odrv4 I__4918 (
            .O(N__28336),
            .I(\current_shift_inst.control_input_1_axb_10 ));
    CascadeMux I__4917 (
            .O(N__28333),
            .I(N__28329));
    InMux I__4916 (
            .O(N__28332),
            .I(N__28326));
    InMux I__4915 (
            .O(N__28329),
            .I(N__28323));
    LocalMux I__4914 (
            .O(N__28326),
            .I(N__28320));
    LocalMux I__4913 (
            .O(N__28323),
            .I(N__28317));
    Span12Mux_s11_h I__4912 (
            .O(N__28320),
            .I(N__28314));
    Span4Mux_h I__4911 (
            .O(N__28317),
            .I(N__28311));
    Odrv12 I__4910 (
            .O(N__28314),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    Odrv4 I__4909 (
            .O(N__28311),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    InMux I__4908 (
            .O(N__28306),
            .I(\current_shift_inst.control_input_1_cry_9 ));
    InMux I__4907 (
            .O(N__28303),
            .I(N__28300));
    LocalMux I__4906 (
            .O(N__28300),
            .I(N__28297));
    Odrv4 I__4905 (
            .O(N__28297),
            .I(\current_shift_inst.control_input_1_axb_11 ));
    CascadeMux I__4904 (
            .O(N__28294),
            .I(N__28290));
    InMux I__4903 (
            .O(N__28293),
            .I(N__28287));
    InMux I__4902 (
            .O(N__28290),
            .I(N__28284));
    LocalMux I__4901 (
            .O(N__28287),
            .I(N__28281));
    LocalMux I__4900 (
            .O(N__28284),
            .I(N__28278));
    Span12Mux_s11_h I__4899 (
            .O(N__28281),
            .I(N__28275));
    Span4Mux_v I__4898 (
            .O(N__28278),
            .I(N__28272));
    Odrv12 I__4897 (
            .O(N__28275),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    Odrv4 I__4896 (
            .O(N__28272),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    InMux I__4895 (
            .O(N__28267),
            .I(\current_shift_inst.control_input_1_cry_10 ));
    InMux I__4894 (
            .O(N__28264),
            .I(N__28261));
    LocalMux I__4893 (
            .O(N__28261),
            .I(N__28258));
    Odrv4 I__4892 (
            .O(N__28258),
            .I(\current_shift_inst.control_input_1_axb_12 ));
    CascadeMux I__4891 (
            .O(N__28255),
            .I(N__28251));
    InMux I__4890 (
            .O(N__28254),
            .I(N__28248));
    InMux I__4889 (
            .O(N__28251),
            .I(N__28245));
    LocalMux I__4888 (
            .O(N__28248),
            .I(N__28240));
    LocalMux I__4887 (
            .O(N__28245),
            .I(N__28240));
    Span4Mux_v I__4886 (
            .O(N__28240),
            .I(N__28237));
    Odrv4 I__4885 (
            .O(N__28237),
            .I(\current_shift_inst.control_inputZ0Z_12 ));
    InMux I__4884 (
            .O(N__28234),
            .I(\current_shift_inst.control_input_1_cry_11 ));
    CascadeMux I__4883 (
            .O(N__28231),
            .I(N__28228));
    InMux I__4882 (
            .O(N__28228),
            .I(N__28225));
    LocalMux I__4881 (
            .O(N__28225),
            .I(N__28222));
    Odrv4 I__4880 (
            .O(N__28222),
            .I(\current_shift_inst.control_input_1_axb_13 ));
    CascadeMux I__4879 (
            .O(N__28219),
            .I(N__28216));
    InMux I__4878 (
            .O(N__28216),
            .I(N__28213));
    LocalMux I__4877 (
            .O(N__28213),
            .I(N__28209));
    InMux I__4876 (
            .O(N__28212),
            .I(N__28206));
    Span4Mux_v I__4875 (
            .O(N__28209),
            .I(N__28203));
    LocalMux I__4874 (
            .O(N__28206),
            .I(N__28200));
    Span4Mux_h I__4873 (
            .O(N__28203),
            .I(N__28197));
    Odrv12 I__4872 (
            .O(N__28200),
            .I(\current_shift_inst.control_inputZ0Z_13 ));
    Odrv4 I__4871 (
            .O(N__28197),
            .I(\current_shift_inst.control_inputZ0Z_13 ));
    InMux I__4870 (
            .O(N__28192),
            .I(\current_shift_inst.control_input_1_cry_12 ));
    InMux I__4869 (
            .O(N__28189),
            .I(N__28186));
    LocalMux I__4868 (
            .O(N__28186),
            .I(\current_shift_inst.control_input_1_axb_0 ));
    InMux I__4867 (
            .O(N__28183),
            .I(N__28180));
    LocalMux I__4866 (
            .O(N__28180),
            .I(N__28176));
    CascadeMux I__4865 (
            .O(N__28179),
            .I(N__28173));
    Span4Mux_v I__4864 (
            .O(N__28176),
            .I(N__28170));
    InMux I__4863 (
            .O(N__28173),
            .I(N__28167));
    Span4Mux_h I__4862 (
            .O(N__28170),
            .I(N__28162));
    LocalMux I__4861 (
            .O(N__28167),
            .I(N__28162));
    Span4Mux_v I__4860 (
            .O(N__28162),
            .I(N__28159));
    Odrv4 I__4859 (
            .O(N__28159),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    InMux I__4858 (
            .O(N__28156),
            .I(N__28153));
    LocalMux I__4857 (
            .O(N__28153),
            .I(N__28150));
    Odrv4 I__4856 (
            .O(N__28150),
            .I(\current_shift_inst.control_input_1_axb_1 ));
    InMux I__4855 (
            .O(N__28147),
            .I(N__28143));
    CascadeMux I__4854 (
            .O(N__28146),
            .I(N__28140));
    LocalMux I__4853 (
            .O(N__28143),
            .I(N__28137));
    InMux I__4852 (
            .O(N__28140),
            .I(N__28134));
    Span4Mux_h I__4851 (
            .O(N__28137),
            .I(N__28131));
    LocalMux I__4850 (
            .O(N__28134),
            .I(N__28128));
    Span4Mux_h I__4849 (
            .O(N__28131),
            .I(N__28125));
    Span4Mux_h I__4848 (
            .O(N__28128),
            .I(N__28122));
    Odrv4 I__4847 (
            .O(N__28125),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    Odrv4 I__4846 (
            .O(N__28122),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    InMux I__4845 (
            .O(N__28117),
            .I(\current_shift_inst.control_input_1_cry_0 ));
    InMux I__4844 (
            .O(N__28114),
            .I(N__28111));
    LocalMux I__4843 (
            .O(N__28111),
            .I(N__28108));
    Odrv4 I__4842 (
            .O(N__28108),
            .I(\current_shift_inst.control_input_1_axb_2 ));
    InMux I__4841 (
            .O(N__28105),
            .I(N__28102));
    LocalMux I__4840 (
            .O(N__28102),
            .I(N__28098));
    CascadeMux I__4839 (
            .O(N__28101),
            .I(N__28095));
    Span4Mux_s3_h I__4838 (
            .O(N__28098),
            .I(N__28092));
    InMux I__4837 (
            .O(N__28095),
            .I(N__28089));
    Span4Mux_h I__4836 (
            .O(N__28092),
            .I(N__28086));
    LocalMux I__4835 (
            .O(N__28089),
            .I(N__28083));
    Span4Mux_h I__4834 (
            .O(N__28086),
            .I(N__28080));
    Span4Mux_v I__4833 (
            .O(N__28083),
            .I(N__28077));
    Odrv4 I__4832 (
            .O(N__28080),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    Odrv4 I__4831 (
            .O(N__28077),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    InMux I__4830 (
            .O(N__28072),
            .I(\current_shift_inst.control_input_1_cry_1 ));
    InMux I__4829 (
            .O(N__28069),
            .I(N__28066));
    LocalMux I__4828 (
            .O(N__28066),
            .I(N__28063));
    Odrv4 I__4827 (
            .O(N__28063),
            .I(\current_shift_inst.control_input_1_axb_3 ));
    InMux I__4826 (
            .O(N__28060),
            .I(N__28057));
    LocalMux I__4825 (
            .O(N__28057),
            .I(N__28053));
    CascadeMux I__4824 (
            .O(N__28056),
            .I(N__28050));
    Span4Mux_h I__4823 (
            .O(N__28053),
            .I(N__28047));
    InMux I__4822 (
            .O(N__28050),
            .I(N__28044));
    Span4Mux_h I__4821 (
            .O(N__28047),
            .I(N__28041));
    LocalMux I__4820 (
            .O(N__28044),
            .I(N__28038));
    Sp12to4 I__4819 (
            .O(N__28041),
            .I(N__28035));
    Span4Mux_v I__4818 (
            .O(N__28038),
            .I(N__28032));
    Odrv12 I__4817 (
            .O(N__28035),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    Odrv4 I__4816 (
            .O(N__28032),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    InMux I__4815 (
            .O(N__28027),
            .I(\current_shift_inst.control_input_1_cry_2 ));
    CascadeMux I__4814 (
            .O(N__28024),
            .I(N__28021));
    InMux I__4813 (
            .O(N__28021),
            .I(N__28018));
    LocalMux I__4812 (
            .O(N__28018),
            .I(N__28015));
    Odrv4 I__4811 (
            .O(N__28015),
            .I(\current_shift_inst.control_input_1_axb_4 ));
    InMux I__4810 (
            .O(N__28012),
            .I(N__28008));
    CascadeMux I__4809 (
            .O(N__28011),
            .I(N__28005));
    LocalMux I__4808 (
            .O(N__28008),
            .I(N__28002));
    InMux I__4807 (
            .O(N__28005),
            .I(N__27999));
    Span4Mux_h I__4806 (
            .O(N__28002),
            .I(N__27996));
    LocalMux I__4805 (
            .O(N__27999),
            .I(N__27993));
    Span4Mux_h I__4804 (
            .O(N__27996),
            .I(N__27990));
    Span4Mux_v I__4803 (
            .O(N__27993),
            .I(N__27987));
    Odrv4 I__4802 (
            .O(N__27990),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    Odrv4 I__4801 (
            .O(N__27987),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    InMux I__4800 (
            .O(N__27982),
            .I(\current_shift_inst.control_input_1_cry_3 ));
    CascadeMux I__4799 (
            .O(N__27979),
            .I(N__27976));
    InMux I__4798 (
            .O(N__27976),
            .I(N__27973));
    LocalMux I__4797 (
            .O(N__27973),
            .I(N__27970));
    Odrv4 I__4796 (
            .O(N__27970),
            .I(\current_shift_inst.control_input_1_axb_5 ));
    InMux I__4795 (
            .O(N__27967),
            .I(N__27964));
    LocalMux I__4794 (
            .O(N__27964),
            .I(N__27960));
    CascadeMux I__4793 (
            .O(N__27963),
            .I(N__27957));
    Span4Mux_h I__4792 (
            .O(N__27960),
            .I(N__27954));
    InMux I__4791 (
            .O(N__27957),
            .I(N__27951));
    Span4Mux_v I__4790 (
            .O(N__27954),
            .I(N__27946));
    LocalMux I__4789 (
            .O(N__27951),
            .I(N__27946));
    Span4Mux_v I__4788 (
            .O(N__27946),
            .I(N__27943));
    Odrv4 I__4787 (
            .O(N__27943),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    InMux I__4786 (
            .O(N__27940),
            .I(\current_shift_inst.control_input_1_cry_4 ));
    InMux I__4785 (
            .O(N__27937),
            .I(N__27931));
    InMux I__4784 (
            .O(N__27936),
            .I(N__27931));
    LocalMux I__4783 (
            .O(N__27931),
            .I(N__27924));
    InMux I__4782 (
            .O(N__27930),
            .I(N__27921));
    InMux I__4781 (
            .O(N__27929),
            .I(N__27916));
    InMux I__4780 (
            .O(N__27928),
            .I(N__27916));
    InMux I__4779 (
            .O(N__27927),
            .I(N__27912));
    Span4Mux_v I__4778 (
            .O(N__27924),
            .I(N__27909));
    LocalMux I__4777 (
            .O(N__27921),
            .I(N__27906));
    LocalMux I__4776 (
            .O(N__27916),
            .I(N__27903));
    InMux I__4775 (
            .O(N__27915),
            .I(N__27900));
    LocalMux I__4774 (
            .O(N__27912),
            .I(N__27897));
    Span4Mux_h I__4773 (
            .O(N__27909),
            .I(N__27894));
    Span4Mux_v I__4772 (
            .O(N__27906),
            .I(N__27891));
    Span4Mux_h I__4771 (
            .O(N__27903),
            .I(N__27888));
    LocalMux I__4770 (
            .O(N__27900),
            .I(N__27885));
    Span4Mux_h I__4769 (
            .O(N__27897),
            .I(N__27882));
    Span4Mux_v I__4768 (
            .O(N__27894),
            .I(N__27879));
    Span4Mux_v I__4767 (
            .O(N__27891),
            .I(N__27876));
    Span4Mux_v I__4766 (
            .O(N__27888),
            .I(N__27873));
    Span4Mux_h I__4765 (
            .O(N__27885),
            .I(N__27868));
    Span4Mux_v I__4764 (
            .O(N__27882),
            .I(N__27868));
    Odrv4 I__4763 (
            .O(N__27879),
            .I(\current_shift_inst.S1_riseZ0 ));
    Odrv4 I__4762 (
            .O(N__27876),
            .I(\current_shift_inst.S1_riseZ0 ));
    Odrv4 I__4761 (
            .O(N__27873),
            .I(\current_shift_inst.S1_riseZ0 ));
    Odrv4 I__4760 (
            .O(N__27868),
            .I(\current_shift_inst.S1_riseZ0 ));
    InMux I__4759 (
            .O(N__27859),
            .I(N__27856));
    LocalMux I__4758 (
            .O(N__27856),
            .I(\current_shift_inst.S1_syncZ0Z0 ));
    InMux I__4757 (
            .O(N__27853),
            .I(N__27850));
    LocalMux I__4756 (
            .O(N__27850),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    InMux I__4755 (
            .O(N__27847),
            .I(N__27841));
    InMux I__4754 (
            .O(N__27846),
            .I(N__27841));
    LocalMux I__4753 (
            .O(N__27841),
            .I(\current_shift_inst.S1_syncZ0Z1 ));
    InMux I__4752 (
            .O(N__27838),
            .I(N__27835));
    LocalMux I__4751 (
            .O(N__27835),
            .I(\current_shift_inst.S1_sync_prevZ0 ));
    CascadeMux I__4750 (
            .O(N__27832),
            .I(N__27829));
    InMux I__4749 (
            .O(N__27829),
            .I(N__27826));
    LocalMux I__4748 (
            .O(N__27826),
            .I(N__27823));
    Span4Mux_v I__4747 (
            .O(N__27823),
            .I(N__27820));
    Odrv4 I__4746 (
            .O(N__27820),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ));
    InMux I__4745 (
            .O(N__27817),
            .I(N__27814));
    LocalMux I__4744 (
            .O(N__27814),
            .I(N__27811));
    Span4Mux_v I__4743 (
            .O(N__27811),
            .I(N__27808));
    Sp12to4 I__4742 (
            .O(N__27808),
            .I(N__27805));
    Odrv12 I__4741 (
            .O(N__27805),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ));
    CascadeMux I__4740 (
            .O(N__27802),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ));
    InMux I__4739 (
            .O(N__27799),
            .I(N__27796));
    LocalMux I__4738 (
            .O(N__27796),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10 ));
    InMux I__4737 (
            .O(N__27793),
            .I(N__27788));
    InMux I__4736 (
            .O(N__27792),
            .I(N__27785));
    InMux I__4735 (
            .O(N__27791),
            .I(N__27782));
    LocalMux I__4734 (
            .O(N__27788),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__4733 (
            .O(N__27785),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__4732 (
            .O(N__27782),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__4731 (
            .O(N__27775),
            .I(N__27770));
    InMux I__4730 (
            .O(N__27774),
            .I(N__27767));
    InMux I__4729 (
            .O(N__27773),
            .I(N__27764));
    LocalMux I__4728 (
            .O(N__27770),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__4727 (
            .O(N__27767),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__4726 (
            .O(N__27764),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__4725 (
            .O(N__27757),
            .I(N__27752));
    InMux I__4724 (
            .O(N__27756),
            .I(N__27749));
    InMux I__4723 (
            .O(N__27755),
            .I(N__27746));
    LocalMux I__4722 (
            .O(N__27752),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__4721 (
            .O(N__27749),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__4720 (
            .O(N__27746),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__4719 (
            .O(N__27739),
            .I(N__27734));
    InMux I__4718 (
            .O(N__27738),
            .I(N__27731));
    InMux I__4717 (
            .O(N__27737),
            .I(N__27728));
    LocalMux I__4716 (
            .O(N__27734),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__4715 (
            .O(N__27731),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__4714 (
            .O(N__27728),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__4713 (
            .O(N__27721),
            .I(N__27716));
    InMux I__4712 (
            .O(N__27720),
            .I(N__27713));
    InMux I__4711 (
            .O(N__27719),
            .I(N__27710));
    LocalMux I__4710 (
            .O(N__27716),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__4709 (
            .O(N__27713),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__4708 (
            .O(N__27710),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    CascadeMux I__4707 (
            .O(N__27703),
            .I(\pwm_generator_inst.un1_counterlto9_2_cascade_ ));
    InMux I__4706 (
            .O(N__27700),
            .I(N__27682));
    InMux I__4705 (
            .O(N__27699),
            .I(N__27682));
    InMux I__4704 (
            .O(N__27698),
            .I(N__27682));
    InMux I__4703 (
            .O(N__27697),
            .I(N__27682));
    InMux I__4702 (
            .O(N__27696),
            .I(N__27677));
    InMux I__4701 (
            .O(N__27695),
            .I(N__27677));
    InMux I__4700 (
            .O(N__27694),
            .I(N__27668));
    InMux I__4699 (
            .O(N__27693),
            .I(N__27668));
    InMux I__4698 (
            .O(N__27692),
            .I(N__27668));
    InMux I__4697 (
            .O(N__27691),
            .I(N__27668));
    LocalMux I__4696 (
            .O(N__27682),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__4695 (
            .O(N__27677),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__4694 (
            .O(N__27668),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__4693 (
            .O(N__27661),
            .I(N__27656));
    InMux I__4692 (
            .O(N__27660),
            .I(N__27653));
    InMux I__4691 (
            .O(N__27659),
            .I(N__27650));
    LocalMux I__4690 (
            .O(N__27656),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__4689 (
            .O(N__27653),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__4688 (
            .O(N__27650),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__4687 (
            .O(N__27643),
            .I(N__27638));
    InMux I__4686 (
            .O(N__27642),
            .I(N__27635));
    InMux I__4685 (
            .O(N__27641),
            .I(N__27632));
    LocalMux I__4684 (
            .O(N__27638),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__4683 (
            .O(N__27635),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__4682 (
            .O(N__27632),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__4681 (
            .O(N__27625),
            .I(N__27620));
    InMux I__4680 (
            .O(N__27624),
            .I(N__27617));
    InMux I__4679 (
            .O(N__27623),
            .I(N__27614));
    LocalMux I__4678 (
            .O(N__27620),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__4677 (
            .O(N__27617),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__4676 (
            .O(N__27614),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__4675 (
            .O(N__27607),
            .I(N__27602));
    InMux I__4674 (
            .O(N__27606),
            .I(N__27599));
    InMux I__4673 (
            .O(N__27605),
            .I(N__27596));
    LocalMux I__4672 (
            .O(N__27602),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__4671 (
            .O(N__27599),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__4670 (
            .O(N__27596),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    CascadeMux I__4669 (
            .O(N__27589),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__4668 (
            .O(N__27586),
            .I(N__27581));
    InMux I__4667 (
            .O(N__27585),
            .I(N__27578));
    InMux I__4666 (
            .O(N__27584),
            .I(N__27575));
    LocalMux I__4665 (
            .O(N__27581),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__4664 (
            .O(N__27578),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__4663 (
            .O(N__27575),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__4662 (
            .O(N__27568),
            .I(N__27565));
    LocalMux I__4661 (
            .O(N__27565),
            .I(\pwm_generator_inst.un1_counterlt9 ));
    InMux I__4660 (
            .O(N__27562),
            .I(N__27559));
    LocalMux I__4659 (
            .O(N__27559),
            .I(N__27556));
    Odrv12 I__4658 (
            .O(N__27556),
            .I(il_min_comp1_D1));
    InMux I__4657 (
            .O(N__27553),
            .I(N__27549));
    InMux I__4656 (
            .O(N__27552),
            .I(N__27546));
    LocalMux I__4655 (
            .O(N__27549),
            .I(N__27543));
    LocalMux I__4654 (
            .O(N__27546),
            .I(N__27540));
    Span4Mux_h I__4653 (
            .O(N__27543),
            .I(N__27537));
    Odrv4 I__4652 (
            .O(N__27540),
            .I(\phase_controller_inst1.N_231 ));
    Odrv4 I__4651 (
            .O(N__27537),
            .I(\phase_controller_inst1.N_231 ));
    InMux I__4650 (
            .O(N__27532),
            .I(N__27529));
    LocalMux I__4649 (
            .O(N__27529),
            .I(N__27523));
    InMux I__4648 (
            .O(N__27528),
            .I(N__27520));
    InMux I__4647 (
            .O(N__27527),
            .I(N__27517));
    InMux I__4646 (
            .O(N__27526),
            .I(N__27514));
    Odrv4 I__4645 (
            .O(N__27523),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__4644 (
            .O(N__27520),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__4643 (
            .O(N__27517),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__4642 (
            .O(N__27514),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    InMux I__4641 (
            .O(N__27505),
            .I(N__27502));
    LocalMux I__4640 (
            .O(N__27502),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2 ));
    InMux I__4639 (
            .O(N__27499),
            .I(N__27496));
    LocalMux I__4638 (
            .O(N__27496),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ));
    CascadeMux I__4637 (
            .O(N__27493),
            .I(N__27490));
    InMux I__4636 (
            .O(N__27490),
            .I(N__27487));
    LocalMux I__4635 (
            .O(N__27487),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1 ));
    CascadeMux I__4634 (
            .O(N__27484),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_ ));
    InMux I__4633 (
            .O(N__27481),
            .I(N__27478));
    LocalMux I__4632 (
            .O(N__27478),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0 ));
    InMux I__4631 (
            .O(N__27475),
            .I(N__27472));
    LocalMux I__4630 (
            .O(N__27472),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ));
    InMux I__4629 (
            .O(N__27469),
            .I(N__27463));
    InMux I__4628 (
            .O(N__27468),
            .I(N__27463));
    LocalMux I__4627 (
            .O(N__27463),
            .I(N__27460));
    Odrv4 I__4626 (
            .O(N__27460),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ));
    InMux I__4625 (
            .O(N__27457),
            .I(N__27454));
    LocalMux I__4624 (
            .O(N__27454),
            .I(N__27449));
    InMux I__4623 (
            .O(N__27453),
            .I(N__27444));
    InMux I__4622 (
            .O(N__27452),
            .I(N__27444));
    Span4Mux_h I__4621 (
            .O(N__27449),
            .I(N__27441));
    LocalMux I__4620 (
            .O(N__27444),
            .I(N__27438));
    Odrv4 I__4619 (
            .O(N__27441),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ));
    Odrv4 I__4618 (
            .O(N__27438),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ));
    InMux I__4617 (
            .O(N__27433),
            .I(N__27430));
    LocalMux I__4616 (
            .O(N__27430),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ));
    InMux I__4615 (
            .O(N__27427),
            .I(N__27424));
    LocalMux I__4614 (
            .O(N__27424),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ));
    CascadeMux I__4613 (
            .O(N__27421),
            .I(N__27418));
    InMux I__4612 (
            .O(N__27418),
            .I(N__27415));
    LocalMux I__4611 (
            .O(N__27415),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ));
    CascadeMux I__4610 (
            .O(N__27412),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_ ));
    InMux I__4609 (
            .O(N__27409),
            .I(N__27406));
    LocalMux I__4608 (
            .O(N__27406),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ));
    InMux I__4607 (
            .O(N__27403),
            .I(N__27400));
    LocalMux I__4606 (
            .O(N__27400),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ));
    CascadeMux I__4605 (
            .O(N__27397),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_ ));
    InMux I__4604 (
            .O(N__27394),
            .I(N__27391));
    LocalMux I__4603 (
            .O(N__27391),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ));
    CascadeMux I__4602 (
            .O(N__27388),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ));
    InMux I__4601 (
            .O(N__27385),
            .I(N__27382));
    LocalMux I__4600 (
            .O(N__27382),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ));
    InMux I__4599 (
            .O(N__27379),
            .I(N__27373));
    InMux I__4598 (
            .O(N__27378),
            .I(N__27373));
    LocalMux I__4597 (
            .O(N__27373),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1 ));
    InMux I__4596 (
            .O(N__27370),
            .I(N__27367));
    LocalMux I__4595 (
            .O(N__27367),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14 ));
    InMux I__4594 (
            .O(N__27364),
            .I(N__27361));
    LocalMux I__4593 (
            .O(N__27361),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ));
    CascadeMux I__4592 (
            .O(N__27358),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0_cascade_ ));
    InMux I__4591 (
            .O(N__27355),
            .I(\current_shift_inst.un38_control_input_0_cry_28 ));
    InMux I__4590 (
            .O(N__27352),
            .I(\current_shift_inst.un38_control_input_0_cry_29 ));
    InMux I__4589 (
            .O(N__27349),
            .I(bfn_10_25_0_));
    CascadeMux I__4588 (
            .O(N__27346),
            .I(N__27338));
    CascadeMux I__4587 (
            .O(N__27345),
            .I(N__27334));
    CascadeMux I__4586 (
            .O(N__27344),
            .I(N__27330));
    InMux I__4585 (
            .O(N__27343),
            .I(N__27327));
    InMux I__4584 (
            .O(N__27342),
            .I(N__27312));
    InMux I__4583 (
            .O(N__27341),
            .I(N__27312));
    InMux I__4582 (
            .O(N__27338),
            .I(N__27312));
    InMux I__4581 (
            .O(N__27337),
            .I(N__27312));
    InMux I__4580 (
            .O(N__27334),
            .I(N__27312));
    InMux I__4579 (
            .O(N__27333),
            .I(N__27312));
    InMux I__4578 (
            .O(N__27330),
            .I(N__27312));
    LocalMux I__4577 (
            .O(N__27327),
            .I(N__27309));
    LocalMux I__4576 (
            .O(N__27312),
            .I(N__27306));
    Span4Mux_h I__4575 (
            .O(N__27309),
            .I(N__27303));
    Span4Mux_v I__4574 (
            .O(N__27306),
            .I(N__27300));
    Span4Mux_h I__4573 (
            .O(N__27303),
            .I(N__27297));
    Span4Mux_v I__4572 (
            .O(N__27300),
            .I(N__27294));
    Odrv4 I__4571 (
            .O(N__27297),
            .I(\current_shift_inst.control_inputZ0Z_25 ));
    Odrv4 I__4570 (
            .O(N__27294),
            .I(\current_shift_inst.control_inputZ0Z_25 ));
    InMux I__4569 (
            .O(N__27289),
            .I(N__27286));
    LocalMux I__4568 (
            .O(N__27286),
            .I(N__27283));
    Span4Mux_h I__4567 (
            .O(N__27283),
            .I(N__27280));
    Span4Mux_h I__4566 (
            .O(N__27280),
            .I(N__27277));
    Odrv4 I__4565 (
            .O(N__27277),
            .I(il_max_comp2_c));
    InMux I__4564 (
            .O(N__27274),
            .I(N__27269));
    InMux I__4563 (
            .O(N__27273),
            .I(N__27266));
    InMux I__4562 (
            .O(N__27272),
            .I(N__27263));
    LocalMux I__4561 (
            .O(N__27269),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    LocalMux I__4560 (
            .O(N__27266),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    LocalMux I__4559 (
            .O(N__27263),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    IoInMux I__4558 (
            .O(N__27256),
            .I(N__27253));
    LocalMux I__4557 (
            .O(N__27253),
            .I(N__27250));
    Span4Mux_s1_v I__4556 (
            .O(N__27250),
            .I(N__27247));
    Odrv4 I__4555 (
            .O(N__27247),
            .I(\delay_measurement_inst.delay_hc_timer.N_336_i ));
    InMux I__4554 (
            .O(N__27244),
            .I(N__27240));
    InMux I__4553 (
            .O(N__27243),
            .I(N__27237));
    LocalMux I__4552 (
            .O(N__27240),
            .I(measured_delay_hc_27));
    LocalMux I__4551 (
            .O(N__27237),
            .I(measured_delay_hc_27));
    InMux I__4550 (
            .O(N__27232),
            .I(N__27228));
    InMux I__4549 (
            .O(N__27231),
            .I(N__27225));
    LocalMux I__4548 (
            .O(N__27228),
            .I(measured_delay_hc_28));
    LocalMux I__4547 (
            .O(N__27225),
            .I(measured_delay_hc_28));
    InMux I__4546 (
            .O(N__27220),
            .I(N__27217));
    LocalMux I__4545 (
            .O(N__27217),
            .I(N__27214));
    Span12Mux_h I__4544 (
            .O(N__27214),
            .I(N__27211));
    Odrv12 I__4543 (
            .O(N__27211),
            .I(il_min_comp1_c));
    InMux I__4542 (
            .O(N__27208),
            .I(N__27205));
    LocalMux I__4541 (
            .O(N__27205),
            .I(N__27202));
    Odrv12 I__4540 (
            .O(N__27202),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ));
    CascadeMux I__4539 (
            .O(N__27199),
            .I(N__27196));
    InMux I__4538 (
            .O(N__27196),
            .I(N__27193));
    LocalMux I__4537 (
            .O(N__27193),
            .I(N__27190));
    Odrv12 I__4536 (
            .O(N__27190),
            .I(\current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ));
    InMux I__4535 (
            .O(N__27187),
            .I(\current_shift_inst.un38_control_input_0_cry_20 ));
    InMux I__4534 (
            .O(N__27184),
            .I(N__27181));
    LocalMux I__4533 (
            .O(N__27181),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ));
    CascadeMux I__4532 (
            .O(N__27178),
            .I(N__27175));
    InMux I__4531 (
            .O(N__27175),
            .I(N__27172));
    LocalMux I__4530 (
            .O(N__27172),
            .I(N__27169));
    Odrv12 I__4529 (
            .O(N__27169),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ));
    InMux I__4528 (
            .O(N__27166),
            .I(\current_shift_inst.un38_control_input_0_cry_21 ));
    InMux I__4527 (
            .O(N__27163),
            .I(N__27160));
    LocalMux I__4526 (
            .O(N__27160),
            .I(N__27157));
    Span4Mux_v I__4525 (
            .O(N__27157),
            .I(N__27154));
    Span4Mux_v I__4524 (
            .O(N__27154),
            .I(N__27151));
    Odrv4 I__4523 (
            .O(N__27151),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ));
    CascadeMux I__4522 (
            .O(N__27148),
            .I(N__27145));
    InMux I__4521 (
            .O(N__27145),
            .I(N__27142));
    LocalMux I__4520 (
            .O(N__27142),
            .I(N__27139));
    Span4Mux_v I__4519 (
            .O(N__27139),
            .I(N__27136));
    Span4Mux_v I__4518 (
            .O(N__27136),
            .I(N__27133));
    Odrv4 I__4517 (
            .O(N__27133),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ));
    InMux I__4516 (
            .O(N__27130),
            .I(bfn_10_24_0_));
    InMux I__4515 (
            .O(N__27127),
            .I(\current_shift_inst.un38_control_input_0_cry_23 ));
    InMux I__4514 (
            .O(N__27124),
            .I(\current_shift_inst.un38_control_input_0_cry_24 ));
    InMux I__4513 (
            .O(N__27121),
            .I(\current_shift_inst.un38_control_input_0_cry_25 ));
    InMux I__4512 (
            .O(N__27118),
            .I(\current_shift_inst.un38_control_input_0_cry_26 ));
    InMux I__4511 (
            .O(N__27115),
            .I(\current_shift_inst.un38_control_input_0_cry_27 ));
    CascadeMux I__4510 (
            .O(N__27112),
            .I(N__27109));
    InMux I__4509 (
            .O(N__27109),
            .I(N__27106));
    LocalMux I__4508 (
            .O(N__27106),
            .I(\current_shift_inst.elapsed_time_ns_1_RNILORI_11 ));
    InMux I__4507 (
            .O(N__27103),
            .I(\current_shift_inst.un38_control_input_0_cry_11 ));
    CascadeMux I__4506 (
            .O(N__27100),
            .I(N__27097));
    InMux I__4505 (
            .O(N__27097),
            .I(N__27094));
    LocalMux I__4504 (
            .O(N__27094),
            .I(N__27091));
    Odrv12 I__4503 (
            .O(N__27091),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ));
    InMux I__4502 (
            .O(N__27088),
            .I(\current_shift_inst.un38_control_input_0_cry_12 ));
    InMux I__4501 (
            .O(N__27085),
            .I(N__27082));
    LocalMux I__4500 (
            .O(N__27082),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ));
    CascadeMux I__4499 (
            .O(N__27079),
            .I(N__27076));
    InMux I__4498 (
            .O(N__27076),
            .I(N__27073));
    LocalMux I__4497 (
            .O(N__27073),
            .I(N__27070));
    Odrv12 I__4496 (
            .O(N__27070),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ));
    InMux I__4495 (
            .O(N__27067),
            .I(\current_shift_inst.un38_control_input_0_cry_13 ));
    CascadeMux I__4494 (
            .O(N__27064),
            .I(N__27061));
    InMux I__4493 (
            .O(N__27061),
            .I(N__27058));
    LocalMux I__4492 (
            .O(N__27058),
            .I(N__27055));
    Odrv12 I__4491 (
            .O(N__27055),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ));
    InMux I__4490 (
            .O(N__27052),
            .I(bfn_10_23_0_));
    InMux I__4489 (
            .O(N__27049),
            .I(N__27046));
    LocalMux I__4488 (
            .O(N__27046),
            .I(N__27043));
    Span4Mux_v I__4487 (
            .O(N__27043),
            .I(N__27040));
    Odrv4 I__4486 (
            .O(N__27040),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ));
    CascadeMux I__4485 (
            .O(N__27037),
            .I(N__27034));
    InMux I__4484 (
            .O(N__27034),
            .I(N__27031));
    LocalMux I__4483 (
            .O(N__27031),
            .I(N__27028));
    Odrv12 I__4482 (
            .O(N__27028),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI190J_15 ));
    InMux I__4481 (
            .O(N__27025),
            .I(\current_shift_inst.un38_control_input_0_cry_15 ));
    InMux I__4480 (
            .O(N__27022),
            .I(\current_shift_inst.un38_control_input_0_cry_16 ));
    InMux I__4479 (
            .O(N__27019),
            .I(N__27016));
    LocalMux I__4478 (
            .O(N__27016),
            .I(N__27013));
    Odrv12 I__4477 (
            .O(N__27013),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ));
    InMux I__4476 (
            .O(N__27010),
            .I(\current_shift_inst.un38_control_input_0_cry_17 ));
    InMux I__4475 (
            .O(N__27007),
            .I(N__27004));
    LocalMux I__4474 (
            .O(N__27004),
            .I(N__27001));
    Odrv12 I__4473 (
            .O(N__27001),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ));
    CascadeMux I__4472 (
            .O(N__26998),
            .I(N__26995));
    InMux I__4471 (
            .O(N__26995),
            .I(N__26992));
    LocalMux I__4470 (
            .O(N__26992),
            .I(N__26989));
    Span4Mux_v I__4469 (
            .O(N__26989),
            .I(N__26986));
    Odrv4 I__4468 (
            .O(N__26986),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ));
    InMux I__4467 (
            .O(N__26983),
            .I(\current_shift_inst.un38_control_input_0_cry_18 ));
    InMux I__4466 (
            .O(N__26980),
            .I(\current_shift_inst.un38_control_input_0_cry_19 ));
    InMux I__4465 (
            .O(N__26977),
            .I(N__26974));
    LocalMux I__4464 (
            .O(N__26974),
            .I(N__26971));
    Odrv4 I__4463 (
            .O(N__26971),
            .I(\current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ));
    InMux I__4462 (
            .O(N__26968),
            .I(N__26965));
    LocalMux I__4461 (
            .O(N__26965),
            .I(N__26962));
    Odrv12 I__4460 (
            .O(N__26962),
            .I(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ));
    CascadeMux I__4459 (
            .O(N__26959),
            .I(N__26956));
    InMux I__4458 (
            .O(N__26956),
            .I(N__26953));
    LocalMux I__4457 (
            .O(N__26953),
            .I(N__26950));
    Odrv4 I__4456 (
            .O(N__26950),
            .I(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ));
    CascadeMux I__4455 (
            .O(N__26947),
            .I(N__26944));
    InMux I__4454 (
            .O(N__26944),
            .I(N__26941));
    LocalMux I__4453 (
            .O(N__26941),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ));
    InMux I__4452 (
            .O(N__26938),
            .I(\current_shift_inst.un38_control_input_0_cry_5 ));
    InMux I__4451 (
            .O(N__26935),
            .I(N__26932));
    LocalMux I__4450 (
            .O(N__26932),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ));
    CascadeMux I__4449 (
            .O(N__26929),
            .I(N__26926));
    InMux I__4448 (
            .O(N__26926),
            .I(N__26923));
    LocalMux I__4447 (
            .O(N__26923),
            .I(N__26920));
    Odrv4 I__4446 (
            .O(N__26920),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ));
    InMux I__4445 (
            .O(N__26917),
            .I(bfn_10_22_0_));
    CascadeMux I__4444 (
            .O(N__26914),
            .I(N__26911));
    InMux I__4443 (
            .O(N__26911),
            .I(N__26908));
    LocalMux I__4442 (
            .O(N__26908),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ));
    InMux I__4441 (
            .O(N__26905),
            .I(\current_shift_inst.un38_control_input_0_cry_7 ));
    InMux I__4440 (
            .O(N__26902),
            .I(N__26899));
    LocalMux I__4439 (
            .O(N__26899),
            .I(N__26896));
    Odrv4 I__4438 (
            .O(N__26896),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ));
    InMux I__4437 (
            .O(N__26893),
            .I(\current_shift_inst.un38_control_input_0_cry_8 ));
    InMux I__4436 (
            .O(N__26890),
            .I(N__26887));
    LocalMux I__4435 (
            .O(N__26887),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ));
    CascadeMux I__4434 (
            .O(N__26884),
            .I(N__26881));
    InMux I__4433 (
            .O(N__26881),
            .I(N__26878));
    LocalMux I__4432 (
            .O(N__26878),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ));
    InMux I__4431 (
            .O(N__26875),
            .I(\current_shift_inst.un38_control_input_0_cry_9 ));
    CascadeMux I__4430 (
            .O(N__26872),
            .I(N__26869));
    InMux I__4429 (
            .O(N__26869),
            .I(N__26866));
    LocalMux I__4428 (
            .O(N__26866),
            .I(N__26863));
    Odrv12 I__4427 (
            .O(N__26863),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ));
    InMux I__4426 (
            .O(N__26860),
            .I(\current_shift_inst.un38_control_input_0_cry_10 ));
    InMux I__4425 (
            .O(N__26857),
            .I(N__26854));
    LocalMux I__4424 (
            .O(N__26854),
            .I(\current_shift_inst.z_i_0_31 ));
    CascadeMux I__4423 (
            .O(N__26851),
            .I(N__26848));
    InMux I__4422 (
            .O(N__26848),
            .I(N__26845));
    LocalMux I__4421 (
            .O(N__26845),
            .I(N__26842));
    Odrv4 I__4420 (
            .O(N__26842),
            .I(\current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ));
    CascadeMux I__4419 (
            .O(N__26839),
            .I(N__26836));
    InMux I__4418 (
            .O(N__26836),
            .I(N__26833));
    LocalMux I__4417 (
            .O(N__26833),
            .I(\current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ));
    CascadeMux I__4416 (
            .O(N__26830),
            .I(N__26827));
    InMux I__4415 (
            .O(N__26827),
            .I(N__26824));
    LocalMux I__4414 (
            .O(N__26824),
            .I(\current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ));
    InMux I__4413 (
            .O(N__26821),
            .I(N__26816));
    InMux I__4412 (
            .O(N__26820),
            .I(N__26813));
    InMux I__4411 (
            .O(N__26819),
            .I(N__26810));
    LocalMux I__4410 (
            .O(N__26816),
            .I(N__26806));
    LocalMux I__4409 (
            .O(N__26813),
            .I(N__26803));
    LocalMux I__4408 (
            .O(N__26810),
            .I(N__26800));
    InMux I__4407 (
            .O(N__26809),
            .I(N__26797));
    Span4Mux_v I__4406 (
            .O(N__26806),
            .I(N__26792));
    Span4Mux_v I__4405 (
            .O(N__26803),
            .I(N__26792));
    Odrv12 I__4404 (
            .O(N__26800),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__4403 (
            .O(N__26797),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__4402 (
            .O(N__26792),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    CascadeMux I__4401 (
            .O(N__26785),
            .I(N__26780));
    InMux I__4400 (
            .O(N__26784),
            .I(N__26777));
    InMux I__4399 (
            .O(N__26783),
            .I(N__26773));
    InMux I__4398 (
            .O(N__26780),
            .I(N__26770));
    LocalMux I__4397 (
            .O(N__26777),
            .I(N__26767));
    InMux I__4396 (
            .O(N__26776),
            .I(N__26764));
    LocalMux I__4395 (
            .O(N__26773),
            .I(N__26761));
    LocalMux I__4394 (
            .O(N__26770),
            .I(N__26758));
    Odrv4 I__4393 (
            .O(N__26767),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__4392 (
            .O(N__26764),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__4391 (
            .O(N__26761),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv12 I__4390 (
            .O(N__26758),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__4389 (
            .O(N__26749),
            .I(N__26746));
    InMux I__4388 (
            .O(N__26746),
            .I(N__26743));
    LocalMux I__4387 (
            .O(N__26743),
            .I(N__26739));
    InMux I__4386 (
            .O(N__26742),
            .I(N__26735));
    Span4Mux_v I__4385 (
            .O(N__26739),
            .I(N__26732));
    CascadeMux I__4384 (
            .O(N__26738),
            .I(N__26729));
    LocalMux I__4383 (
            .O(N__26735),
            .I(N__26725));
    Span4Mux_h I__4382 (
            .O(N__26732),
            .I(N__26722));
    InMux I__4381 (
            .O(N__26729),
            .I(N__26719));
    InMux I__4380 (
            .O(N__26728),
            .I(N__26716));
    Span4Mux_h I__4379 (
            .O(N__26725),
            .I(N__26713));
    Odrv4 I__4378 (
            .O(N__26722),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__4377 (
            .O(N__26719),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__4376 (
            .O(N__26716),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__4375 (
            .O(N__26713),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__4374 (
            .O(N__26704),
            .I(N__26701));
    LocalMux I__4373 (
            .O(N__26701),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ));
    CascadeMux I__4372 (
            .O(N__26698),
            .I(\phase_controller_inst1.stoper_tr.N_21_cascade_ ));
    CascadeMux I__4371 (
            .O(N__26695),
            .I(N__26692));
    InMux I__4370 (
            .O(N__26692),
            .I(N__26688));
    InMux I__4369 (
            .O(N__26691),
            .I(N__26684));
    LocalMux I__4368 (
            .O(N__26688),
            .I(N__26681));
    InMux I__4367 (
            .O(N__26687),
            .I(N__26678));
    LocalMux I__4366 (
            .O(N__26684),
            .I(N__26674));
    Span4Mux_h I__4365 (
            .O(N__26681),
            .I(N__26671));
    LocalMux I__4364 (
            .O(N__26678),
            .I(N__26668));
    InMux I__4363 (
            .O(N__26677),
            .I(N__26665));
    Span4Mux_h I__4362 (
            .O(N__26674),
            .I(N__26662));
    Odrv4 I__4361 (
            .O(N__26671),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__4360 (
            .O(N__26668),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__4359 (
            .O(N__26665),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__4358 (
            .O(N__26662),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__4357 (
            .O(N__26653),
            .I(N__26650));
    LocalMux I__4356 (
            .O(N__26650),
            .I(N__26647));
    Span4Mux_h I__4355 (
            .O(N__26647),
            .I(N__26643));
    InMux I__4354 (
            .O(N__26646),
            .I(N__26638));
    Span4Mux_h I__4353 (
            .O(N__26643),
            .I(N__26635));
    InMux I__4352 (
            .O(N__26642),
            .I(N__26632));
    InMux I__4351 (
            .O(N__26641),
            .I(N__26629));
    LocalMux I__4350 (
            .O(N__26638),
            .I(N__26626));
    Odrv4 I__4349 (
            .O(N__26635),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__4348 (
            .O(N__26632),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__4347 (
            .O(N__26629),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__4346 (
            .O(N__26626),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__4345 (
            .O(N__26617),
            .I(N__26614));
    InMux I__4344 (
            .O(N__26614),
            .I(N__26609));
    CascadeMux I__4343 (
            .O(N__26613),
            .I(N__26606));
    InMux I__4342 (
            .O(N__26612),
            .I(N__26603));
    LocalMux I__4341 (
            .O(N__26609),
            .I(N__26599));
    InMux I__4340 (
            .O(N__26606),
            .I(N__26596));
    LocalMux I__4339 (
            .O(N__26603),
            .I(N__26593));
    InMux I__4338 (
            .O(N__26602),
            .I(N__26590));
    Span4Mux_h I__4337 (
            .O(N__26599),
            .I(N__26587));
    LocalMux I__4336 (
            .O(N__26596),
            .I(N__26584));
    Odrv4 I__4335 (
            .O(N__26593),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__4334 (
            .O(N__26590),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__4333 (
            .O(N__26587),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__4332 (
            .O(N__26584),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__4331 (
            .O(N__26575),
            .I(N__26571));
    InMux I__4330 (
            .O(N__26574),
            .I(N__26568));
    LocalMux I__4329 (
            .O(N__26571),
            .I(N__26564));
    LocalMux I__4328 (
            .O(N__26568),
            .I(N__26560));
    InMux I__4327 (
            .O(N__26567),
            .I(N__26557));
    Span4Mux_h I__4326 (
            .O(N__26564),
            .I(N__26554));
    InMux I__4325 (
            .O(N__26563),
            .I(N__26551));
    Odrv4 I__4324 (
            .O(N__26560),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__4323 (
            .O(N__26557),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__4322 (
            .O(N__26554),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__4321 (
            .O(N__26551),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    CascadeMux I__4320 (
            .O(N__26542),
            .I(N__26539));
    InMux I__4319 (
            .O(N__26539),
            .I(N__26536));
    LocalMux I__4318 (
            .O(N__26536),
            .I(N__26533));
    Odrv4 I__4317 (
            .O(N__26533),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31 ));
    InMux I__4316 (
            .O(N__26530),
            .I(N__26527));
    LocalMux I__4315 (
            .O(N__26527),
            .I(N__26522));
    InMux I__4314 (
            .O(N__26526),
            .I(N__26519));
    InMux I__4313 (
            .O(N__26525),
            .I(N__26515));
    Span4Mux_v I__4312 (
            .O(N__26522),
            .I(N__26512));
    LocalMux I__4311 (
            .O(N__26519),
            .I(N__26509));
    InMux I__4310 (
            .O(N__26518),
            .I(N__26506));
    LocalMux I__4309 (
            .O(N__26515),
            .I(N__26503));
    Span4Mux_h I__4308 (
            .O(N__26512),
            .I(N__26498));
    Span4Mux_h I__4307 (
            .O(N__26509),
            .I(N__26498));
    LocalMux I__4306 (
            .O(N__26506),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__4305 (
            .O(N__26503),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__4304 (
            .O(N__26498),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__4303 (
            .O(N__26491),
            .I(N__26486));
    InMux I__4302 (
            .O(N__26490),
            .I(N__26483));
    InMux I__4301 (
            .O(N__26489),
            .I(N__26479));
    LocalMux I__4300 (
            .O(N__26486),
            .I(N__26476));
    LocalMux I__4299 (
            .O(N__26483),
            .I(N__26473));
    InMux I__4298 (
            .O(N__26482),
            .I(N__26470));
    LocalMux I__4297 (
            .O(N__26479),
            .I(N__26467));
    Span4Mux_h I__4296 (
            .O(N__26476),
            .I(N__26464));
    Odrv12 I__4295 (
            .O(N__26473),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__4294 (
            .O(N__26470),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__4293 (
            .O(N__26467),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__4292 (
            .O(N__26464),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    CascadeMux I__4291 (
            .O(N__26455),
            .I(N__26450));
    CascadeMux I__4290 (
            .O(N__26454),
            .I(N__26447));
    CascadeMux I__4289 (
            .O(N__26453),
            .I(N__26444));
    InMux I__4288 (
            .O(N__26450),
            .I(N__26441));
    InMux I__4287 (
            .O(N__26447),
            .I(N__26437));
    InMux I__4286 (
            .O(N__26444),
            .I(N__26434));
    LocalMux I__4285 (
            .O(N__26441),
            .I(N__26431));
    CascadeMux I__4284 (
            .O(N__26440),
            .I(N__26428));
    LocalMux I__4283 (
            .O(N__26437),
            .I(N__26423));
    LocalMux I__4282 (
            .O(N__26434),
            .I(N__26423));
    Span4Mux_h I__4281 (
            .O(N__26431),
            .I(N__26420));
    InMux I__4280 (
            .O(N__26428),
            .I(N__26417));
    Span4Mux_v I__4279 (
            .O(N__26423),
            .I(N__26414));
    Odrv4 I__4278 (
            .O(N__26420),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__4277 (
            .O(N__26417),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__4276 (
            .O(N__26414),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__4275 (
            .O(N__26407),
            .I(N__26403));
    InMux I__4274 (
            .O(N__26406),
            .I(N__26398));
    LocalMux I__4273 (
            .O(N__26403),
            .I(N__26395));
    InMux I__4272 (
            .O(N__26402),
            .I(N__26392));
    InMux I__4271 (
            .O(N__26401),
            .I(N__26389));
    LocalMux I__4270 (
            .O(N__26398),
            .I(N__26386));
    Odrv12 I__4269 (
            .O(N__26395),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__4268 (
            .O(N__26392),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__4267 (
            .O(N__26389),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__4266 (
            .O(N__26386),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__4265 (
            .O(N__26377),
            .I(N__26372));
    InMux I__4264 (
            .O(N__26376),
            .I(N__26369));
    InMux I__4263 (
            .O(N__26375),
            .I(N__26366));
    LocalMux I__4262 (
            .O(N__26372),
            .I(N__26362));
    LocalMux I__4261 (
            .O(N__26369),
            .I(N__26359));
    LocalMux I__4260 (
            .O(N__26366),
            .I(N__26356));
    InMux I__4259 (
            .O(N__26365),
            .I(N__26353));
    Span4Mux_h I__4258 (
            .O(N__26362),
            .I(N__26350));
    Span4Mux_h I__4257 (
            .O(N__26359),
            .I(N__26347));
    Odrv4 I__4256 (
            .O(N__26356),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__4255 (
            .O(N__26353),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__4254 (
            .O(N__26350),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__4253 (
            .O(N__26347),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__4252 (
            .O(N__26338),
            .I(N__26333));
    InMux I__4251 (
            .O(N__26337),
            .I(N__26330));
    InMux I__4250 (
            .O(N__26336),
            .I(N__26326));
    LocalMux I__4249 (
            .O(N__26333),
            .I(N__26323));
    LocalMux I__4248 (
            .O(N__26330),
            .I(N__26320));
    InMux I__4247 (
            .O(N__26329),
            .I(N__26317));
    LocalMux I__4246 (
            .O(N__26326),
            .I(N__26314));
    Span4Mux_h I__4245 (
            .O(N__26323),
            .I(N__26311));
    Odrv4 I__4244 (
            .O(N__26320),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__4243 (
            .O(N__26317),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__4242 (
            .O(N__26314),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__4241 (
            .O(N__26311),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__4240 (
            .O(N__26302),
            .I(N__26298));
    CascadeMux I__4239 (
            .O(N__26301),
            .I(N__26295));
    InMux I__4238 (
            .O(N__26298),
            .I(N__26291));
    InMux I__4237 (
            .O(N__26295),
            .I(N__26288));
    InMux I__4236 (
            .O(N__26294),
            .I(N__26285));
    LocalMux I__4235 (
            .O(N__26291),
            .I(N__26281));
    LocalMux I__4234 (
            .O(N__26288),
            .I(N__26278));
    LocalMux I__4233 (
            .O(N__26285),
            .I(N__26275));
    InMux I__4232 (
            .O(N__26284),
            .I(N__26272));
    Span4Mux_h I__4231 (
            .O(N__26281),
            .I(N__26269));
    Span4Mux_h I__4230 (
            .O(N__26278),
            .I(N__26266));
    Odrv12 I__4229 (
            .O(N__26275),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__4228 (
            .O(N__26272),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__4227 (
            .O(N__26269),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__4226 (
            .O(N__26266),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__4225 (
            .O(N__26257),
            .I(N__26252));
    InMux I__4224 (
            .O(N__26256),
            .I(N__26249));
    InMux I__4223 (
            .O(N__26255),
            .I(N__26245));
    LocalMux I__4222 (
            .O(N__26252),
            .I(N__26242));
    LocalMux I__4221 (
            .O(N__26249),
            .I(N__26239));
    InMux I__4220 (
            .O(N__26248),
            .I(N__26236));
    LocalMux I__4219 (
            .O(N__26245),
            .I(N__26233));
    Span4Mux_h I__4218 (
            .O(N__26242),
            .I(N__26230));
    Odrv4 I__4217 (
            .O(N__26239),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__4216 (
            .O(N__26236),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__4215 (
            .O(N__26233),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__4214 (
            .O(N__26230),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__4213 (
            .O(N__26221),
            .I(N__26218));
    LocalMux I__4212 (
            .O(N__26218),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ));
    InMux I__4211 (
            .O(N__26215),
            .I(N__26212));
    LocalMux I__4210 (
            .O(N__26212),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ));
    CascadeMux I__4209 (
            .O(N__26209),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ));
    InMux I__4208 (
            .O(N__26206),
            .I(N__26200));
    InMux I__4207 (
            .O(N__26205),
            .I(N__26200));
    LocalMux I__4206 (
            .O(N__26200),
            .I(N__26197));
    Span4Mux_h I__4205 (
            .O(N__26197),
            .I(N__26194));
    Odrv4 I__4204 (
            .O(N__26194),
            .I(\current_shift_inst.PI_CTRL.N_46_21 ));
    CascadeMux I__4203 (
            .O(N__26191),
            .I(N__26187));
    CascadeMux I__4202 (
            .O(N__26190),
            .I(N__26184));
    InMux I__4201 (
            .O(N__26187),
            .I(N__26181));
    InMux I__4200 (
            .O(N__26184),
            .I(N__26177));
    LocalMux I__4199 (
            .O(N__26181),
            .I(N__26173));
    CascadeMux I__4198 (
            .O(N__26180),
            .I(N__26170));
    LocalMux I__4197 (
            .O(N__26177),
            .I(N__26167));
    InMux I__4196 (
            .O(N__26176),
            .I(N__26164));
    Span4Mux_h I__4195 (
            .O(N__26173),
            .I(N__26161));
    InMux I__4194 (
            .O(N__26170),
            .I(N__26158));
    Span4Mux_h I__4193 (
            .O(N__26167),
            .I(N__26153));
    LocalMux I__4192 (
            .O(N__26164),
            .I(N__26153));
    Odrv4 I__4191 (
            .O(N__26161),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__4190 (
            .O(N__26158),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__4189 (
            .O(N__26153),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    CascadeMux I__4188 (
            .O(N__26146),
            .I(\phase_controller_inst1.N_232_cascade_ ));
    InMux I__4187 (
            .O(N__26143),
            .I(N__26140));
    LocalMux I__4186 (
            .O(N__26140),
            .I(N__26135));
    InMux I__4185 (
            .O(N__26139),
            .I(N__26132));
    InMux I__4184 (
            .O(N__26138),
            .I(N__26129));
    Span4Mux_v I__4183 (
            .O(N__26135),
            .I(N__26126));
    LocalMux I__4182 (
            .O(N__26132),
            .I(N__26121));
    LocalMux I__4181 (
            .O(N__26129),
            .I(N__26121));
    Span4Mux_v I__4180 (
            .O(N__26126),
            .I(N__26118));
    Span12Mux_h I__4179 (
            .O(N__26121),
            .I(N__26115));
    Odrv4 I__4178 (
            .O(N__26118),
            .I(il_max_comp1_D2));
    Odrv12 I__4177 (
            .O(N__26115),
            .I(il_max_comp1_D2));
    InMux I__4176 (
            .O(N__26110),
            .I(N__26107));
    LocalMux I__4175 (
            .O(N__26107),
            .I(N__26104));
    Odrv4 I__4174 (
            .O(N__26104),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__4173 (
            .O(N__26101),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__4172 (
            .O(N__26098),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__4171 (
            .O(N__26095),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__4170 (
            .O(N__26092),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__4169 (
            .O(N__26089),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__4168 (
            .O(N__26086),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__4167 (
            .O(N__26083),
            .I(bfn_10_13_0_));
    InMux I__4166 (
            .O(N__26080),
            .I(\pwm_generator_inst.counter_cry_8 ));
    CascadeMux I__4165 (
            .O(N__26077),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_ ));
    InMux I__4164 (
            .O(N__26074),
            .I(N__26071));
    LocalMux I__4163 (
            .O(N__26071),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto13 ));
    InMux I__4162 (
            .O(N__26068),
            .I(N__26063));
    InMux I__4161 (
            .O(N__26067),
            .I(N__26060));
    InMux I__4160 (
            .O(N__26066),
            .I(N__26057));
    LocalMux I__4159 (
            .O(N__26063),
            .I(measured_delay_hc_19));
    LocalMux I__4158 (
            .O(N__26060),
            .I(measured_delay_hc_19));
    LocalMux I__4157 (
            .O(N__26057),
            .I(measured_delay_hc_19));
    CascadeMux I__4156 (
            .O(N__26050),
            .I(N__26047));
    InMux I__4155 (
            .O(N__26047),
            .I(N__26044));
    LocalMux I__4154 (
            .O(N__26044),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ));
    InMux I__4153 (
            .O(N__26041),
            .I(bfn_10_12_0_));
    InMux I__4152 (
            .O(N__26038),
            .I(\pwm_generator_inst.counter_cry_0 ));
    CascadeMux I__4151 (
            .O(N__26035),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_ ));
    InMux I__4150 (
            .O(N__26032),
            .I(N__26029));
    LocalMux I__4149 (
            .O(N__26029),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz ));
    CascadeMux I__4148 (
            .O(N__26026),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30_cascade_ ));
    InMux I__4147 (
            .O(N__26023),
            .I(N__26020));
    LocalMux I__4146 (
            .O(N__26020),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ));
    InMux I__4145 (
            .O(N__26017),
            .I(N__26014));
    LocalMux I__4144 (
            .O(N__26014),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    CascadeMux I__4143 (
            .O(N__26011),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_ ));
    InMux I__4142 (
            .O(N__26008),
            .I(N__26003));
    InMux I__4141 (
            .O(N__26007),
            .I(N__26000));
    InMux I__4140 (
            .O(N__26006),
            .I(N__25997));
    LocalMux I__4139 (
            .O(N__26003),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__4138 (
            .O(N__26000),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__4137 (
            .O(N__25997),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    InMux I__4136 (
            .O(N__25990),
            .I(N__25985));
    InMux I__4135 (
            .O(N__25989),
            .I(N__25982));
    InMux I__4134 (
            .O(N__25988),
            .I(N__25979));
    LocalMux I__4133 (
            .O(N__25985),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__4132 (
            .O(N__25982),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__4131 (
            .O(N__25979),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    InMux I__4130 (
            .O(N__25972),
            .I(N__25966));
    InMux I__4129 (
            .O(N__25971),
            .I(N__25963));
    InMux I__4128 (
            .O(N__25970),
            .I(N__25960));
    InMux I__4127 (
            .O(N__25969),
            .I(N__25957));
    LocalMux I__4126 (
            .O(N__25966),
            .I(N__25952));
    LocalMux I__4125 (
            .O(N__25963),
            .I(N__25952));
    LocalMux I__4124 (
            .O(N__25960),
            .I(delay_hc_d2));
    LocalMux I__4123 (
            .O(N__25957),
            .I(delay_hc_d2));
    Odrv4 I__4122 (
            .O(N__25952),
            .I(delay_hc_d2));
    InMux I__4121 (
            .O(N__25945),
            .I(N__25941));
    InMux I__4120 (
            .O(N__25944),
            .I(N__25938));
    LocalMux I__4119 (
            .O(N__25941),
            .I(measured_delay_hc_26));
    LocalMux I__4118 (
            .O(N__25938),
            .I(measured_delay_hc_26));
    CascadeMux I__4117 (
            .O(N__25933),
            .I(N__25929));
    InMux I__4116 (
            .O(N__25932),
            .I(N__25926));
    InMux I__4115 (
            .O(N__25929),
            .I(N__25923));
    LocalMux I__4114 (
            .O(N__25926),
            .I(measured_delay_hc_30));
    LocalMux I__4113 (
            .O(N__25923),
            .I(measured_delay_hc_30));
    InMux I__4112 (
            .O(N__25918),
            .I(N__25914));
    InMux I__4111 (
            .O(N__25917),
            .I(N__25911));
    LocalMux I__4110 (
            .O(N__25914),
            .I(measured_delay_hc_25));
    LocalMux I__4109 (
            .O(N__25911),
            .I(measured_delay_hc_25));
    InMux I__4108 (
            .O(N__25906),
            .I(N__25902));
    InMux I__4107 (
            .O(N__25905),
            .I(N__25899));
    LocalMux I__4106 (
            .O(N__25902),
            .I(measured_delay_hc_23));
    LocalMux I__4105 (
            .O(N__25899),
            .I(measured_delay_hc_23));
    InMux I__4104 (
            .O(N__25894),
            .I(N__25890));
    InMux I__4103 (
            .O(N__25893),
            .I(N__25887));
    LocalMux I__4102 (
            .O(N__25890),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__4101 (
            .O(N__25887),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__4100 (
            .O(N__25882),
            .I(N__25878));
    InMux I__4099 (
            .O(N__25881),
            .I(N__25875));
    LocalMux I__4098 (
            .O(N__25878),
            .I(measured_delay_hc_24));
    LocalMux I__4097 (
            .O(N__25875),
            .I(measured_delay_hc_24));
    InMux I__4096 (
            .O(N__25870),
            .I(N__25866));
    InMux I__4095 (
            .O(N__25869),
            .I(N__25863));
    LocalMux I__4094 (
            .O(N__25866),
            .I(measured_delay_hc_29));
    LocalMux I__4093 (
            .O(N__25863),
            .I(measured_delay_hc_29));
    InMux I__4092 (
            .O(N__25858),
            .I(N__25855));
    LocalMux I__4091 (
            .O(N__25855),
            .I(N__25852));
    Odrv4 I__4090 (
            .O(N__25852),
            .I(\current_shift_inst.S3_syncZ0Z0 ));
    InMux I__4089 (
            .O(N__25849),
            .I(N__25843));
    InMux I__4088 (
            .O(N__25848),
            .I(N__25843));
    LocalMux I__4087 (
            .O(N__25843),
            .I(\current_shift_inst.S3_syncZ0Z1 ));
    InMux I__4086 (
            .O(N__25840),
            .I(N__25837));
    LocalMux I__4085 (
            .O(N__25837),
            .I(\current_shift_inst.S3_sync_prevZ0 ));
    InMux I__4084 (
            .O(N__25834),
            .I(N__25831));
    LocalMux I__4083 (
            .O(N__25831),
            .I(N__25828));
    IoSpan4Mux I__4082 (
            .O(N__25828),
            .I(N__25825));
    Odrv4 I__4081 (
            .O(N__25825),
            .I(il_min_comp2_c));
    CascadeMux I__4080 (
            .O(N__25822),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3_cascade_ ));
    InMux I__4079 (
            .O(N__25819),
            .I(N__25816));
    LocalMux I__4078 (
            .O(N__25816),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4 ));
    InMux I__4077 (
            .O(N__25813),
            .I(N__25809));
    CascadeMux I__4076 (
            .O(N__25812),
            .I(N__25806));
    LocalMux I__4075 (
            .O(N__25809),
            .I(N__25802));
    InMux I__4074 (
            .O(N__25806),
            .I(N__25796));
    InMux I__4073 (
            .O(N__25805),
            .I(N__25796));
    Span4Mux_v I__4072 (
            .O(N__25802),
            .I(N__25790));
    InMux I__4071 (
            .O(N__25801),
            .I(N__25787));
    LocalMux I__4070 (
            .O(N__25796),
            .I(N__25784));
    InMux I__4069 (
            .O(N__25795),
            .I(N__25779));
    InMux I__4068 (
            .O(N__25794),
            .I(N__25779));
    InMux I__4067 (
            .O(N__25793),
            .I(N__25776));
    Odrv4 I__4066 (
            .O(N__25790),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    LocalMux I__4065 (
            .O(N__25787),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    Odrv4 I__4064 (
            .O(N__25784),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    LocalMux I__4063 (
            .O(N__25779),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    LocalMux I__4062 (
            .O(N__25776),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    CascadeMux I__4061 (
            .O(N__25765),
            .I(N__25762));
    InMux I__4060 (
            .O(N__25762),
            .I(N__25758));
    CascadeMux I__4059 (
            .O(N__25761),
            .I(N__25754));
    LocalMux I__4058 (
            .O(N__25758),
            .I(N__25751));
    InMux I__4057 (
            .O(N__25757),
            .I(N__25748));
    InMux I__4056 (
            .O(N__25754),
            .I(N__25745));
    Odrv12 I__4055 (
            .O(N__25751),
            .I(\current_shift_inst.S3_riseZ0 ));
    LocalMux I__4054 (
            .O(N__25748),
            .I(\current_shift_inst.S3_riseZ0 ));
    LocalMux I__4053 (
            .O(N__25745),
            .I(\current_shift_inst.S3_riseZ0 ));
    InMux I__4052 (
            .O(N__25738),
            .I(N__25735));
    LocalMux I__4051 (
            .O(N__25735),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__4050 (
            .O(N__25732),
            .I(N__25729));
    InMux I__4049 (
            .O(N__25729),
            .I(N__25726));
    LocalMux I__4048 (
            .O(N__25726),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__4047 (
            .O(N__25723),
            .I(N__25720));
    LocalMux I__4046 (
            .O(N__25720),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    CascadeMux I__4045 (
            .O(N__25717),
            .I(N__25714));
    InMux I__4044 (
            .O(N__25714),
            .I(N__25711));
    LocalMux I__4043 (
            .O(N__25711),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    CascadeMux I__4042 (
            .O(N__25708),
            .I(N__25700));
    InMux I__4041 (
            .O(N__25707),
            .I(N__25685));
    InMux I__4040 (
            .O(N__25706),
            .I(N__25685));
    InMux I__4039 (
            .O(N__25705),
            .I(N__25685));
    InMux I__4038 (
            .O(N__25704),
            .I(N__25685));
    InMux I__4037 (
            .O(N__25703),
            .I(N__25685));
    InMux I__4036 (
            .O(N__25700),
            .I(N__25678));
    InMux I__4035 (
            .O(N__25699),
            .I(N__25678));
    InMux I__4034 (
            .O(N__25698),
            .I(N__25678));
    CascadeMux I__4033 (
            .O(N__25697),
            .I(N__25673));
    InMux I__4032 (
            .O(N__25696),
            .I(N__25667));
    LocalMux I__4031 (
            .O(N__25685),
            .I(N__25662));
    LocalMux I__4030 (
            .O(N__25678),
            .I(N__25662));
    InMux I__4029 (
            .O(N__25677),
            .I(N__25659));
    InMux I__4028 (
            .O(N__25676),
            .I(N__25646));
    InMux I__4027 (
            .O(N__25673),
            .I(N__25637));
    InMux I__4026 (
            .O(N__25672),
            .I(N__25637));
    InMux I__4025 (
            .O(N__25671),
            .I(N__25637));
    InMux I__4024 (
            .O(N__25670),
            .I(N__25637));
    LocalMux I__4023 (
            .O(N__25667),
            .I(N__25634));
    Span4Mux_v I__4022 (
            .O(N__25662),
            .I(N__25631));
    LocalMux I__4021 (
            .O(N__25659),
            .I(N__25628));
    InMux I__4020 (
            .O(N__25658),
            .I(N__25623));
    InMux I__4019 (
            .O(N__25657),
            .I(N__25623));
    CascadeMux I__4018 (
            .O(N__25656),
            .I(N__25618));
    CascadeMux I__4017 (
            .O(N__25655),
            .I(N__25615));
    InMux I__4016 (
            .O(N__25654),
            .I(N__25607));
    InMux I__4015 (
            .O(N__25653),
            .I(N__25607));
    InMux I__4014 (
            .O(N__25652),
            .I(N__25607));
    InMux I__4013 (
            .O(N__25651),
            .I(N__25600));
    InMux I__4012 (
            .O(N__25650),
            .I(N__25600));
    InMux I__4011 (
            .O(N__25649),
            .I(N__25600));
    LocalMux I__4010 (
            .O(N__25646),
            .I(N__25595));
    LocalMux I__4009 (
            .O(N__25637),
            .I(N__25595));
    Span4Mux_v I__4008 (
            .O(N__25634),
            .I(N__25586));
    Span4Mux_h I__4007 (
            .O(N__25631),
            .I(N__25586));
    Span4Mux_v I__4006 (
            .O(N__25628),
            .I(N__25586));
    LocalMux I__4005 (
            .O(N__25623),
            .I(N__25586));
    InMux I__4004 (
            .O(N__25622),
            .I(N__25575));
    InMux I__4003 (
            .O(N__25621),
            .I(N__25575));
    InMux I__4002 (
            .O(N__25618),
            .I(N__25575));
    InMux I__4001 (
            .O(N__25615),
            .I(N__25575));
    InMux I__4000 (
            .O(N__25614),
            .I(N__25575));
    LocalMux I__3999 (
            .O(N__25607),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    LocalMux I__3998 (
            .O(N__25600),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__3997 (
            .O(N__25595),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__3996 (
            .O(N__25586),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    LocalMux I__3995 (
            .O(N__25575),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    InMux I__3994 (
            .O(N__25564),
            .I(N__25561));
    LocalMux I__3993 (
            .O(N__25561),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    CascadeMux I__3992 (
            .O(N__25558),
            .I(N__25555));
    InMux I__3991 (
            .O(N__25555),
            .I(N__25541));
    CascadeMux I__3990 (
            .O(N__25554),
            .I(N__25538));
    CascadeMux I__3989 (
            .O(N__25553),
            .I(N__25535));
    CascadeMux I__3988 (
            .O(N__25552),
            .I(N__25532));
    CascadeMux I__3987 (
            .O(N__25551),
            .I(N__25529));
    CascadeMux I__3986 (
            .O(N__25550),
            .I(N__25523));
    CascadeMux I__3985 (
            .O(N__25549),
            .I(N__25517));
    CascadeMux I__3984 (
            .O(N__25548),
            .I(N__25514));
    CascadeMux I__3983 (
            .O(N__25547),
            .I(N__25511));
    CascadeMux I__3982 (
            .O(N__25546),
            .I(N__25506));
    CascadeMux I__3981 (
            .O(N__25545),
            .I(N__25503));
    CascadeMux I__3980 (
            .O(N__25544),
            .I(N__25500));
    LocalMux I__3979 (
            .O(N__25541),
            .I(N__25496));
    InMux I__3978 (
            .O(N__25538),
            .I(N__25493));
    InMux I__3977 (
            .O(N__25535),
            .I(N__25482));
    InMux I__3976 (
            .O(N__25532),
            .I(N__25482));
    InMux I__3975 (
            .O(N__25529),
            .I(N__25482));
    InMux I__3974 (
            .O(N__25528),
            .I(N__25482));
    InMux I__3973 (
            .O(N__25527),
            .I(N__25482));
    CascadeMux I__3972 (
            .O(N__25526),
            .I(N__25479));
    InMux I__3971 (
            .O(N__25523),
            .I(N__25470));
    CascadeMux I__3970 (
            .O(N__25522),
            .I(N__25467));
    CascadeMux I__3969 (
            .O(N__25521),
            .I(N__25463));
    InMux I__3968 (
            .O(N__25520),
            .I(N__25460));
    InMux I__3967 (
            .O(N__25517),
            .I(N__25449));
    InMux I__3966 (
            .O(N__25514),
            .I(N__25449));
    InMux I__3965 (
            .O(N__25511),
            .I(N__25449));
    InMux I__3964 (
            .O(N__25510),
            .I(N__25449));
    InMux I__3963 (
            .O(N__25509),
            .I(N__25449));
    InMux I__3962 (
            .O(N__25506),
            .I(N__25440));
    InMux I__3961 (
            .O(N__25503),
            .I(N__25440));
    InMux I__3960 (
            .O(N__25500),
            .I(N__25440));
    InMux I__3959 (
            .O(N__25499),
            .I(N__25440));
    Span4Mux_h I__3958 (
            .O(N__25496),
            .I(N__25433));
    LocalMux I__3957 (
            .O(N__25493),
            .I(N__25433));
    LocalMux I__3956 (
            .O(N__25482),
            .I(N__25433));
    InMux I__3955 (
            .O(N__25479),
            .I(N__25428));
    InMux I__3954 (
            .O(N__25478),
            .I(N__25428));
    CascadeMux I__3953 (
            .O(N__25477),
            .I(N__25425));
    CascadeMux I__3952 (
            .O(N__25476),
            .I(N__25422));
    CascadeMux I__3951 (
            .O(N__25475),
            .I(N__25418));
    CascadeMux I__3950 (
            .O(N__25474),
            .I(N__25414));
    CascadeMux I__3949 (
            .O(N__25473),
            .I(N__25411));
    LocalMux I__3948 (
            .O(N__25470),
            .I(N__25407));
    InMux I__3947 (
            .O(N__25467),
            .I(N__25402));
    InMux I__3946 (
            .O(N__25466),
            .I(N__25402));
    InMux I__3945 (
            .O(N__25463),
            .I(N__25398));
    LocalMux I__3944 (
            .O(N__25460),
            .I(N__25395));
    LocalMux I__3943 (
            .O(N__25449),
            .I(N__25386));
    LocalMux I__3942 (
            .O(N__25440),
            .I(N__25386));
    Span4Mux_h I__3941 (
            .O(N__25433),
            .I(N__25386));
    LocalMux I__3940 (
            .O(N__25428),
            .I(N__25386));
    InMux I__3939 (
            .O(N__25425),
            .I(N__25379));
    InMux I__3938 (
            .O(N__25422),
            .I(N__25379));
    InMux I__3937 (
            .O(N__25421),
            .I(N__25379));
    InMux I__3936 (
            .O(N__25418),
            .I(N__25374));
    InMux I__3935 (
            .O(N__25417),
            .I(N__25374));
    InMux I__3934 (
            .O(N__25414),
            .I(N__25367));
    InMux I__3933 (
            .O(N__25411),
            .I(N__25367));
    InMux I__3932 (
            .O(N__25410),
            .I(N__25367));
    Span4Mux_h I__3931 (
            .O(N__25407),
            .I(N__25364));
    LocalMux I__3930 (
            .O(N__25402),
            .I(N__25361));
    InMux I__3929 (
            .O(N__25401),
            .I(N__25358));
    LocalMux I__3928 (
            .O(N__25398),
            .I(N__25351));
    Span4Mux_h I__3927 (
            .O(N__25395),
            .I(N__25351));
    Span4Mux_v I__3926 (
            .O(N__25386),
            .I(N__25351));
    LocalMux I__3925 (
            .O(N__25379),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3924 (
            .O(N__25374),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3923 (
            .O(N__25367),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3922 (
            .O(N__25364),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__3921 (
            .O(N__25361),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3920 (
            .O(N__25358),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3919 (
            .O(N__25351),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__3918 (
            .O(N__25336),
            .I(N__25318));
    InMux I__3917 (
            .O(N__25335),
            .I(N__25307));
    InMux I__3916 (
            .O(N__25334),
            .I(N__25307));
    InMux I__3915 (
            .O(N__25333),
            .I(N__25307));
    InMux I__3914 (
            .O(N__25332),
            .I(N__25307));
    InMux I__3913 (
            .O(N__25331),
            .I(N__25307));
    InMux I__3912 (
            .O(N__25330),
            .I(N__25300));
    InMux I__3911 (
            .O(N__25329),
            .I(N__25300));
    InMux I__3910 (
            .O(N__25328),
            .I(N__25300));
    InMux I__3909 (
            .O(N__25327),
            .I(N__25295));
    InMux I__3908 (
            .O(N__25326),
            .I(N__25295));
    InMux I__3907 (
            .O(N__25325),
            .I(N__25286));
    InMux I__3906 (
            .O(N__25324),
            .I(N__25277));
    InMux I__3905 (
            .O(N__25323),
            .I(N__25277));
    InMux I__3904 (
            .O(N__25322),
            .I(N__25277));
    InMux I__3903 (
            .O(N__25321),
            .I(N__25277));
    LocalMux I__3902 (
            .O(N__25318),
            .I(N__25274));
    LocalMux I__3901 (
            .O(N__25307),
            .I(N__25267));
    LocalMux I__3900 (
            .O(N__25300),
            .I(N__25267));
    LocalMux I__3899 (
            .O(N__25295),
            .I(N__25267));
    InMux I__3898 (
            .O(N__25294),
            .I(N__25264));
    InMux I__3897 (
            .O(N__25293),
            .I(N__25253));
    InMux I__3896 (
            .O(N__25292),
            .I(N__25253));
    InMux I__3895 (
            .O(N__25291),
            .I(N__25253));
    InMux I__3894 (
            .O(N__25290),
            .I(N__25253));
    InMux I__3893 (
            .O(N__25289),
            .I(N__25253));
    LocalMux I__3892 (
            .O(N__25286),
            .I(N__25242));
    LocalMux I__3891 (
            .O(N__25277),
            .I(N__25242));
    Span4Mux_v I__3890 (
            .O(N__25274),
            .I(N__25235));
    Span4Mux_v I__3889 (
            .O(N__25267),
            .I(N__25235));
    LocalMux I__3888 (
            .O(N__25264),
            .I(N__25235));
    LocalMux I__3887 (
            .O(N__25253),
            .I(N__25232));
    InMux I__3886 (
            .O(N__25252),
            .I(N__25219));
    InMux I__3885 (
            .O(N__25251),
            .I(N__25219));
    InMux I__3884 (
            .O(N__25250),
            .I(N__25219));
    InMux I__3883 (
            .O(N__25249),
            .I(N__25219));
    InMux I__3882 (
            .O(N__25248),
            .I(N__25219));
    InMux I__3881 (
            .O(N__25247),
            .I(N__25219));
    Odrv12 I__3880 (
            .O(N__25242),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    Odrv4 I__3879 (
            .O(N__25235),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    Odrv4 I__3878 (
            .O(N__25232),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    LocalMux I__3877 (
            .O(N__25219),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    CEMux I__3876 (
            .O(N__25210),
            .I(N__25204));
    CEMux I__3875 (
            .O(N__25209),
            .I(N__25201));
    CEMux I__3874 (
            .O(N__25208),
            .I(N__25198));
    CEMux I__3873 (
            .O(N__25207),
            .I(N__25191));
    LocalMux I__3872 (
            .O(N__25204),
            .I(N__25188));
    LocalMux I__3871 (
            .O(N__25201),
            .I(N__25183));
    LocalMux I__3870 (
            .O(N__25198),
            .I(N__25183));
    CEMux I__3869 (
            .O(N__25197),
            .I(N__25180));
    CEMux I__3868 (
            .O(N__25196),
            .I(N__25175));
    CEMux I__3867 (
            .O(N__25195),
            .I(N__25169));
    CEMux I__3866 (
            .O(N__25194),
            .I(N__25166));
    LocalMux I__3865 (
            .O(N__25191),
            .I(N__25163));
    Span4Mux_h I__3864 (
            .O(N__25188),
            .I(N__25156));
    Span4Mux_v I__3863 (
            .O(N__25183),
            .I(N__25156));
    LocalMux I__3862 (
            .O(N__25180),
            .I(N__25156));
    CEMux I__3861 (
            .O(N__25179),
            .I(N__25149));
    CEMux I__3860 (
            .O(N__25178),
            .I(N__25146));
    LocalMux I__3859 (
            .O(N__25175),
            .I(N__25142));
    CEMux I__3858 (
            .O(N__25174),
            .I(N__25139));
    CEMux I__3857 (
            .O(N__25173),
            .I(N__25136));
    CEMux I__3856 (
            .O(N__25172),
            .I(N__25129));
    LocalMux I__3855 (
            .O(N__25169),
            .I(N__25124));
    LocalMux I__3854 (
            .O(N__25166),
            .I(N__25124));
    Span4Mux_h I__3853 (
            .O(N__25163),
            .I(N__25119));
    Span4Mux_v I__3852 (
            .O(N__25156),
            .I(N__25119));
    CEMux I__3851 (
            .O(N__25155),
            .I(N__25116));
    CEMux I__3850 (
            .O(N__25154),
            .I(N__25113));
    CEMux I__3849 (
            .O(N__25153),
            .I(N__25110));
    CEMux I__3848 (
            .O(N__25152),
            .I(N__25107));
    LocalMux I__3847 (
            .O(N__25149),
            .I(N__25101));
    LocalMux I__3846 (
            .O(N__25146),
            .I(N__25101));
    CEMux I__3845 (
            .O(N__25145),
            .I(N__25098));
    Span4Mux_v I__3844 (
            .O(N__25142),
            .I(N__25091));
    LocalMux I__3843 (
            .O(N__25139),
            .I(N__25091));
    LocalMux I__3842 (
            .O(N__25136),
            .I(N__25091));
    CEMux I__3841 (
            .O(N__25135),
            .I(N__25088));
    CEMux I__3840 (
            .O(N__25134),
            .I(N__25085));
    CEMux I__3839 (
            .O(N__25133),
            .I(N__25082));
    CEMux I__3838 (
            .O(N__25132),
            .I(N__25078));
    LocalMux I__3837 (
            .O(N__25129),
            .I(N__25074));
    Span4Mux_h I__3836 (
            .O(N__25124),
            .I(N__25065));
    Span4Mux_h I__3835 (
            .O(N__25119),
            .I(N__25065));
    LocalMux I__3834 (
            .O(N__25116),
            .I(N__25065));
    LocalMux I__3833 (
            .O(N__25113),
            .I(N__25065));
    LocalMux I__3832 (
            .O(N__25110),
            .I(N__25061));
    LocalMux I__3831 (
            .O(N__25107),
            .I(N__25058));
    CEMux I__3830 (
            .O(N__25106),
            .I(N__25055));
    Span4Mux_v I__3829 (
            .O(N__25101),
            .I(N__25049));
    LocalMux I__3828 (
            .O(N__25098),
            .I(N__25049));
    Span4Mux_h I__3827 (
            .O(N__25091),
            .I(N__25042));
    LocalMux I__3826 (
            .O(N__25088),
            .I(N__25042));
    LocalMux I__3825 (
            .O(N__25085),
            .I(N__25042));
    LocalMux I__3824 (
            .O(N__25082),
            .I(N__25039));
    CEMux I__3823 (
            .O(N__25081),
            .I(N__25036));
    LocalMux I__3822 (
            .O(N__25078),
            .I(N__25033));
    CEMux I__3821 (
            .O(N__25077),
            .I(N__25030));
    Span4Mux_v I__3820 (
            .O(N__25074),
            .I(N__25025));
    Span4Mux_v I__3819 (
            .O(N__25065),
            .I(N__25025));
    CEMux I__3818 (
            .O(N__25064),
            .I(N__25022));
    Span4Mux_v I__3817 (
            .O(N__25061),
            .I(N__25015));
    Span4Mux_h I__3816 (
            .O(N__25058),
            .I(N__25015));
    LocalMux I__3815 (
            .O(N__25055),
            .I(N__25015));
    CEMux I__3814 (
            .O(N__25054),
            .I(N__25012));
    Span4Mux_v I__3813 (
            .O(N__25049),
            .I(N__25007));
    Span4Mux_v I__3812 (
            .O(N__25042),
            .I(N__25007));
    Span4Mux_v I__3811 (
            .O(N__25039),
            .I(N__25002));
    LocalMux I__3810 (
            .O(N__25036),
            .I(N__25002));
    Span4Mux_v I__3809 (
            .O(N__25033),
            .I(N__24997));
    LocalMux I__3808 (
            .O(N__25030),
            .I(N__24997));
    Span4Mux_v I__3807 (
            .O(N__25025),
            .I(N__24994));
    LocalMux I__3806 (
            .O(N__25022),
            .I(N__24987));
    Sp12to4 I__3805 (
            .O(N__25015),
            .I(N__24987));
    LocalMux I__3804 (
            .O(N__25012),
            .I(N__24987));
    Span4Mux_v I__3803 (
            .O(N__25007),
            .I(N__24980));
    Span4Mux_v I__3802 (
            .O(N__25002),
            .I(N__24980));
    Span4Mux_s2_h I__3801 (
            .O(N__24997),
            .I(N__24980));
    Odrv4 I__3800 (
            .O(N__24994),
            .I(N_717_g));
    Odrv12 I__3799 (
            .O(N__24987),
            .I(N_717_g));
    Odrv4 I__3798 (
            .O(N__24980),
            .I(N_717_g));
    InMux I__3797 (
            .O(N__24973),
            .I(N__24969));
    InMux I__3796 (
            .O(N__24972),
            .I(N__24965));
    LocalMux I__3795 (
            .O(N__24969),
            .I(N__24961));
    InMux I__3794 (
            .O(N__24968),
            .I(N__24958));
    LocalMux I__3793 (
            .O(N__24965),
            .I(N__24955));
    InMux I__3792 (
            .O(N__24964),
            .I(N__24952));
    Span4Mux_h I__3791 (
            .O(N__24961),
            .I(N__24949));
    LocalMux I__3790 (
            .O(N__24958),
            .I(N__24946));
    Odrv12 I__3789 (
            .O(N__24955),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__3788 (
            .O(N__24952),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__3787 (
            .O(N__24949),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__3786 (
            .O(N__24946),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    InMux I__3785 (
            .O(N__24937),
            .I(N__24934));
    LocalMux I__3784 (
            .O(N__24934),
            .I(N__24931));
    Span4Mux_v I__3783 (
            .O(N__24931),
            .I(N__24927));
    InMux I__3782 (
            .O(N__24930),
            .I(N__24924));
    Span4Mux_h I__3781 (
            .O(N__24927),
            .I(N__24919));
    LocalMux I__3780 (
            .O(N__24924),
            .I(N__24916));
    InMux I__3779 (
            .O(N__24923),
            .I(N__24913));
    InMux I__3778 (
            .O(N__24922),
            .I(N__24910));
    Odrv4 I__3777 (
            .O(N__24919),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv12 I__3776 (
            .O(N__24916),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__3775 (
            .O(N__24913),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__3774 (
            .O(N__24910),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    CascadeMux I__3773 (
            .O(N__24901),
            .I(N__24896));
    CascadeMux I__3772 (
            .O(N__24900),
            .I(N__24893));
    InMux I__3771 (
            .O(N__24899),
            .I(N__24890));
    InMux I__3770 (
            .O(N__24896),
            .I(N__24887));
    InMux I__3769 (
            .O(N__24893),
            .I(N__24884));
    LocalMux I__3768 (
            .O(N__24890),
            .I(N__24880));
    LocalMux I__3767 (
            .O(N__24887),
            .I(N__24875));
    LocalMux I__3766 (
            .O(N__24884),
            .I(N__24875));
    InMux I__3765 (
            .O(N__24883),
            .I(N__24872));
    Span4Mux_h I__3764 (
            .O(N__24880),
            .I(N__24869));
    Span4Mux_h I__3763 (
            .O(N__24875),
            .I(N__24866));
    LocalMux I__3762 (
            .O(N__24872),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__3761 (
            .O(N__24869),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__3760 (
            .O(N__24866),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__3759 (
            .O(N__24859),
            .I(N__24853));
    InMux I__3758 (
            .O(N__24858),
            .I(N__24853));
    LocalMux I__3757 (
            .O(N__24853),
            .I(N__24850));
    Span4Mux_h I__3756 (
            .O(N__24850),
            .I(N__24847));
    Odrv4 I__3755 (
            .O(N__24847),
            .I(\current_shift_inst.PI_CTRL.N_46_16 ));
    InMux I__3754 (
            .O(N__24844),
            .I(N__24841));
    LocalMux I__3753 (
            .O(N__24841),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    CascadeMux I__3752 (
            .O(N__24838),
            .I(N__24835));
    InMux I__3751 (
            .O(N__24835),
            .I(N__24832));
    LocalMux I__3750 (
            .O(N__24832),
            .I(N__24829));
    Odrv4 I__3749 (
            .O(N__24829),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__3748 (
            .O(N__24826),
            .I(N__24822));
    CascadeMux I__3747 (
            .O(N__24825),
            .I(N__24818));
    LocalMux I__3746 (
            .O(N__24822),
            .I(N__24815));
    InMux I__3745 (
            .O(N__24821),
            .I(N__24812));
    InMux I__3744 (
            .O(N__24818),
            .I(N__24808));
    Span4Mux_v I__3743 (
            .O(N__24815),
            .I(N__24803));
    LocalMux I__3742 (
            .O(N__24812),
            .I(N__24803));
    InMux I__3741 (
            .O(N__24811),
            .I(N__24800));
    LocalMux I__3740 (
            .O(N__24808),
            .I(N__24795));
    Span4Mux_h I__3739 (
            .O(N__24803),
            .I(N__24795));
    LocalMux I__3738 (
            .O(N__24800),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__3737 (
            .O(N__24795),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__3736 (
            .O(N__24790),
            .I(N__24787));
    LocalMux I__3735 (
            .O(N__24787),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__3734 (
            .O(N__24784),
            .I(N__24781));
    LocalMux I__3733 (
            .O(N__24781),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__3732 (
            .O(N__24778),
            .I(N__24775));
    LocalMux I__3731 (
            .O(N__24775),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    CascadeMux I__3730 (
            .O(N__24772),
            .I(N__24769));
    InMux I__3729 (
            .O(N__24769),
            .I(N__24766));
    LocalMux I__3728 (
            .O(N__24766),
            .I(N__24763));
    Span4Mux_h I__3727 (
            .O(N__24763),
            .I(N__24760));
    Span4Mux_v I__3726 (
            .O(N__24760),
            .I(N__24757));
    Odrv4 I__3725 (
            .O(N__24757),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    InMux I__3724 (
            .O(N__24754),
            .I(N__24751));
    LocalMux I__3723 (
            .O(N__24751),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__3722 (
            .O(N__24748),
            .I(N__24745));
    InMux I__3721 (
            .O(N__24745),
            .I(N__24742));
    LocalMux I__3720 (
            .O(N__24742),
            .I(N__24739));
    Span4Mux_h I__3719 (
            .O(N__24739),
            .I(N__24736));
    Span4Mux_h I__3718 (
            .O(N__24736),
            .I(N__24733));
    Odrv4 I__3717 (
            .O(N__24733),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    InMux I__3716 (
            .O(N__24730),
            .I(N__24727));
    LocalMux I__3715 (
            .O(N__24727),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__3714 (
            .O(N__24724),
            .I(N__24721));
    InMux I__3713 (
            .O(N__24721),
            .I(N__24718));
    LocalMux I__3712 (
            .O(N__24718),
            .I(N__24715));
    Span4Mux_v I__3711 (
            .O(N__24715),
            .I(N__24712));
    Span4Mux_h I__3710 (
            .O(N__24712),
            .I(N__24709));
    Odrv4 I__3709 (
            .O(N__24709),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    InMux I__3708 (
            .O(N__24706),
            .I(N__24703));
    LocalMux I__3707 (
            .O(N__24703),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__3706 (
            .O(N__24700),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__3705 (
            .O(N__24697),
            .I(N__24694));
    LocalMux I__3704 (
            .O(N__24694),
            .I(N__24691));
    Span4Mux_s1_v I__3703 (
            .O(N__24691),
            .I(N__24688));
    Sp12to4 I__3702 (
            .O(N__24688),
            .I(N__24685));
    Span12Mux_h I__3701 (
            .O(N__24685),
            .I(N__24682));
    Odrv12 I__3700 (
            .O(N__24682),
            .I(pwm_output_c));
    CascadeMux I__3699 (
            .O(N__24679),
            .I(N__24676));
    InMux I__3698 (
            .O(N__24676),
            .I(N__24673));
    LocalMux I__3697 (
            .O(N__24673),
            .I(N__24670));
    Odrv12 I__3696 (
            .O(N__24670),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ));
    CascadeMux I__3695 (
            .O(N__24667),
            .I(N__24664));
    InMux I__3694 (
            .O(N__24664),
            .I(N__24661));
    LocalMux I__3693 (
            .O(N__24661),
            .I(N__24658));
    Span4Mux_h I__3692 (
            .O(N__24658),
            .I(N__24655));
    Odrv4 I__3691 (
            .O(N__24655),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__3690 (
            .O(N__24652),
            .I(N__24649));
    InMux I__3689 (
            .O(N__24649),
            .I(N__24646));
    LocalMux I__3688 (
            .O(N__24646),
            .I(N__24643));
    Span4Mux_h I__3687 (
            .O(N__24643),
            .I(N__24640));
    Odrv4 I__3686 (
            .O(N__24640),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CEMux I__3685 (
            .O(N__24637),
            .I(N__24633));
    CEMux I__3684 (
            .O(N__24636),
            .I(N__24630));
    LocalMux I__3683 (
            .O(N__24633),
            .I(N__24627));
    LocalMux I__3682 (
            .O(N__24630),
            .I(N__24623));
    Span4Mux_v I__3681 (
            .O(N__24627),
            .I(N__24618));
    CEMux I__3680 (
            .O(N__24626),
            .I(N__24615));
    Span4Mux_v I__3679 (
            .O(N__24623),
            .I(N__24612));
    CEMux I__3678 (
            .O(N__24622),
            .I(N__24609));
    CEMux I__3677 (
            .O(N__24621),
            .I(N__24606));
    Odrv4 I__3676 (
            .O(N__24618),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    LocalMux I__3675 (
            .O(N__24615),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__3674 (
            .O(N__24612),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    LocalMux I__3673 (
            .O(N__24609),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    LocalMux I__3672 (
            .O(N__24606),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__3671 (
            .O(N__24595),
            .I(N__24591));
    InMux I__3670 (
            .O(N__24594),
            .I(N__24588));
    LocalMux I__3669 (
            .O(N__24591),
            .I(N__24583));
    LocalMux I__3668 (
            .O(N__24588),
            .I(N__24580));
    InMux I__3667 (
            .O(N__24587),
            .I(N__24577));
    InMux I__3666 (
            .O(N__24586),
            .I(N__24574));
    Odrv4 I__3665 (
            .O(N__24583),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    Odrv4 I__3664 (
            .O(N__24580),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    LocalMux I__3663 (
            .O(N__24577),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    LocalMux I__3662 (
            .O(N__24574),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    CascadeMux I__3661 (
            .O(N__24565),
            .I(N__24562));
    InMux I__3660 (
            .O(N__24562),
            .I(N__24559));
    LocalMux I__3659 (
            .O(N__24559),
            .I(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__3658 (
            .O(N__24556),
            .I(N__24550));
    InMux I__3657 (
            .O(N__24555),
            .I(N__24543));
    InMux I__3656 (
            .O(N__24554),
            .I(N__24543));
    InMux I__3655 (
            .O(N__24553),
            .I(N__24543));
    LocalMux I__3654 (
            .O(N__24550),
            .I(N__24536));
    LocalMux I__3653 (
            .O(N__24543),
            .I(N__24536));
    InMux I__3652 (
            .O(N__24542),
            .I(N__24533));
    InMux I__3651 (
            .O(N__24541),
            .I(N__24530));
    Span4Mux_v I__3650 (
            .O(N__24536),
            .I(N__24525));
    LocalMux I__3649 (
            .O(N__24533),
            .I(N__24525));
    LocalMux I__3648 (
            .O(N__24530),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__3647 (
            .O(N__24525),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__3646 (
            .O(N__24520),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt8_cascade_ ));
    InMux I__3645 (
            .O(N__24517),
            .I(N__24514));
    LocalMux I__3644 (
            .O(N__24514),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt15 ));
    CascadeMux I__3643 (
            .O(N__24511),
            .I(N__24508));
    InMux I__3642 (
            .O(N__24508),
            .I(N__24505));
    LocalMux I__3641 (
            .O(N__24505),
            .I(N__24502));
    Span4Mux_h I__3640 (
            .O(N__24502),
            .I(N__24499));
    Span4Mux_v I__3639 (
            .O(N__24499),
            .I(N__24496));
    Odrv4 I__3638 (
            .O(N__24496),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    InMux I__3637 (
            .O(N__24493),
            .I(N__24490));
    LocalMux I__3636 (
            .O(N__24490),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__3635 (
            .O(N__24487),
            .I(N__24484));
    InMux I__3634 (
            .O(N__24484),
            .I(N__24481));
    LocalMux I__3633 (
            .O(N__24481),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    InMux I__3632 (
            .O(N__24478),
            .I(N__24475));
    LocalMux I__3631 (
            .O(N__24475),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__3630 (
            .O(N__24472),
            .I(N__24469));
    InMux I__3629 (
            .O(N__24469),
            .I(N__24466));
    LocalMux I__3628 (
            .O(N__24466),
            .I(N__24463));
    Span4Mux_v I__3627 (
            .O(N__24463),
            .I(N__24460));
    Odrv4 I__3626 (
            .O(N__24460),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    InMux I__3625 (
            .O(N__24457),
            .I(N__24454));
    LocalMux I__3624 (
            .O(N__24454),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__3623 (
            .O(N__24451),
            .I(N__24448));
    InMux I__3622 (
            .O(N__24448),
            .I(N__24445));
    LocalMux I__3621 (
            .O(N__24445),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    InMux I__3620 (
            .O(N__24442),
            .I(N__24439));
    LocalMux I__3619 (
            .O(N__24439),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__3618 (
            .O(N__24436),
            .I(N__24433));
    InMux I__3617 (
            .O(N__24433),
            .I(N__24430));
    LocalMux I__3616 (
            .O(N__24430),
            .I(N__24427));
    Odrv4 I__3615 (
            .O(N__24427),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    InMux I__3614 (
            .O(N__24424),
            .I(N__24421));
    LocalMux I__3613 (
            .O(N__24421),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__3612 (
            .O(N__24418),
            .I(N__24415));
    InMux I__3611 (
            .O(N__24415),
            .I(N__24412));
    LocalMux I__3610 (
            .O(N__24412),
            .I(N__24409));
    Span4Mux_v I__3609 (
            .O(N__24409),
            .I(N__24406));
    Odrv4 I__3608 (
            .O(N__24406),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    InMux I__3607 (
            .O(N__24403),
            .I(N__24400));
    LocalMux I__3606 (
            .O(N__24400),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__3605 (
            .O(N__24397),
            .I(N__24394));
    InMux I__3604 (
            .O(N__24394),
            .I(N__24391));
    LocalMux I__3603 (
            .O(N__24391),
            .I(N__24388));
    Span4Mux_v I__3602 (
            .O(N__24388),
            .I(N__24385));
    Span4Mux_h I__3601 (
            .O(N__24385),
            .I(N__24382));
    Odrv4 I__3600 (
            .O(N__24382),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    InMux I__3599 (
            .O(N__24379),
            .I(N__24376));
    LocalMux I__3598 (
            .O(N__24376),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__3597 (
            .O(N__24373),
            .I(N__24370));
    LocalMux I__3596 (
            .O(N__24370),
            .I(N__24366));
    InMux I__3595 (
            .O(N__24369),
            .I(N__24362));
    Span4Mux_v I__3594 (
            .O(N__24366),
            .I(N__24359));
    InMux I__3593 (
            .O(N__24365),
            .I(N__24356));
    LocalMux I__3592 (
            .O(N__24362),
            .I(measured_delay_hc_21));
    Odrv4 I__3591 (
            .O(N__24359),
            .I(measured_delay_hc_21));
    LocalMux I__3590 (
            .O(N__24356),
            .I(measured_delay_hc_21));
    InMux I__3589 (
            .O(N__24349),
            .I(N__24344));
    InMux I__3588 (
            .O(N__24348),
            .I(N__24341));
    InMux I__3587 (
            .O(N__24347),
            .I(N__24338));
    LocalMux I__3586 (
            .O(N__24344),
            .I(measured_delay_hc_20));
    LocalMux I__3585 (
            .O(N__24341),
            .I(measured_delay_hc_20));
    LocalMux I__3584 (
            .O(N__24338),
            .I(measured_delay_hc_20));
    CascadeMux I__3583 (
            .O(N__24331),
            .I(N__24326));
    CascadeMux I__3582 (
            .O(N__24330),
            .I(N__24323));
    InMux I__3581 (
            .O(N__24329),
            .I(N__24320));
    InMux I__3580 (
            .O(N__24326),
            .I(N__24317));
    InMux I__3579 (
            .O(N__24323),
            .I(N__24314));
    LocalMux I__3578 (
            .O(N__24320),
            .I(measured_delay_hc_22));
    LocalMux I__3577 (
            .O(N__24317),
            .I(measured_delay_hc_22));
    LocalMux I__3576 (
            .O(N__24314),
            .I(measured_delay_hc_22));
    InMux I__3575 (
            .O(N__24307),
            .I(N__24304));
    LocalMux I__3574 (
            .O(N__24304),
            .I(N__24301));
    Span12Mux_h I__3573 (
            .O(N__24301),
            .I(N__24298));
    Odrv12 I__3572 (
            .O(N__24298),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    InMux I__3571 (
            .O(N__24295),
            .I(N__24292));
    LocalMux I__3570 (
            .O(N__24292),
            .I(N__24289));
    Odrv4 I__3569 (
            .O(N__24289),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_2 ));
    CascadeMux I__3568 (
            .O(N__24286),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_ ));
    InMux I__3567 (
            .O(N__24283),
            .I(N__24280));
    LocalMux I__3566 (
            .O(N__24280),
            .I(\current_shift_inst.N_199 ));
    InMux I__3565 (
            .O(N__24277),
            .I(N__24274));
    LocalMux I__3564 (
            .O(N__24274),
            .I(N__24271));
    Span4Mux_v I__3563 (
            .O(N__24271),
            .I(N__24266));
    CascadeMux I__3562 (
            .O(N__24270),
            .I(N__24263));
    InMux I__3561 (
            .O(N__24269),
            .I(N__24259));
    Span4Mux_v I__3560 (
            .O(N__24266),
            .I(N__24256));
    InMux I__3559 (
            .O(N__24263),
            .I(N__24250));
    InMux I__3558 (
            .O(N__24262),
            .I(N__24250));
    LocalMux I__3557 (
            .O(N__24259),
            .I(N__24245));
    Span4Mux_h I__3556 (
            .O(N__24256),
            .I(N__24245));
    InMux I__3555 (
            .O(N__24255),
            .I(N__24242));
    LocalMux I__3554 (
            .O(N__24250),
            .I(\current_shift_inst.phase_validZ0 ));
    Odrv4 I__3553 (
            .O(N__24245),
            .I(\current_shift_inst.phase_validZ0 ));
    LocalMux I__3552 (
            .O(N__24242),
            .I(\current_shift_inst.phase_validZ0 ));
    CascadeMux I__3551 (
            .O(N__24235),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4_cascade_ ));
    InMux I__3550 (
            .O(N__24232),
            .I(N__24229));
    LocalMux I__3549 (
            .O(N__24229),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3 ));
    InMux I__3548 (
            .O(N__24226),
            .I(bfn_8_20_0_));
    InMux I__3547 (
            .O(N__24223),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ));
    InMux I__3546 (
            .O(N__24220),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    InMux I__3545 (
            .O(N__24217),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    InMux I__3544 (
            .O(N__24214),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    InMux I__3543 (
            .O(N__24211),
            .I(N__24208));
    LocalMux I__3542 (
            .O(N__24208),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__3541 (
            .O(N__24205),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    InMux I__3540 (
            .O(N__24202),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__3539 (
            .O(N__24199),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__3538 (
            .O(N__24196),
            .I(N__24193));
    LocalMux I__3537 (
            .O(N__24193),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__3536 (
            .O(N__24190),
            .I(bfn_8_19_0_));
    InMux I__3535 (
            .O(N__24187),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ));
    InMux I__3534 (
            .O(N__24184),
            .I(N__24180));
    InMux I__3533 (
            .O(N__24183),
            .I(N__24176));
    LocalMux I__3532 (
            .O(N__24180),
            .I(N__24173));
    CascadeMux I__3531 (
            .O(N__24179),
            .I(N__24170));
    LocalMux I__3530 (
            .O(N__24176),
            .I(N__24164));
    Span4Mux_h I__3529 (
            .O(N__24173),
            .I(N__24161));
    InMux I__3528 (
            .O(N__24170),
            .I(N__24156));
    InMux I__3527 (
            .O(N__24169),
            .I(N__24156));
    InMux I__3526 (
            .O(N__24168),
            .I(N__24153));
    InMux I__3525 (
            .O(N__24167),
            .I(N__24150));
    Odrv4 I__3524 (
            .O(N__24164),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__3523 (
            .O(N__24161),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__3522 (
            .O(N__24156),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__3521 (
            .O(N__24153),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__3520 (
            .O(N__24150),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__3519 (
            .O(N__24139),
            .I(N__24136));
    LocalMux I__3518 (
            .O(N__24136),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__3517 (
            .O(N__24133),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__3516 (
            .O(N__24130),
            .I(N__24127));
    InMux I__3515 (
            .O(N__24127),
            .I(N__24124));
    LocalMux I__3514 (
            .O(N__24124),
            .I(N__24121));
    Odrv4 I__3513 (
            .O(N__24121),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__3512 (
            .O(N__24118),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    InMux I__3511 (
            .O(N__24115),
            .I(N__24112));
    LocalMux I__3510 (
            .O(N__24112),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__3509 (
            .O(N__24109),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    InMux I__3508 (
            .O(N__24106),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    InMux I__3507 (
            .O(N__24103),
            .I(N__24100));
    LocalMux I__3506 (
            .O(N__24100),
            .I(N__24097));
    Odrv4 I__3505 (
            .O(N__24097),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__3504 (
            .O(N__24094),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    InMux I__3503 (
            .O(N__24091),
            .I(N__24088));
    LocalMux I__3502 (
            .O(N__24088),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__3501 (
            .O(N__24085),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    InMux I__3500 (
            .O(N__24082),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    InMux I__3499 (
            .O(N__24079),
            .I(N__24074));
    InMux I__3498 (
            .O(N__24078),
            .I(N__24068));
    InMux I__3497 (
            .O(N__24077),
            .I(N__24068));
    LocalMux I__3496 (
            .O(N__24074),
            .I(N__24065));
    InMux I__3495 (
            .O(N__24073),
            .I(N__24062));
    LocalMux I__3494 (
            .O(N__24068),
            .I(N__24059));
    Span4Mux_h I__3493 (
            .O(N__24065),
            .I(N__24054));
    LocalMux I__3492 (
            .O(N__24062),
            .I(N__24054));
    Span4Mux_h I__3491 (
            .O(N__24059),
            .I(N__24051));
    Odrv4 I__3490 (
            .O(N__24054),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__3489 (
            .O(N__24051),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__3488 (
            .O(N__24046),
            .I(N__24043));
    LocalMux I__3487 (
            .O(N__24043),
            .I(N__24040));
    Odrv4 I__3486 (
            .O(N__24040),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__3485 (
            .O(N__24037),
            .I(bfn_8_18_0_));
    InMux I__3484 (
            .O(N__24034),
            .I(N__24029));
    InMux I__3483 (
            .O(N__24033),
            .I(N__24024));
    InMux I__3482 (
            .O(N__24032),
            .I(N__24024));
    LocalMux I__3481 (
            .O(N__24029),
            .I(N__24021));
    LocalMux I__3480 (
            .O(N__24024),
            .I(N__24017));
    Span4Mux_h I__3479 (
            .O(N__24021),
            .I(N__24014));
    InMux I__3478 (
            .O(N__24020),
            .I(N__24011));
    Span4Mux_h I__3477 (
            .O(N__24017),
            .I(N__24008));
    Odrv4 I__3476 (
            .O(N__24014),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__3475 (
            .O(N__24011),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__3474 (
            .O(N__24008),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__3473 (
            .O(N__24001),
            .I(N__23998));
    LocalMux I__3472 (
            .O(N__23998),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__3471 (
            .O(N__23995),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ));
    InMux I__3470 (
            .O(N__23992),
            .I(N__23989));
    LocalMux I__3469 (
            .O(N__23989),
            .I(N__23986));
    Odrv4 I__3468 (
            .O(N__23986),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__3467 (
            .O(N__23983),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    InMux I__3466 (
            .O(N__23980),
            .I(N__23977));
    LocalMux I__3465 (
            .O(N__23977),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__3464 (
            .O(N__23974),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    InMux I__3463 (
            .O(N__23971),
            .I(N__23968));
    LocalMux I__3462 (
            .O(N__23968),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__3461 (
            .O(N__23965),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    InMux I__3460 (
            .O(N__23962),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    InMux I__3459 (
            .O(N__23959),
            .I(N__23956));
    LocalMux I__3458 (
            .O(N__23956),
            .I(N__23953));
    Odrv4 I__3457 (
            .O(N__23953),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__3456 (
            .O(N__23950),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    InMux I__3455 (
            .O(N__23947),
            .I(N__23944));
    LocalMux I__3454 (
            .O(N__23944),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__3453 (
            .O(N__23941),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    InMux I__3452 (
            .O(N__23938),
            .I(N__23934));
    InMux I__3451 (
            .O(N__23937),
            .I(N__23931));
    LocalMux I__3450 (
            .O(N__23934),
            .I(N__23925));
    LocalMux I__3449 (
            .O(N__23931),
            .I(N__23925));
    InMux I__3448 (
            .O(N__23930),
            .I(N__23922));
    Span4Mux_h I__3447 (
            .O(N__23925),
            .I(N__23919));
    LocalMux I__3446 (
            .O(N__23922),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    Odrv4 I__3445 (
            .O(N__23919),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    InMux I__3444 (
            .O(N__23914),
            .I(N__23909));
    InMux I__3443 (
            .O(N__23913),
            .I(N__23906));
    InMux I__3442 (
            .O(N__23912),
            .I(N__23903));
    LocalMux I__3441 (
            .O(N__23909),
            .I(N__23898));
    LocalMux I__3440 (
            .O(N__23906),
            .I(N__23898));
    LocalMux I__3439 (
            .O(N__23903),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv12 I__3438 (
            .O(N__23898),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__3437 (
            .O(N__23893),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ));
    CascadeMux I__3436 (
            .O(N__23890),
            .I(N__23886));
    InMux I__3435 (
            .O(N__23889),
            .I(N__23882));
    InMux I__3434 (
            .O(N__23886),
            .I(N__23879));
    InMux I__3433 (
            .O(N__23885),
            .I(N__23876));
    LocalMux I__3432 (
            .O(N__23882),
            .I(N__23871));
    LocalMux I__3431 (
            .O(N__23879),
            .I(N__23871));
    LocalMux I__3430 (
            .O(N__23876),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv12 I__3429 (
            .O(N__23871),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__3428 (
            .O(N__23866),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    InMux I__3427 (
            .O(N__23863),
            .I(N__23857));
    InMux I__3426 (
            .O(N__23862),
            .I(N__23850));
    InMux I__3425 (
            .O(N__23861),
            .I(N__23850));
    InMux I__3424 (
            .O(N__23860),
            .I(N__23850));
    LocalMux I__3423 (
            .O(N__23857),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    LocalMux I__3422 (
            .O(N__23850),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    InMux I__3421 (
            .O(N__23845),
            .I(N__23839));
    InMux I__3420 (
            .O(N__23844),
            .I(N__23834));
    InMux I__3419 (
            .O(N__23843),
            .I(N__23834));
    InMux I__3418 (
            .O(N__23842),
            .I(N__23831));
    LocalMux I__3417 (
            .O(N__23839),
            .I(N__23826));
    LocalMux I__3416 (
            .O(N__23834),
            .I(N__23826));
    LocalMux I__3415 (
            .O(N__23831),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv12 I__3414 (
            .O(N__23826),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__3413 (
            .O(N__23821),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CascadeMux I__3412 (
            .O(N__23818),
            .I(N__23813));
    InMux I__3411 (
            .O(N__23817),
            .I(N__23808));
    InMux I__3410 (
            .O(N__23816),
            .I(N__23808));
    InMux I__3409 (
            .O(N__23813),
            .I(N__23805));
    LocalMux I__3408 (
            .O(N__23808),
            .I(N__23800));
    LocalMux I__3407 (
            .O(N__23805),
            .I(N__23800));
    Span4Mux_h I__3406 (
            .O(N__23800),
            .I(N__23797));
    Span4Mux_h I__3405 (
            .O(N__23797),
            .I(N__23793));
    InMux I__3404 (
            .O(N__23796),
            .I(N__23790));
    Odrv4 I__3403 (
            .O(N__23793),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__3402 (
            .O(N__23790),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__3401 (
            .O(N__23785),
            .I(N__23782));
    InMux I__3400 (
            .O(N__23782),
            .I(N__23779));
    LocalMux I__3399 (
            .O(N__23779),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__3398 (
            .O(N__23776),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    InMux I__3397 (
            .O(N__23773),
            .I(N__23770));
    LocalMux I__3396 (
            .O(N__23770),
            .I(N__23766));
    InMux I__3395 (
            .O(N__23769),
            .I(N__23761));
    Span4Mux_h I__3394 (
            .O(N__23766),
            .I(N__23758));
    InMux I__3393 (
            .O(N__23765),
            .I(N__23753));
    InMux I__3392 (
            .O(N__23764),
            .I(N__23753));
    LocalMux I__3391 (
            .O(N__23761),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__3390 (
            .O(N__23758),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__3389 (
            .O(N__23753),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__3388 (
            .O(N__23746),
            .I(N__23743));
    LocalMux I__3387 (
            .O(N__23743),
            .I(N__23740));
    Span4Mux_h I__3386 (
            .O(N__23740),
            .I(N__23737));
    Odrv4 I__3385 (
            .O(N__23737),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__3384 (
            .O(N__23734),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    InMux I__3383 (
            .O(N__23731),
            .I(N__23726));
    InMux I__3382 (
            .O(N__23730),
            .I(N__23721));
    InMux I__3381 (
            .O(N__23729),
            .I(N__23721));
    LocalMux I__3380 (
            .O(N__23726),
            .I(N__23715));
    LocalMux I__3379 (
            .O(N__23721),
            .I(N__23715));
    InMux I__3378 (
            .O(N__23720),
            .I(N__23712));
    Span4Mux_h I__3377 (
            .O(N__23715),
            .I(N__23709));
    LocalMux I__3376 (
            .O(N__23712),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__3375 (
            .O(N__23709),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__3374 (
            .O(N__23704),
            .I(N__23701));
    LocalMux I__3373 (
            .O(N__23701),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__3372 (
            .O(N__23698),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    InMux I__3371 (
            .O(N__23695),
            .I(N__23691));
    CascadeMux I__3370 (
            .O(N__23694),
            .I(N__23687));
    LocalMux I__3369 (
            .O(N__23691),
            .I(N__23684));
    InMux I__3368 (
            .O(N__23690),
            .I(N__23679));
    InMux I__3367 (
            .O(N__23687),
            .I(N__23679));
    Span4Mux_h I__3366 (
            .O(N__23684),
            .I(N__23673));
    LocalMux I__3365 (
            .O(N__23679),
            .I(N__23673));
    InMux I__3364 (
            .O(N__23678),
            .I(N__23670));
    Span4Mux_h I__3363 (
            .O(N__23673),
            .I(N__23667));
    LocalMux I__3362 (
            .O(N__23670),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__3361 (
            .O(N__23667),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__3360 (
            .O(N__23662),
            .I(N__23659));
    LocalMux I__3359 (
            .O(N__23659),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    CascadeMux I__3358 (
            .O(N__23656),
            .I(\phase_controller_inst1.N_228_cascade_ ));
    InMux I__3357 (
            .O(N__23653),
            .I(N__23650));
    LocalMux I__3356 (
            .O(N__23650),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ));
    InMux I__3355 (
            .O(N__23647),
            .I(N__23643));
    InMux I__3354 (
            .O(N__23646),
            .I(N__23640));
    LocalMux I__3353 (
            .O(N__23643),
            .I(N__23637));
    LocalMux I__3352 (
            .O(N__23640),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__3351 (
            .O(N__23637),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__3350 (
            .O(N__23632),
            .I(N__23622));
    CascadeMux I__3349 (
            .O(N__23631),
            .I(N__23618));
    CascadeMux I__3348 (
            .O(N__23630),
            .I(N__23614));
    CascadeMux I__3347 (
            .O(N__23629),
            .I(N__23610));
    CascadeMux I__3346 (
            .O(N__23628),
            .I(N__23606));
    CascadeMux I__3345 (
            .O(N__23627),
            .I(N__23601));
    CascadeMux I__3344 (
            .O(N__23626),
            .I(N__23598));
    CascadeMux I__3343 (
            .O(N__23625),
            .I(N__23594));
    InMux I__3342 (
            .O(N__23622),
            .I(N__23579));
    InMux I__3341 (
            .O(N__23621),
            .I(N__23579));
    InMux I__3340 (
            .O(N__23618),
            .I(N__23579));
    InMux I__3339 (
            .O(N__23617),
            .I(N__23579));
    InMux I__3338 (
            .O(N__23614),
            .I(N__23579));
    InMux I__3337 (
            .O(N__23613),
            .I(N__23579));
    InMux I__3336 (
            .O(N__23610),
            .I(N__23579));
    InMux I__3335 (
            .O(N__23609),
            .I(N__23560));
    InMux I__3334 (
            .O(N__23606),
            .I(N__23560));
    InMux I__3333 (
            .O(N__23605),
            .I(N__23560));
    InMux I__3332 (
            .O(N__23604),
            .I(N__23560));
    InMux I__3331 (
            .O(N__23601),
            .I(N__23560));
    InMux I__3330 (
            .O(N__23598),
            .I(N__23560));
    InMux I__3329 (
            .O(N__23597),
            .I(N__23560));
    InMux I__3328 (
            .O(N__23594),
            .I(N__23560));
    LocalMux I__3327 (
            .O(N__23579),
            .I(N__23557));
    CascadeMux I__3326 (
            .O(N__23578),
            .I(N__23553));
    CascadeMux I__3325 (
            .O(N__23577),
            .I(N__23547));
    LocalMux I__3324 (
            .O(N__23560),
            .I(N__23544));
    Span4Mux_v I__3323 (
            .O(N__23557),
            .I(N__23541));
    InMux I__3322 (
            .O(N__23556),
            .I(N__23532));
    InMux I__3321 (
            .O(N__23553),
            .I(N__23532));
    InMux I__3320 (
            .O(N__23552),
            .I(N__23532));
    InMux I__3319 (
            .O(N__23551),
            .I(N__23532));
    InMux I__3318 (
            .O(N__23550),
            .I(N__23524));
    InMux I__3317 (
            .O(N__23547),
            .I(N__23524));
    Span4Mux_h I__3316 (
            .O(N__23544),
            .I(N__23517));
    Span4Mux_h I__3315 (
            .O(N__23541),
            .I(N__23517));
    LocalMux I__3314 (
            .O(N__23532),
            .I(N__23517));
    InMux I__3313 (
            .O(N__23531),
            .I(N__23510));
    InMux I__3312 (
            .O(N__23530),
            .I(N__23510));
    InMux I__3311 (
            .O(N__23529),
            .I(N__23510));
    LocalMux I__3310 (
            .O(N__23524),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__3309 (
            .O(N__23517),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__3308 (
            .O(N__23510),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    CascadeMux I__3307 (
            .O(N__23503),
            .I(N__23489));
    CascadeMux I__3306 (
            .O(N__23502),
            .I(N__23485));
    InMux I__3305 (
            .O(N__23501),
            .I(N__23466));
    InMux I__3304 (
            .O(N__23500),
            .I(N__23466));
    InMux I__3303 (
            .O(N__23499),
            .I(N__23466));
    InMux I__3302 (
            .O(N__23498),
            .I(N__23466));
    InMux I__3301 (
            .O(N__23497),
            .I(N__23466));
    InMux I__3300 (
            .O(N__23496),
            .I(N__23466));
    InMux I__3299 (
            .O(N__23495),
            .I(N__23466));
    InMux I__3298 (
            .O(N__23494),
            .I(N__23466));
    InMux I__3297 (
            .O(N__23493),
            .I(N__23461));
    InMux I__3296 (
            .O(N__23492),
            .I(N__23448));
    InMux I__3295 (
            .O(N__23489),
            .I(N__23448));
    InMux I__3294 (
            .O(N__23488),
            .I(N__23448));
    InMux I__3293 (
            .O(N__23485),
            .I(N__23448));
    InMux I__3292 (
            .O(N__23484),
            .I(N__23448));
    InMux I__3291 (
            .O(N__23483),
            .I(N__23448));
    LocalMux I__3290 (
            .O(N__23466),
            .I(N__23445));
    InMux I__3289 (
            .O(N__23465),
            .I(N__23433));
    InMux I__3288 (
            .O(N__23464),
            .I(N__23433));
    LocalMux I__3287 (
            .O(N__23461),
            .I(N__23428));
    LocalMux I__3286 (
            .O(N__23448),
            .I(N__23428));
    Span4Mux_h I__3285 (
            .O(N__23445),
            .I(N__23425));
    InMux I__3284 (
            .O(N__23444),
            .I(N__23420));
    InMux I__3283 (
            .O(N__23443),
            .I(N__23420));
    InMux I__3282 (
            .O(N__23442),
            .I(N__23411));
    InMux I__3281 (
            .O(N__23441),
            .I(N__23411));
    InMux I__3280 (
            .O(N__23440),
            .I(N__23411));
    InMux I__3279 (
            .O(N__23439),
            .I(N__23411));
    InMux I__3278 (
            .O(N__23438),
            .I(N__23408));
    LocalMux I__3277 (
            .O(N__23433),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv12 I__3276 (
            .O(N__23428),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__3275 (
            .O(N__23425),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__3274 (
            .O(N__23420),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__3273 (
            .O(N__23411),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__3272 (
            .O(N__23408),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__3271 (
            .O(N__23395),
            .I(N__23388));
    CascadeMux I__3270 (
            .O(N__23394),
            .I(N__23385));
    CascadeMux I__3269 (
            .O(N__23393),
            .I(N__23382));
    CascadeMux I__3268 (
            .O(N__23392),
            .I(N__23379));
    CascadeMux I__3267 (
            .O(N__23391),
            .I(N__23371));
    InMux I__3266 (
            .O(N__23388),
            .I(N__23356));
    InMux I__3265 (
            .O(N__23385),
            .I(N__23356));
    InMux I__3264 (
            .O(N__23382),
            .I(N__23356));
    InMux I__3263 (
            .O(N__23379),
            .I(N__23356));
    InMux I__3262 (
            .O(N__23378),
            .I(N__23347));
    InMux I__3261 (
            .O(N__23377),
            .I(N__23347));
    InMux I__3260 (
            .O(N__23376),
            .I(N__23347));
    InMux I__3259 (
            .O(N__23375),
            .I(N__23347));
    CascadeMux I__3258 (
            .O(N__23374),
            .I(N__23341));
    InMux I__3257 (
            .O(N__23371),
            .I(N__23332));
    InMux I__3256 (
            .O(N__23370),
            .I(N__23332));
    InMux I__3255 (
            .O(N__23369),
            .I(N__23332));
    InMux I__3254 (
            .O(N__23368),
            .I(N__23323));
    InMux I__3253 (
            .O(N__23367),
            .I(N__23323));
    InMux I__3252 (
            .O(N__23366),
            .I(N__23323));
    InMux I__3251 (
            .O(N__23365),
            .I(N__23323));
    LocalMux I__3250 (
            .O(N__23356),
            .I(N__23318));
    LocalMux I__3249 (
            .O(N__23347),
            .I(N__23318));
    CascadeMux I__3248 (
            .O(N__23346),
            .I(N__23315));
    CascadeMux I__3247 (
            .O(N__23345),
            .I(N__23311));
    CascadeMux I__3246 (
            .O(N__23344),
            .I(N__23308));
    InMux I__3245 (
            .O(N__23341),
            .I(N__23301));
    InMux I__3244 (
            .O(N__23340),
            .I(N__23301));
    InMux I__3243 (
            .O(N__23339),
            .I(N__23298));
    LocalMux I__3242 (
            .O(N__23332),
            .I(N__23293));
    LocalMux I__3241 (
            .O(N__23323),
            .I(N__23293));
    Span4Mux_h I__3240 (
            .O(N__23318),
            .I(N__23290));
    InMux I__3239 (
            .O(N__23315),
            .I(N__23285));
    InMux I__3238 (
            .O(N__23314),
            .I(N__23285));
    InMux I__3237 (
            .O(N__23311),
            .I(N__23278));
    InMux I__3236 (
            .O(N__23308),
            .I(N__23278));
    InMux I__3235 (
            .O(N__23307),
            .I(N__23278));
    InMux I__3234 (
            .O(N__23306),
            .I(N__23275));
    LocalMux I__3233 (
            .O(N__23301),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__3232 (
            .O(N__23298),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv12 I__3231 (
            .O(N__23293),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__3230 (
            .O(N__23290),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__3229 (
            .O(N__23285),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__3228 (
            .O(N__23278),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__3227 (
            .O(N__23275),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    InMux I__3226 (
            .O(N__23260),
            .I(N__23257));
    LocalMux I__3225 (
            .O(N__23257),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ));
    InMux I__3224 (
            .O(N__23254),
            .I(N__23251));
    LocalMux I__3223 (
            .O(N__23251),
            .I(N__23247));
    InMux I__3222 (
            .O(N__23250),
            .I(N__23244));
    Span4Mux_h I__3221 (
            .O(N__23247),
            .I(N__23241));
    LocalMux I__3220 (
            .O(N__23244),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__3219 (
            .O(N__23241),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__3218 (
            .O(N__23236),
            .I(N__23233));
    LocalMux I__3217 (
            .O(N__23233),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ));
    InMux I__3216 (
            .O(N__23230),
            .I(N__23226));
    InMux I__3215 (
            .O(N__23229),
            .I(N__23223));
    LocalMux I__3214 (
            .O(N__23226),
            .I(N__23220));
    LocalMux I__3213 (
            .O(N__23223),
            .I(N__23217));
    Span4Mux_h I__3212 (
            .O(N__23220),
            .I(N__23214));
    Odrv4 I__3211 (
            .O(N__23217),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__3210 (
            .O(N__23214),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__3209 (
            .O(N__23209),
            .I(N__23206));
    LocalMux I__3208 (
            .O(N__23206),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ));
    InMux I__3207 (
            .O(N__23203),
            .I(N__23200));
    LocalMux I__3206 (
            .O(N__23200),
            .I(N__23196));
    InMux I__3205 (
            .O(N__23199),
            .I(N__23193));
    Span4Mux_h I__3204 (
            .O(N__23196),
            .I(N__23190));
    LocalMux I__3203 (
            .O(N__23193),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__3202 (
            .O(N__23190),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__3201 (
            .O(N__23185),
            .I(N__23182));
    LocalMux I__3200 (
            .O(N__23182),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ));
    InMux I__3199 (
            .O(N__23179),
            .I(N__23176));
    LocalMux I__3198 (
            .O(N__23176),
            .I(N__23173));
    Span4Mux_h I__3197 (
            .O(N__23173),
            .I(N__23170));
    Span4Mux_h I__3196 (
            .O(N__23170),
            .I(N__23167));
    Odrv4 I__3195 (
            .O(N__23167),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    InMux I__3194 (
            .O(N__23164),
            .I(N__23161));
    LocalMux I__3193 (
            .O(N__23161),
            .I(N__23158));
    Span4Mux_h I__3192 (
            .O(N__23158),
            .I(N__23155));
    Span4Mux_h I__3191 (
            .O(N__23155),
            .I(N__23152));
    Odrv4 I__3190 (
            .O(N__23152),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    InMux I__3189 (
            .O(N__23149),
            .I(N__23146));
    LocalMux I__3188 (
            .O(N__23146),
            .I(N__23143));
    Span4Mux_v I__3187 (
            .O(N__23143),
            .I(N__23140));
    Span4Mux_h I__3186 (
            .O(N__23140),
            .I(N__23137));
    Odrv4 I__3185 (
            .O(N__23137),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__3184 (
            .O(N__23134),
            .I(N__23131));
    InMux I__3183 (
            .O(N__23131),
            .I(N__23128));
    LocalMux I__3182 (
            .O(N__23128),
            .I(N__23125));
    Span4Mux_v I__3181 (
            .O(N__23125),
            .I(N__23122));
    Odrv4 I__3180 (
            .O(N__23122),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__3179 (
            .O(N__23119),
            .I(N__23116));
    InMux I__3178 (
            .O(N__23116),
            .I(N__23113));
    LocalMux I__3177 (
            .O(N__23113),
            .I(N__23110));
    Span4Mux_v I__3176 (
            .O(N__23110),
            .I(N__23107));
    Odrv4 I__3175 (
            .O(N__23107),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__3174 (
            .O(N__23104),
            .I(N__23101));
    InMux I__3173 (
            .O(N__23101),
            .I(N__23098));
    LocalMux I__3172 (
            .O(N__23098),
            .I(N__23095));
    Span4Mux_h I__3171 (
            .O(N__23095),
            .I(N__23092));
    Odrv4 I__3170 (
            .O(N__23092),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__3169 (
            .O(N__23089),
            .I(N__23086));
    InMux I__3168 (
            .O(N__23086),
            .I(N__23083));
    LocalMux I__3167 (
            .O(N__23083),
            .I(N__23080));
    Span4Mux_v I__3166 (
            .O(N__23080),
            .I(N__23077));
    Span4Mux_h I__3165 (
            .O(N__23077),
            .I(N__23074));
    Odrv4 I__3164 (
            .O(N__23074),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__3163 (
            .O(N__23071),
            .I(N__23068));
    InMux I__3162 (
            .O(N__23068),
            .I(N__23065));
    LocalMux I__3161 (
            .O(N__23065),
            .I(N__23062));
    Span4Mux_h I__3160 (
            .O(N__23062),
            .I(N__23059));
    Odrv4 I__3159 (
            .O(N__23059),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    IoInMux I__3158 (
            .O(N__23056),
            .I(N__23053));
    LocalMux I__3157 (
            .O(N__23053),
            .I(N__23050));
    IoSpan4Mux I__3156 (
            .O(N__23050),
            .I(N__23047));
    Span4Mux_s2_v I__3155 (
            .O(N__23047),
            .I(N__23044));
    Span4Mux_v I__3154 (
            .O(N__23044),
            .I(N__23041));
    Odrv4 I__3153 (
            .O(N__23041),
            .I(\current_shift_inst.timer_s1.N_187_i ));
    InMux I__3152 (
            .O(N__23038),
            .I(N__23035));
    LocalMux I__3151 (
            .O(N__23035),
            .I(N__23032));
    Odrv12 I__3150 (
            .O(N__23032),
            .I(il_max_comp1_c));
    InMux I__3149 (
            .O(N__23029),
            .I(N__23026));
    LocalMux I__3148 (
            .O(N__23026),
            .I(N__23023));
    Odrv12 I__3147 (
            .O(N__23023),
            .I(il_max_comp1_D1));
    InMux I__3146 (
            .O(N__23020),
            .I(N__23017));
    LocalMux I__3145 (
            .O(N__23017),
            .I(N__23014));
    Odrv12 I__3144 (
            .O(N__23014),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__3143 (
            .O(N__23011),
            .I(N__23008));
    LocalMux I__3142 (
            .O(N__23008),
            .I(N__23005));
    Odrv12 I__3141 (
            .O(N__23005),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    CascadeMux I__3140 (
            .O(N__23002),
            .I(N__22999));
    InMux I__3139 (
            .O(N__22999),
            .I(N__22996));
    LocalMux I__3138 (
            .O(N__22996),
            .I(N__22993));
    Span4Mux_v I__3137 (
            .O(N__22993),
            .I(N__22990));
    Span4Mux_h I__3136 (
            .O(N__22990),
            .I(N__22987));
    Odrv4 I__3135 (
            .O(N__22987),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__3134 (
            .O(N__22984),
            .I(N__22981));
    InMux I__3133 (
            .O(N__22981),
            .I(N__22978));
    LocalMux I__3132 (
            .O(N__22978),
            .I(N__22975));
    Span4Mux_h I__3131 (
            .O(N__22975),
            .I(N__22972));
    Odrv4 I__3130 (
            .O(N__22972),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    CascadeMux I__3129 (
            .O(N__22969),
            .I(N__22966));
    InMux I__3128 (
            .O(N__22966),
            .I(N__22963));
    LocalMux I__3127 (
            .O(N__22963),
            .I(N__22960));
    Span4Mux_v I__3126 (
            .O(N__22960),
            .I(N__22957));
    Odrv4 I__3125 (
            .O(N__22957),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__3124 (
            .O(N__22954),
            .I(N__22951));
    InMux I__3123 (
            .O(N__22951),
            .I(N__22948));
    LocalMux I__3122 (
            .O(N__22948),
            .I(N__22945));
    Span4Mux_h I__3121 (
            .O(N__22945),
            .I(N__22942));
    Odrv4 I__3120 (
            .O(N__22942),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    CascadeMux I__3119 (
            .O(N__22939),
            .I(N__22936));
    InMux I__3118 (
            .O(N__22936),
            .I(N__22933));
    LocalMux I__3117 (
            .O(N__22933),
            .I(N__22930));
    Span4Mux_h I__3116 (
            .O(N__22930),
            .I(N__22927));
    Odrv4 I__3115 (
            .O(N__22927),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__3114 (
            .O(N__22924),
            .I(N__22921));
    LocalMux I__3113 (
            .O(N__22921),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31 ));
    InMux I__3112 (
            .O(N__22918),
            .I(N__22915));
    LocalMux I__3111 (
            .O(N__22915),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2 ));
    InMux I__3110 (
            .O(N__22912),
            .I(N__22909));
    LocalMux I__3109 (
            .O(N__22909),
            .I(N__22905));
    InMux I__3108 (
            .O(N__22908),
            .I(N__22902));
    Span4Mux_v I__3107 (
            .O(N__22905),
            .I(N__22897));
    LocalMux I__3106 (
            .O(N__22902),
            .I(N__22897));
    Odrv4 I__3105 (
            .O(N__22897),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    CascadeMux I__3104 (
            .O(N__22894),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_ ));
    InMux I__3103 (
            .O(N__22891),
            .I(N__22885));
    InMux I__3102 (
            .O(N__22890),
            .I(N__22885));
    LocalMux I__3101 (
            .O(N__22885),
            .I(N__22882));
    Odrv4 I__3100 (
            .O(N__22882),
            .I(\current_shift_inst.PI_CTRL.N_44 ));
    InMux I__3099 (
            .O(N__22879),
            .I(N__22876));
    LocalMux I__3098 (
            .O(N__22876),
            .I(N__22872));
    InMux I__3097 (
            .O(N__22875),
            .I(N__22869));
    Span4Mux_v I__3096 (
            .O(N__22872),
            .I(N__22866));
    LocalMux I__3095 (
            .O(N__22869),
            .I(N__22863));
    Odrv4 I__3094 (
            .O(N__22866),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv12 I__3093 (
            .O(N__22863),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__3092 (
            .O(N__22858),
            .I(N__22855));
    LocalMux I__3091 (
            .O(N__22855),
            .I(N__22852));
    Span4Mux_h I__3090 (
            .O(N__22852),
            .I(N__22849));
    Odrv4 I__3089 (
            .O(N__22849),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ));
    InMux I__3088 (
            .O(N__22846),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__3087 (
            .O(N__22843),
            .I(N__22840));
    LocalMux I__3086 (
            .O(N__22840),
            .I(N__22836));
    InMux I__3085 (
            .O(N__22839),
            .I(N__22833));
    Span4Mux_h I__3084 (
            .O(N__22836),
            .I(N__22828));
    LocalMux I__3083 (
            .O(N__22833),
            .I(N__22828));
    Odrv4 I__3082 (
            .O(N__22828),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__3081 (
            .O(N__22825),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__3080 (
            .O(N__22822),
            .I(N__22819));
    LocalMux I__3079 (
            .O(N__22819),
            .I(N__22816));
    Span4Mux_h I__3078 (
            .O(N__22816),
            .I(N__22813));
    Odrv4 I__3077 (
            .O(N__22813),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ));
    InMux I__3076 (
            .O(N__22810),
            .I(N__22807));
    LocalMux I__3075 (
            .O(N__22807),
            .I(N__22804));
    Odrv4 I__3074 (
            .O(N__22804),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    CascadeMux I__3073 (
            .O(N__22801),
            .I(\current_shift_inst.PI_CTRL.N_47_16_cascade_ ));
    InMux I__3072 (
            .O(N__22798),
            .I(N__22795));
    LocalMux I__3071 (
            .O(N__22795),
            .I(N__22792));
    Odrv12 I__3070 (
            .O(N__22792),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31 ));
    InMux I__3069 (
            .O(N__22789),
            .I(N__22786));
    LocalMux I__3068 (
            .O(N__22786),
            .I(\current_shift_inst.PI_CTRL.N_47_21 ));
    InMux I__3067 (
            .O(N__22783),
            .I(N__22780));
    LocalMux I__3066 (
            .O(N__22780),
            .I(\current_shift_inst.PI_CTRL.N_47_16 ));
    CascadeMux I__3065 (
            .O(N__22777),
            .I(\current_shift_inst.PI_CTRL.N_47_21_cascade_ ));
    InMux I__3064 (
            .O(N__22774),
            .I(N__22771));
    LocalMux I__3063 (
            .O(N__22771),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31 ));
    InMux I__3062 (
            .O(N__22768),
            .I(N__22765));
    LocalMux I__3061 (
            .O(N__22765),
            .I(N__22761));
    InMux I__3060 (
            .O(N__22764),
            .I(N__22758));
    Odrv4 I__3059 (
            .O(N__22761),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__3058 (
            .O(N__22758),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__3057 (
            .O(N__22753),
            .I(N__22750));
    LocalMux I__3056 (
            .O(N__22750),
            .I(N__22747));
    Odrv12 I__3055 (
            .O(N__22747),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ));
    InMux I__3054 (
            .O(N__22744),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__3053 (
            .O(N__22741),
            .I(N__22738));
    LocalMux I__3052 (
            .O(N__22738),
            .I(N__22734));
    InMux I__3051 (
            .O(N__22737),
            .I(N__22731));
    Odrv4 I__3050 (
            .O(N__22734),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__3049 (
            .O(N__22731),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__3048 (
            .O(N__22726),
            .I(N__22723));
    LocalMux I__3047 (
            .O(N__22723),
            .I(N__22720));
    Odrv4 I__3046 (
            .O(N__22720),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ));
    InMux I__3045 (
            .O(N__22717),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__3044 (
            .O(N__22714),
            .I(N__22711));
    LocalMux I__3043 (
            .O(N__22711),
            .I(N__22707));
    InMux I__3042 (
            .O(N__22710),
            .I(N__22704));
    Odrv4 I__3041 (
            .O(N__22707),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__3040 (
            .O(N__22704),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__3039 (
            .O(N__22699),
            .I(N__22696));
    LocalMux I__3038 (
            .O(N__22696),
            .I(N__22693));
    Odrv4 I__3037 (
            .O(N__22693),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ));
    InMux I__3036 (
            .O(N__22690),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__3035 (
            .O(N__22687),
            .I(N__22683));
    InMux I__3034 (
            .O(N__22686),
            .I(N__22680));
    LocalMux I__3033 (
            .O(N__22683),
            .I(N__22677));
    LocalMux I__3032 (
            .O(N__22680),
            .I(N__22674));
    Odrv4 I__3031 (
            .O(N__22677),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__3030 (
            .O(N__22674),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__3029 (
            .O(N__22669),
            .I(N__22666));
    LocalMux I__3028 (
            .O(N__22666),
            .I(N__22663));
    Odrv4 I__3027 (
            .O(N__22663),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ));
    InMux I__3026 (
            .O(N__22660),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__3025 (
            .O(N__22657),
            .I(N__22654));
    LocalMux I__3024 (
            .O(N__22654),
            .I(N__22650));
    InMux I__3023 (
            .O(N__22653),
            .I(N__22647));
    Odrv12 I__3022 (
            .O(N__22650),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__3021 (
            .O(N__22647),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__3020 (
            .O(N__22642),
            .I(N__22639));
    LocalMux I__3019 (
            .O(N__22639),
            .I(N__22636));
    Odrv4 I__3018 (
            .O(N__22636),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ));
    InMux I__3017 (
            .O(N__22633),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__3016 (
            .O(N__22630),
            .I(N__22627));
    LocalMux I__3015 (
            .O(N__22627),
            .I(N__22624));
    Span4Mux_h I__3014 (
            .O(N__22624),
            .I(N__22620));
    InMux I__3013 (
            .O(N__22623),
            .I(N__22617));
    Odrv4 I__3012 (
            .O(N__22620),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__3011 (
            .O(N__22617),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__3010 (
            .O(N__22612),
            .I(N__22609));
    LocalMux I__3009 (
            .O(N__22609),
            .I(N__22606));
    Odrv4 I__3008 (
            .O(N__22606),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ));
    InMux I__3007 (
            .O(N__22603),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__3006 (
            .O(N__22600),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__3005 (
            .O(N__22597),
            .I(N__22594));
    LocalMux I__3004 (
            .O(N__22594),
            .I(N__22590));
    InMux I__3003 (
            .O(N__22593),
            .I(N__22587));
    Span4Mux_v I__3002 (
            .O(N__22590),
            .I(N__22584));
    LocalMux I__3001 (
            .O(N__22587),
            .I(N__22581));
    Odrv4 I__3000 (
            .O(N__22584),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv12 I__2999 (
            .O(N__22581),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__2998 (
            .O(N__22576),
            .I(N__22573));
    LocalMux I__2997 (
            .O(N__22573),
            .I(N__22570));
    Span4Mux_h I__2996 (
            .O(N__22570),
            .I(N__22567));
    Odrv4 I__2995 (
            .O(N__22567),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ));
    InMux I__2994 (
            .O(N__22564),
            .I(bfn_7_15_0_));
    InMux I__2993 (
            .O(N__22561),
            .I(N__22558));
    LocalMux I__2992 (
            .O(N__22558),
            .I(N__22555));
    Span4Mux_h I__2991 (
            .O(N__22555),
            .I(N__22551));
    InMux I__2990 (
            .O(N__22554),
            .I(N__22548));
    Odrv4 I__2989 (
            .O(N__22551),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__2988 (
            .O(N__22548),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__2987 (
            .O(N__22543),
            .I(N__22540));
    LocalMux I__2986 (
            .O(N__22540),
            .I(N__22537));
    Span4Mux_v I__2985 (
            .O(N__22537),
            .I(N__22534));
    Odrv4 I__2984 (
            .O(N__22534),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ));
    InMux I__2983 (
            .O(N__22531),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    CascadeMux I__2982 (
            .O(N__22528),
            .I(N__22525));
    InMux I__2981 (
            .O(N__22525),
            .I(N__22522));
    LocalMux I__2980 (
            .O(N__22522),
            .I(N__22519));
    Span4Mux_v I__2979 (
            .O(N__22519),
            .I(N__22515));
    InMux I__2978 (
            .O(N__22518),
            .I(N__22512));
    Odrv4 I__2977 (
            .O(N__22515),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__2976 (
            .O(N__22512),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__2975 (
            .O(N__22507),
            .I(N__22504));
    LocalMux I__2974 (
            .O(N__22504),
            .I(N__22501));
    Span4Mux_h I__2973 (
            .O(N__22501),
            .I(N__22498));
    Odrv4 I__2972 (
            .O(N__22498),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ));
    InMux I__2971 (
            .O(N__22495),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__2970 (
            .O(N__22492),
            .I(N__22489));
    LocalMux I__2969 (
            .O(N__22489),
            .I(N__22486));
    Span4Mux_v I__2968 (
            .O(N__22486),
            .I(N__22482));
    InMux I__2967 (
            .O(N__22485),
            .I(N__22479));
    Odrv4 I__2966 (
            .O(N__22482),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__2965 (
            .O(N__22479),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__2964 (
            .O(N__22474),
            .I(N__22471));
    LocalMux I__2963 (
            .O(N__22471),
            .I(N__22468));
    Span4Mux_h I__2962 (
            .O(N__22468),
            .I(N__22465));
    Odrv4 I__2961 (
            .O(N__22465),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ));
    InMux I__2960 (
            .O(N__22462),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__2959 (
            .O(N__22459),
            .I(N__22456));
    LocalMux I__2958 (
            .O(N__22456),
            .I(N__22453));
    Span4Mux_h I__2957 (
            .O(N__22453),
            .I(N__22449));
    InMux I__2956 (
            .O(N__22452),
            .I(N__22446));
    Odrv4 I__2955 (
            .O(N__22449),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__2954 (
            .O(N__22446),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__2953 (
            .O(N__22441),
            .I(N__22438));
    LocalMux I__2952 (
            .O(N__22438),
            .I(N__22435));
    Span4Mux_v I__2951 (
            .O(N__22435),
            .I(N__22432));
    Odrv4 I__2950 (
            .O(N__22432),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ));
    InMux I__2949 (
            .O(N__22429),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__2948 (
            .O(N__22426),
            .I(N__22423));
    LocalMux I__2947 (
            .O(N__22423),
            .I(N__22420));
    Span4Mux_h I__2946 (
            .O(N__22420),
            .I(N__22416));
    InMux I__2945 (
            .O(N__22419),
            .I(N__22413));
    Odrv4 I__2944 (
            .O(N__22416),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__2943 (
            .O(N__22413),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__2942 (
            .O(N__22408),
            .I(N__22405));
    LocalMux I__2941 (
            .O(N__22405),
            .I(N__22402));
    Span4Mux_h I__2940 (
            .O(N__22402),
            .I(N__22399));
    Odrv4 I__2939 (
            .O(N__22399),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ));
    InMux I__2938 (
            .O(N__22396),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__2937 (
            .O(N__22393),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__2936 (
            .O(N__22390),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__2935 (
            .O(N__22387),
            .I(bfn_7_14_0_));
    InMux I__2934 (
            .O(N__22384),
            .I(N__22381));
    LocalMux I__2933 (
            .O(N__22381),
            .I(N__22378));
    Odrv12 I__2932 (
            .O(N__22378),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__2931 (
            .O(N__22375),
            .I(N__22372));
    LocalMux I__2930 (
            .O(N__22372),
            .I(N__22369));
    Span4Mux_h I__2929 (
            .O(N__22369),
            .I(N__22366));
    Odrv4 I__2928 (
            .O(N__22366),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    CascadeMux I__2927 (
            .O(N__22363),
            .I(N__22360));
    InMux I__2926 (
            .O(N__22360),
            .I(N__22357));
    LocalMux I__2925 (
            .O(N__22357),
            .I(N__22354));
    Span4Mux_h I__2924 (
            .O(N__22354),
            .I(N__22351));
    Odrv4 I__2923 (
            .O(N__22351),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__2922 (
            .O(N__22348),
            .I(N__22345));
    InMux I__2921 (
            .O(N__22345),
            .I(N__22342));
    LocalMux I__2920 (
            .O(N__22342),
            .I(N__22339));
    Span4Mux_v I__2919 (
            .O(N__22339),
            .I(N__22336));
    Span4Mux_h I__2918 (
            .O(N__22336),
            .I(N__22333));
    Odrv4 I__2917 (
            .O(N__22333),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__2916 (
            .O(N__22330),
            .I(N__22327));
    InMux I__2915 (
            .O(N__22327),
            .I(N__22324));
    LocalMux I__2914 (
            .O(N__22324),
            .I(N__22321));
    Span4Mux_h I__2913 (
            .O(N__22321),
            .I(N__22318));
    Odrv4 I__2912 (
            .O(N__22318),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__2911 (
            .O(N__22315),
            .I(N__22312));
    InMux I__2910 (
            .O(N__22312),
            .I(N__22309));
    LocalMux I__2909 (
            .O(N__22309),
            .I(N__22306));
    Span4Mux_h I__2908 (
            .O(N__22306),
            .I(N__22303));
    Odrv4 I__2907 (
            .O(N__22303),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__2906 (
            .O(N__22300),
            .I(N__22297));
    InMux I__2905 (
            .O(N__22297),
            .I(N__22293));
    InMux I__2904 (
            .O(N__22296),
            .I(N__22290));
    LocalMux I__2903 (
            .O(N__22293),
            .I(N__22287));
    LocalMux I__2902 (
            .O(N__22290),
            .I(N__22283));
    Span4Mux_v I__2901 (
            .O(N__22287),
            .I(N__22280));
    InMux I__2900 (
            .O(N__22286),
            .I(N__22277));
    Odrv4 I__2899 (
            .O(N__22283),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__2898 (
            .O(N__22280),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__2897 (
            .O(N__22277),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__2896 (
            .O(N__22270),
            .I(N__22267));
    InMux I__2895 (
            .O(N__22267),
            .I(N__22264));
    LocalMux I__2894 (
            .O(N__22264),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    CascadeMux I__2893 (
            .O(N__22261),
            .I(N__22258));
    InMux I__2892 (
            .O(N__22258),
            .I(N__22255));
    LocalMux I__2891 (
            .O(N__22255),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    CascadeMux I__2890 (
            .O(N__22252),
            .I(N__22249));
    InMux I__2889 (
            .O(N__22249),
            .I(N__22246));
    LocalMux I__2888 (
            .O(N__22246),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    CascadeMux I__2887 (
            .O(N__22243),
            .I(N__22240));
    InMux I__2886 (
            .O(N__22240),
            .I(N__22237));
    LocalMux I__2885 (
            .O(N__22237),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    CascadeMux I__2884 (
            .O(N__22234),
            .I(N__22231));
    InMux I__2883 (
            .O(N__22231),
            .I(N__22228));
    LocalMux I__2882 (
            .O(N__22228),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    CascadeMux I__2881 (
            .O(N__22225),
            .I(N__22222));
    InMux I__2880 (
            .O(N__22222),
            .I(N__22219));
    LocalMux I__2879 (
            .O(N__22219),
            .I(N__22216));
    Odrv4 I__2878 (
            .O(N__22216),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__2877 (
            .O(N__22213),
            .I(N__22210));
    InMux I__2876 (
            .O(N__22210),
            .I(N__22207));
    LocalMux I__2875 (
            .O(N__22207),
            .I(N__22204));
    Odrv4 I__2874 (
            .O(N__22204),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    CascadeMux I__2873 (
            .O(N__22201),
            .I(N__22194));
    CascadeMux I__2872 (
            .O(N__22200),
            .I(N__22190));
    CascadeMux I__2871 (
            .O(N__22199),
            .I(N__22186));
    InMux I__2870 (
            .O(N__22198),
            .I(N__22171));
    InMux I__2869 (
            .O(N__22197),
            .I(N__22171));
    InMux I__2868 (
            .O(N__22194),
            .I(N__22171));
    InMux I__2867 (
            .O(N__22193),
            .I(N__22171));
    InMux I__2866 (
            .O(N__22190),
            .I(N__22171));
    InMux I__2865 (
            .O(N__22189),
            .I(N__22171));
    InMux I__2864 (
            .O(N__22186),
            .I(N__22171));
    LocalMux I__2863 (
            .O(N__22171),
            .I(N__22168));
    Odrv4 I__2862 (
            .O(N__22168),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    CascadeMux I__2861 (
            .O(N__22165),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ));
    InMux I__2860 (
            .O(N__22162),
            .I(N__22159));
    LocalMux I__2859 (
            .O(N__22159),
            .I(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ));
    CascadeMux I__2858 (
            .O(N__22156),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    CascadeMux I__2857 (
            .O(N__22153),
            .I(N__22150));
    InMux I__2856 (
            .O(N__22150),
            .I(N__22147));
    LocalMux I__2855 (
            .O(N__22147),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__2854 (
            .O(N__22144),
            .I(N__22141));
    LocalMux I__2853 (
            .O(N__22141),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__2852 (
            .O(N__22138),
            .I(N__22135));
    InMux I__2851 (
            .O(N__22135),
            .I(N__22132));
    LocalMux I__2850 (
            .O(N__22132),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__2849 (
            .O(N__22129),
            .I(N__22126));
    LocalMux I__2848 (
            .O(N__22126),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__2847 (
            .O(N__22123),
            .I(N__22120));
    InMux I__2846 (
            .O(N__22120),
            .I(N__22117));
    LocalMux I__2845 (
            .O(N__22117),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__2844 (
            .O(N__22114),
            .I(N__22111));
    InMux I__2843 (
            .O(N__22111),
            .I(N__22108));
    LocalMux I__2842 (
            .O(N__22108),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__2841 (
            .O(N__22105),
            .I(N__22102));
    LocalMux I__2840 (
            .O(N__22102),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    InMux I__2839 (
            .O(N__22099),
            .I(N__22096));
    LocalMux I__2838 (
            .O(N__22096),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__2837 (
            .O(N__22093),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__2836 (
            .O(N__22090),
            .I(N__22087));
    LocalMux I__2835 (
            .O(N__22087),
            .I(N__22084));
    Odrv12 I__2834 (
            .O(N__22084),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__2833 (
            .O(N__22081),
            .I(N__22078));
    InMux I__2832 (
            .O(N__22078),
            .I(N__22075));
    LocalMux I__2831 (
            .O(N__22075),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__2830 (
            .O(N__22072),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ));
    InMux I__2829 (
            .O(N__22069),
            .I(N__22066));
    LocalMux I__2828 (
            .O(N__22066),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__2827 (
            .O(N__22063),
            .I(N__22060));
    LocalMux I__2826 (
            .O(N__22060),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__2825 (
            .O(N__22057),
            .I(N__22054));
    LocalMux I__2824 (
            .O(N__22054),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__2823 (
            .O(N__22051),
            .I(N__22048));
    LocalMux I__2822 (
            .O(N__22048),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__2821 (
            .O(N__22045),
            .I(N__22042));
    LocalMux I__2820 (
            .O(N__22042),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__2819 (
            .O(N__22039),
            .I(N__22036));
    LocalMux I__2818 (
            .O(N__22036),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__2817 (
            .O(N__22033),
            .I(N__22030));
    InMux I__2816 (
            .O(N__22030),
            .I(N__22027));
    LocalMux I__2815 (
            .O(N__22027),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__2814 (
            .O(N__22024),
            .I(N__22021));
    LocalMux I__2813 (
            .O(N__22021),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    InMux I__2812 (
            .O(N__22018),
            .I(N__22015));
    LocalMux I__2811 (
            .O(N__22015),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    CascadeMux I__2810 (
            .O(N__22012),
            .I(N__22009));
    InMux I__2809 (
            .O(N__22009),
            .I(N__22006));
    LocalMux I__2808 (
            .O(N__22006),
            .I(N__22003));
    Odrv4 I__2807 (
            .O(N__22003),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__2806 (
            .O(N__22000),
            .I(N__21997));
    LocalMux I__2805 (
            .O(N__21997),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__2804 (
            .O(N__21994),
            .I(N__21991));
    InMux I__2803 (
            .O(N__21991),
            .I(N__21988));
    LocalMux I__2802 (
            .O(N__21988),
            .I(N__21985));
    Odrv4 I__2801 (
            .O(N__21985),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    InMux I__2800 (
            .O(N__21982),
            .I(N__21979));
    LocalMux I__2799 (
            .O(N__21979),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__2798 (
            .O(N__21976),
            .I(N__21973));
    InMux I__2797 (
            .O(N__21973),
            .I(N__21970));
    LocalMux I__2796 (
            .O(N__21970),
            .I(N__21967));
    Odrv12 I__2795 (
            .O(N__21967),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__2794 (
            .O(N__21964),
            .I(N__21961));
    LocalMux I__2793 (
            .O(N__21961),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__2792 (
            .O(N__21958),
            .I(N__21955));
    InMux I__2791 (
            .O(N__21955),
            .I(N__21952));
    LocalMux I__2790 (
            .O(N__21952),
            .I(N__21949));
    Odrv12 I__2789 (
            .O(N__21949),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__2788 (
            .O(N__21946),
            .I(N__21943));
    LocalMux I__2787 (
            .O(N__21943),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__2786 (
            .O(N__21940),
            .I(N__21937));
    InMux I__2785 (
            .O(N__21937),
            .I(N__21934));
    LocalMux I__2784 (
            .O(N__21934),
            .I(N__21931));
    Span4Mux_h I__2783 (
            .O(N__21931),
            .I(N__21928));
    Odrv4 I__2782 (
            .O(N__21928),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__2781 (
            .O(N__21925),
            .I(N__21922));
    LocalMux I__2780 (
            .O(N__21922),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__2779 (
            .O(N__21919),
            .I(N__21916));
    LocalMux I__2778 (
            .O(N__21916),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__2777 (
            .O(N__21913),
            .I(N__21910));
    LocalMux I__2776 (
            .O(N__21910),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__2775 (
            .O(N__21907),
            .I(N__21904));
    InMux I__2774 (
            .O(N__21904),
            .I(N__21901));
    LocalMux I__2773 (
            .O(N__21901),
            .I(N__21898));
    Span4Mux_h I__2772 (
            .O(N__21898),
            .I(N__21895));
    Odrv4 I__2771 (
            .O(N__21895),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    InMux I__2770 (
            .O(N__21892),
            .I(N__21889));
    LocalMux I__2769 (
            .O(N__21889),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__2768 (
            .O(N__21886),
            .I(N__21883));
    LocalMux I__2767 (
            .O(N__21883),
            .I(N__21880));
    Odrv4 I__2766 (
            .O(N__21880),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ));
    CascadeMux I__2765 (
            .O(N__21877),
            .I(un2_counter_5_cascade_));
    CascadeMux I__2764 (
            .O(N__21874),
            .I(N__21869));
    InMux I__2763 (
            .O(N__21873),
            .I(N__21866));
    InMux I__2762 (
            .O(N__21872),
            .I(N__21860));
    InMux I__2761 (
            .O(N__21869),
            .I(N__21860));
    LocalMux I__2760 (
            .O(N__21866),
            .I(N__21857));
    InMux I__2759 (
            .O(N__21865),
            .I(N__21854));
    LocalMux I__2758 (
            .O(N__21860),
            .I(counterZ0Z_0));
    Odrv4 I__2757 (
            .O(N__21857),
            .I(counterZ0Z_0));
    LocalMux I__2756 (
            .O(N__21854),
            .I(counterZ0Z_0));
    InMux I__2755 (
            .O(N__21847),
            .I(N__21843));
    InMux I__2754 (
            .O(N__21846),
            .I(N__21840));
    LocalMux I__2753 (
            .O(N__21843),
            .I(counterZ0Z_11));
    LocalMux I__2752 (
            .O(N__21840),
            .I(counterZ0Z_11));
    InMux I__2751 (
            .O(N__21835),
            .I(N__21831));
    InMux I__2750 (
            .O(N__21834),
            .I(N__21828));
    LocalMux I__2749 (
            .O(N__21831),
            .I(counterZ0Z_9));
    LocalMux I__2748 (
            .O(N__21828),
            .I(counterZ0Z_9));
    CascadeMux I__2747 (
            .O(N__21823),
            .I(N__21819));
    InMux I__2746 (
            .O(N__21822),
            .I(N__21816));
    InMux I__2745 (
            .O(N__21819),
            .I(N__21813));
    LocalMux I__2744 (
            .O(N__21816),
            .I(counterZ0Z_12));
    LocalMux I__2743 (
            .O(N__21813),
            .I(counterZ0Z_12));
    InMux I__2742 (
            .O(N__21808),
            .I(N__21804));
    InMux I__2741 (
            .O(N__21807),
            .I(N__21801));
    LocalMux I__2740 (
            .O(N__21804),
            .I(N__21798));
    LocalMux I__2739 (
            .O(N__21801),
            .I(counterZ0Z_8));
    Odrv4 I__2738 (
            .O(N__21798),
            .I(counterZ0Z_8));
    InMux I__2737 (
            .O(N__21793),
            .I(N__21787));
    InMux I__2736 (
            .O(N__21792),
            .I(N__21782));
    InMux I__2735 (
            .O(N__21791),
            .I(N__21779));
    InMux I__2734 (
            .O(N__21790),
            .I(N__21776));
    LocalMux I__2733 (
            .O(N__21787),
            .I(N__21773));
    InMux I__2732 (
            .O(N__21786),
            .I(N__21770));
    InMux I__2731 (
            .O(N__21785),
            .I(N__21767));
    LocalMux I__2730 (
            .O(N__21782),
            .I(N__21760));
    LocalMux I__2729 (
            .O(N__21779),
            .I(N__21760));
    LocalMux I__2728 (
            .O(N__21776),
            .I(N__21760));
    Odrv4 I__2727 (
            .O(N__21773),
            .I(un2_counter_7));
    LocalMux I__2726 (
            .O(N__21770),
            .I(un2_counter_7));
    LocalMux I__2725 (
            .O(N__21767),
            .I(un2_counter_7));
    Odrv4 I__2724 (
            .O(N__21760),
            .I(un2_counter_7));
    InMux I__2723 (
            .O(N__21751),
            .I(N__21741));
    InMux I__2722 (
            .O(N__21750),
            .I(N__21741));
    InMux I__2721 (
            .O(N__21749),
            .I(N__21736));
    InMux I__2720 (
            .O(N__21748),
            .I(N__21736));
    InMux I__2719 (
            .O(N__21747),
            .I(N__21733));
    InMux I__2718 (
            .O(N__21746),
            .I(N__21730));
    LocalMux I__2717 (
            .O(N__21741),
            .I(un2_counter_8));
    LocalMux I__2716 (
            .O(N__21736),
            .I(un2_counter_8));
    LocalMux I__2715 (
            .O(N__21733),
            .I(un2_counter_8));
    LocalMux I__2714 (
            .O(N__21730),
            .I(un2_counter_8));
    InMux I__2713 (
            .O(N__21721),
            .I(N__21711));
    InMux I__2712 (
            .O(N__21720),
            .I(N__21711));
    InMux I__2711 (
            .O(N__21719),
            .I(N__21706));
    InMux I__2710 (
            .O(N__21718),
            .I(N__21706));
    InMux I__2709 (
            .O(N__21717),
            .I(N__21703));
    InMux I__2708 (
            .O(N__21716),
            .I(N__21700));
    LocalMux I__2707 (
            .O(N__21711),
            .I(un2_counter_9));
    LocalMux I__2706 (
            .O(N__21706),
            .I(un2_counter_9));
    LocalMux I__2705 (
            .O(N__21703),
            .I(un2_counter_9));
    LocalMux I__2704 (
            .O(N__21700),
            .I(un2_counter_9));
    CascadeMux I__2703 (
            .O(N__21691),
            .I(N__21686));
    InMux I__2702 (
            .O(N__21690),
            .I(N__21683));
    CascadeMux I__2701 (
            .O(N__21689),
            .I(N__21679));
    InMux I__2700 (
            .O(N__21686),
            .I(N__21676));
    LocalMux I__2699 (
            .O(N__21683),
            .I(N__21673));
    InMux I__2698 (
            .O(N__21682),
            .I(N__21670));
    InMux I__2697 (
            .O(N__21679),
            .I(N__21667));
    LocalMux I__2696 (
            .O(N__21676),
            .I(clk_10khz_i));
    Odrv4 I__2695 (
            .O(N__21673),
            .I(clk_10khz_i));
    LocalMux I__2694 (
            .O(N__21670),
            .I(clk_10khz_i));
    LocalMux I__2693 (
            .O(N__21667),
            .I(clk_10khz_i));
    CascadeMux I__2692 (
            .O(N__21658),
            .I(N__21654));
    InMux I__2691 (
            .O(N__21657),
            .I(N__21651));
    InMux I__2690 (
            .O(N__21654),
            .I(N__21648));
    LocalMux I__2689 (
            .O(N__21651),
            .I(counterZ0Z_6));
    LocalMux I__2688 (
            .O(N__21648),
            .I(counterZ0Z_6));
    InMux I__2687 (
            .O(N__21643),
            .I(un5_counter_cry_5));
    CascadeMux I__2686 (
            .O(N__21640),
            .I(N__21637));
    InMux I__2685 (
            .O(N__21637),
            .I(N__21634));
    LocalMux I__2684 (
            .O(N__21634),
            .I(counter_RNO_0Z0Z_7));
    InMux I__2683 (
            .O(N__21631),
            .I(un5_counter_cry_6));
    InMux I__2682 (
            .O(N__21628),
            .I(un5_counter_cry_7));
    InMux I__2681 (
            .O(N__21625),
            .I(bfn_5_8_0_));
    CascadeMux I__2680 (
            .O(N__21622),
            .I(N__21619));
    InMux I__2679 (
            .O(N__21619),
            .I(N__21616));
    LocalMux I__2678 (
            .O(N__21616),
            .I(counter_RNO_0Z0Z_10));
    InMux I__2677 (
            .O(N__21613),
            .I(un5_counter_cry_9));
    InMux I__2676 (
            .O(N__21610),
            .I(un5_counter_cry_10));
    InMux I__2675 (
            .O(N__21607),
            .I(un5_counter_cry_11));
    CascadeMux I__2674 (
            .O(N__21604),
            .I(N__21601));
    InMux I__2673 (
            .O(N__21601),
            .I(N__21598));
    LocalMux I__2672 (
            .O(N__21598),
            .I(counter_RNO_0Z0Z_12));
    InMux I__2671 (
            .O(N__21595),
            .I(N__21591));
    InMux I__2670 (
            .O(N__21594),
            .I(N__21588));
    LocalMux I__2669 (
            .O(N__21591),
            .I(counterZ0Z_10));
    LocalMux I__2668 (
            .O(N__21588),
            .I(counterZ0Z_10));
    InMux I__2667 (
            .O(N__21583),
            .I(N__21579));
    InMux I__2666 (
            .O(N__21582),
            .I(N__21576));
    LocalMux I__2665 (
            .O(N__21579),
            .I(counterZ0Z_7));
    LocalMux I__2664 (
            .O(N__21576),
            .I(counterZ0Z_7));
    InMux I__2663 (
            .O(N__21571),
            .I(N__21567));
    InMux I__2662 (
            .O(N__21570),
            .I(N__21564));
    LocalMux I__2661 (
            .O(N__21567),
            .I(N__21561));
    LocalMux I__2660 (
            .O(N__21564),
            .I(counterZ0Z_2));
    Odrv12 I__2659 (
            .O(N__21561),
            .I(counterZ0Z_2));
    CascadeMux I__2658 (
            .O(N__21556),
            .I(N__21553));
    InMux I__2657 (
            .O(N__21553),
            .I(N__21549));
    InMux I__2656 (
            .O(N__21552),
            .I(N__21545));
    LocalMux I__2655 (
            .O(N__21549),
            .I(N__21542));
    InMux I__2654 (
            .O(N__21548),
            .I(N__21539));
    LocalMux I__2653 (
            .O(N__21545),
            .I(counterZ0Z_1));
    Odrv4 I__2652 (
            .O(N__21542),
            .I(counterZ0Z_1));
    LocalMux I__2651 (
            .O(N__21539),
            .I(counterZ0Z_1));
    InMux I__2650 (
            .O(N__21532),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    CascadeMux I__2649 (
            .O(N__21529),
            .I(N__21523));
    InMux I__2648 (
            .O(N__21528),
            .I(N__21518));
    CascadeMux I__2647 (
            .O(N__21527),
            .I(N__21515));
    CascadeMux I__2646 (
            .O(N__21526),
            .I(N__21509));
    InMux I__2645 (
            .O(N__21523),
            .I(N__21506));
    InMux I__2644 (
            .O(N__21522),
            .I(N__21500));
    InMux I__2643 (
            .O(N__21521),
            .I(N__21500));
    LocalMux I__2642 (
            .O(N__21518),
            .I(N__21497));
    InMux I__2641 (
            .O(N__21515),
            .I(N__21494));
    InMux I__2640 (
            .O(N__21514),
            .I(N__21485));
    InMux I__2639 (
            .O(N__21513),
            .I(N__21485));
    InMux I__2638 (
            .O(N__21512),
            .I(N__21485));
    InMux I__2637 (
            .O(N__21509),
            .I(N__21485));
    LocalMux I__2636 (
            .O(N__21506),
            .I(N__21482));
    InMux I__2635 (
            .O(N__21505),
            .I(N__21479));
    LocalMux I__2634 (
            .O(N__21500),
            .I(N__21476));
    Span12Mux_s7_v I__2633 (
            .O(N__21497),
            .I(N__21469));
    LocalMux I__2632 (
            .O(N__21494),
            .I(N__21469));
    LocalMux I__2631 (
            .O(N__21485),
            .I(N__21469));
    Span4Mux_h I__2630 (
            .O(N__21482),
            .I(N__21466));
    LocalMux I__2629 (
            .O(N__21479),
            .I(N__21463));
    Span4Mux_h I__2628 (
            .O(N__21476),
            .I(N__21460));
    Span12Mux_v I__2627 (
            .O(N__21469),
            .I(N__21457));
    Span4Mux_v I__2626 (
            .O(N__21466),
            .I(N__21454));
    Span12Mux_s4_h I__2625 (
            .O(N__21463),
            .I(N__21451));
    Span4Mux_v I__2624 (
            .O(N__21460),
            .I(N__21448));
    Odrv12 I__2623 (
            .O(N__21457),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2622 (
            .O(N__21454),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv12 I__2621 (
            .O(N__21451),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2620 (
            .O(N__21448),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    CascadeMux I__2619 (
            .O(N__21439),
            .I(N__21436));
    InMux I__2618 (
            .O(N__21436),
            .I(N__21433));
    LocalMux I__2617 (
            .O(N__21433),
            .I(N__21430));
    Odrv4 I__2616 (
            .O(N__21430),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__2615 (
            .O(N__21427),
            .I(N__21424));
    InMux I__2614 (
            .O(N__21424),
            .I(N__21421));
    LocalMux I__2613 (
            .O(N__21421),
            .I(N__21418));
    Odrv4 I__2612 (
            .O(N__21418),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    InMux I__2611 (
            .O(N__21415),
            .I(N__21412));
    LocalMux I__2610 (
            .O(N__21412),
            .I(N__21409));
    Span4Mux_s2_v I__2609 (
            .O(N__21409),
            .I(N__21406));
    Odrv4 I__2608 (
            .O(N__21406),
            .I(un7_start_stop_0_a3));
    InMux I__2607 (
            .O(N__21403),
            .I(un5_counter_cry_1));
    InMux I__2606 (
            .O(N__21400),
            .I(N__21396));
    InMux I__2605 (
            .O(N__21399),
            .I(N__21393));
    LocalMux I__2604 (
            .O(N__21396),
            .I(counterZ0Z_3));
    LocalMux I__2603 (
            .O(N__21393),
            .I(counterZ0Z_3));
    InMux I__2602 (
            .O(N__21388),
            .I(un5_counter_cry_2));
    InMux I__2601 (
            .O(N__21385),
            .I(N__21381));
    InMux I__2600 (
            .O(N__21384),
            .I(N__21378));
    LocalMux I__2599 (
            .O(N__21381),
            .I(counterZ0Z_4));
    LocalMux I__2598 (
            .O(N__21378),
            .I(counterZ0Z_4));
    InMux I__2597 (
            .O(N__21373),
            .I(un5_counter_cry_3));
    InMux I__2596 (
            .O(N__21370),
            .I(N__21366));
    InMux I__2595 (
            .O(N__21369),
            .I(N__21363));
    LocalMux I__2594 (
            .O(N__21366),
            .I(counterZ0Z_5));
    LocalMux I__2593 (
            .O(N__21363),
            .I(counterZ0Z_5));
    InMux I__2592 (
            .O(N__21358),
            .I(un5_counter_cry_4));
    InMux I__2591 (
            .O(N__21355),
            .I(N__21351));
    InMux I__2590 (
            .O(N__21354),
            .I(N__21348));
    LocalMux I__2589 (
            .O(N__21351),
            .I(N__21345));
    LocalMux I__2588 (
            .O(N__21348),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    Odrv4 I__2587 (
            .O(N__21345),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2586 (
            .O(N__21340),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__2585 (
            .O(N__21337),
            .I(N__21333));
    InMux I__2584 (
            .O(N__21336),
            .I(N__21330));
    LocalMux I__2583 (
            .O(N__21333),
            .I(N__21325));
    LocalMux I__2582 (
            .O(N__21330),
            .I(N__21325));
    Span4Mux_h I__2581 (
            .O(N__21325),
            .I(N__21322));
    Odrv4 I__2580 (
            .O(N__21322),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2579 (
            .O(N__21319),
            .I(bfn_4_20_0_));
    InMux I__2578 (
            .O(N__21316),
            .I(N__21312));
    InMux I__2577 (
            .O(N__21315),
            .I(N__21309));
    LocalMux I__2576 (
            .O(N__21312),
            .I(N__21306));
    LocalMux I__2575 (
            .O(N__21309),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    Odrv4 I__2574 (
            .O(N__21306),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2573 (
            .O(N__21301),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    InMux I__2572 (
            .O(N__21298),
            .I(N__21292));
    InMux I__2571 (
            .O(N__21297),
            .I(N__21292));
    LocalMux I__2570 (
            .O(N__21292),
            .I(N__21289));
    Odrv4 I__2569 (
            .O(N__21289),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2568 (
            .O(N__21286),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2567 (
            .O(N__21283),
            .I(N__21280));
    LocalMux I__2566 (
            .O(N__21280),
            .I(N__21276));
    InMux I__2565 (
            .O(N__21279),
            .I(N__21273));
    Odrv4 I__2564 (
            .O(N__21276),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    LocalMux I__2563 (
            .O(N__21273),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2562 (
            .O(N__21268),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2561 (
            .O(N__21265),
            .I(N__21262));
    LocalMux I__2560 (
            .O(N__21262),
            .I(N__21258));
    InMux I__2559 (
            .O(N__21261),
            .I(N__21255));
    Odrv4 I__2558 (
            .O(N__21258),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    LocalMux I__2557 (
            .O(N__21255),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2556 (
            .O(N__21250),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2555 (
            .O(N__21247),
            .I(N__21243));
    InMux I__2554 (
            .O(N__21246),
            .I(N__21240));
    LocalMux I__2553 (
            .O(N__21243),
            .I(N__21235));
    LocalMux I__2552 (
            .O(N__21240),
            .I(N__21235));
    Odrv4 I__2551 (
            .O(N__21235),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2550 (
            .O(N__21232),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    CascadeMux I__2549 (
            .O(N__21229),
            .I(N__21226));
    InMux I__2548 (
            .O(N__21226),
            .I(N__21222));
    InMux I__2547 (
            .O(N__21225),
            .I(N__21219));
    LocalMux I__2546 (
            .O(N__21222),
            .I(N__21216));
    LocalMux I__2545 (
            .O(N__21219),
            .I(N__21211));
    Span4Mux_h I__2544 (
            .O(N__21216),
            .I(N__21211));
    Odrv4 I__2543 (
            .O(N__21211),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2542 (
            .O(N__21208),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2541 (
            .O(N__21205),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    CascadeMux I__2540 (
            .O(N__21202),
            .I(N__21199));
    InMux I__2539 (
            .O(N__21199),
            .I(N__21196));
    LocalMux I__2538 (
            .O(N__21196),
            .I(N__21193));
    Span4Mux_h I__2537 (
            .O(N__21193),
            .I(N__21190));
    Odrv4 I__2536 (
            .O(N__21190),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    CascadeMux I__2535 (
            .O(N__21187),
            .I(N__21184));
    InMux I__2534 (
            .O(N__21184),
            .I(N__21180));
    InMux I__2533 (
            .O(N__21183),
            .I(N__21177));
    LocalMux I__2532 (
            .O(N__21180),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__2531 (
            .O(N__21177),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2530 (
            .O(N__21172),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__2529 (
            .O(N__21169),
            .I(N__21166));
    LocalMux I__2528 (
            .O(N__21166),
            .I(N__21163));
    Span4Mux_v I__2527 (
            .O(N__21163),
            .I(N__21159));
    InMux I__2526 (
            .O(N__21162),
            .I(N__21156));
    Odrv4 I__2525 (
            .O(N__21159),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    LocalMux I__2524 (
            .O(N__21156),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2523 (
            .O(N__21151),
            .I(bfn_4_19_0_));
    CascadeMux I__2522 (
            .O(N__21148),
            .I(N__21145));
    InMux I__2521 (
            .O(N__21145),
            .I(N__21142));
    LocalMux I__2520 (
            .O(N__21142),
            .I(N__21139));
    Odrv4 I__2519 (
            .O(N__21139),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    CascadeMux I__2518 (
            .O(N__21136),
            .I(N__21133));
    InMux I__2517 (
            .O(N__21133),
            .I(N__21130));
    LocalMux I__2516 (
            .O(N__21130),
            .I(N__21126));
    InMux I__2515 (
            .O(N__21129),
            .I(N__21123));
    Odrv4 I__2514 (
            .O(N__21126),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    LocalMux I__2513 (
            .O(N__21123),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2512 (
            .O(N__21118),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    InMux I__2511 (
            .O(N__21115),
            .I(N__21111));
    CascadeMux I__2510 (
            .O(N__21114),
            .I(N__21108));
    LocalMux I__2509 (
            .O(N__21111),
            .I(N__21105));
    InMux I__2508 (
            .O(N__21108),
            .I(N__21102));
    Odrv4 I__2507 (
            .O(N__21105),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    LocalMux I__2506 (
            .O(N__21102),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2505 (
            .O(N__21097),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2504 (
            .O(N__21094),
            .I(N__21088));
    InMux I__2503 (
            .O(N__21093),
            .I(N__21088));
    LocalMux I__2502 (
            .O(N__21088),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2501 (
            .O(N__21085),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    CascadeMux I__2500 (
            .O(N__21082),
            .I(N__21079));
    InMux I__2499 (
            .O(N__21079),
            .I(N__21073));
    InMux I__2498 (
            .O(N__21078),
            .I(N__21073));
    LocalMux I__2497 (
            .O(N__21073),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2496 (
            .O(N__21070),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__2495 (
            .O(N__21067),
            .I(N__21063));
    InMux I__2494 (
            .O(N__21066),
            .I(N__21060));
    LocalMux I__2493 (
            .O(N__21063),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    LocalMux I__2492 (
            .O(N__21060),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2491 (
            .O(N__21055),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    CascadeMux I__2490 (
            .O(N__21052),
            .I(N__21048));
    InMux I__2489 (
            .O(N__21051),
            .I(N__21043));
    InMux I__2488 (
            .O(N__21048),
            .I(N__21043));
    LocalMux I__2487 (
            .O(N__21043),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2486 (
            .O(N__21040),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    CascadeMux I__2485 (
            .O(N__21037),
            .I(N__21034));
    InMux I__2484 (
            .O(N__21034),
            .I(N__21030));
    InMux I__2483 (
            .O(N__21033),
            .I(N__21026));
    LocalMux I__2482 (
            .O(N__21030),
            .I(N__21023));
    InMux I__2481 (
            .O(N__21029),
            .I(N__21020));
    LocalMux I__2480 (
            .O(N__21026),
            .I(N__21017));
    Span4Mux_h I__2479 (
            .O(N__21023),
            .I(N__21012));
    LocalMux I__2478 (
            .O(N__21020),
            .I(N__21012));
    Span4Mux_h I__2477 (
            .O(N__21017),
            .I(N__21009));
    Span4Mux_v I__2476 (
            .O(N__21012),
            .I(N__21006));
    Odrv4 I__2475 (
            .O(N__21009),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2474 (
            .O(N__21006),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2473 (
            .O(N__21001),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    CascadeMux I__2472 (
            .O(N__20998),
            .I(N__20995));
    InMux I__2471 (
            .O(N__20995),
            .I(N__20991));
    InMux I__2470 (
            .O(N__20994),
            .I(N__20987));
    LocalMux I__2469 (
            .O(N__20991),
            .I(N__20984));
    InMux I__2468 (
            .O(N__20990),
            .I(N__20981));
    LocalMux I__2467 (
            .O(N__20987),
            .I(N__20978));
    Span4Mux_h I__2466 (
            .O(N__20984),
            .I(N__20973));
    LocalMux I__2465 (
            .O(N__20981),
            .I(N__20973));
    Span4Mux_h I__2464 (
            .O(N__20978),
            .I(N__20970));
    Span4Mux_v I__2463 (
            .O(N__20973),
            .I(N__20967));
    Odrv4 I__2462 (
            .O(N__20970),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__2461 (
            .O(N__20967),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2460 (
            .O(N__20962),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    CascadeMux I__2459 (
            .O(N__20959),
            .I(N__20956));
    InMux I__2458 (
            .O(N__20956),
            .I(N__20953));
    LocalMux I__2457 (
            .O(N__20953),
            .I(N__20949));
    InMux I__2456 (
            .O(N__20952),
            .I(N__20946));
    Span4Mux_h I__2455 (
            .O(N__20949),
            .I(N__20942));
    LocalMux I__2454 (
            .O(N__20946),
            .I(N__20939));
    InMux I__2453 (
            .O(N__20945),
            .I(N__20936));
    Span4Mux_v I__2452 (
            .O(N__20942),
            .I(N__20933));
    Span4Mux_h I__2451 (
            .O(N__20939),
            .I(N__20930));
    LocalMux I__2450 (
            .O(N__20936),
            .I(N__20927));
    Odrv4 I__2449 (
            .O(N__20933),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2448 (
            .O(N__20930),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv12 I__2447 (
            .O(N__20927),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2446 (
            .O(N__20920),
            .I(bfn_4_18_0_));
    InMux I__2445 (
            .O(N__20917),
            .I(N__20914));
    LocalMux I__2444 (
            .O(N__20914),
            .I(N__20911));
    Span4Mux_v I__2443 (
            .O(N__20911),
            .I(N__20907));
    InMux I__2442 (
            .O(N__20910),
            .I(N__20904));
    Span4Mux_v I__2441 (
            .O(N__20907),
            .I(N__20900));
    LocalMux I__2440 (
            .O(N__20904),
            .I(N__20897));
    InMux I__2439 (
            .O(N__20903),
            .I(N__20894));
    Span4Mux_h I__2438 (
            .O(N__20900),
            .I(N__20891));
    Span4Mux_h I__2437 (
            .O(N__20897),
            .I(N__20888));
    LocalMux I__2436 (
            .O(N__20894),
            .I(N__20885));
    Odrv4 I__2435 (
            .O(N__20891),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv4 I__2434 (
            .O(N__20888),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv12 I__2433 (
            .O(N__20885),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2432 (
            .O(N__20878),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    CascadeMux I__2431 (
            .O(N__20875),
            .I(N__20871));
    InMux I__2430 (
            .O(N__20874),
            .I(N__20868));
    InMux I__2429 (
            .O(N__20871),
            .I(N__20865));
    LocalMux I__2428 (
            .O(N__20868),
            .I(N__20860));
    LocalMux I__2427 (
            .O(N__20865),
            .I(N__20860));
    Odrv4 I__2426 (
            .O(N__20860),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2425 (
            .O(N__20857),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2424 (
            .O(N__20854),
            .I(N__20851));
    LocalMux I__2423 (
            .O(N__20851),
            .I(N__20847));
    InMux I__2422 (
            .O(N__20850),
            .I(N__20844));
    Odrv4 I__2421 (
            .O(N__20847),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    LocalMux I__2420 (
            .O(N__20844),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2419 (
            .O(N__20839),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2418 (
            .O(N__20836),
            .I(N__20830));
    InMux I__2417 (
            .O(N__20835),
            .I(N__20830));
    LocalMux I__2416 (
            .O(N__20830),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2415 (
            .O(N__20827),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2414 (
            .O(N__20824),
            .I(N__20821));
    LocalMux I__2413 (
            .O(N__20821),
            .I(N__20817));
    InMux I__2412 (
            .O(N__20820),
            .I(N__20814));
    Odrv4 I__2411 (
            .O(N__20817),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    LocalMux I__2410 (
            .O(N__20814),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2409 (
            .O(N__20809),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__2408 (
            .O(N__20806),
            .I(N__20800));
    InMux I__2407 (
            .O(N__20805),
            .I(N__20800));
    LocalMux I__2406 (
            .O(N__20800),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    CascadeMux I__2405 (
            .O(N__20797),
            .I(N__20794));
    InMux I__2404 (
            .O(N__20794),
            .I(N__20791));
    LocalMux I__2403 (
            .O(N__20791),
            .I(N__20788));
    Span4Mux_h I__2402 (
            .O(N__20788),
            .I(N__20785));
    Odrv4 I__2401 (
            .O(N__20785),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    CascadeMux I__2400 (
            .O(N__20782),
            .I(N__20779));
    InMux I__2399 (
            .O(N__20779),
            .I(N__20776));
    LocalMux I__2398 (
            .O(N__20776),
            .I(N__20773));
    Span4Mux_h I__2397 (
            .O(N__20773),
            .I(N__20770));
    Span4Mux_v I__2396 (
            .O(N__20770),
            .I(N__20767));
    Odrv4 I__2395 (
            .O(N__20767),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    CascadeMux I__2394 (
            .O(N__20764),
            .I(N__20761));
    InMux I__2393 (
            .O(N__20761),
            .I(N__20758));
    LocalMux I__2392 (
            .O(N__20758),
            .I(N__20755));
    Span4Mux_h I__2391 (
            .O(N__20755),
            .I(N__20752));
    Span4Mux_v I__2390 (
            .O(N__20752),
            .I(N__20749));
    Odrv4 I__2389 (
            .O(N__20749),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2388 (
            .O(N__20746),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    CascadeMux I__2387 (
            .O(N__20743),
            .I(N__20740));
    InMux I__2386 (
            .O(N__20740),
            .I(N__20737));
    LocalMux I__2385 (
            .O(N__20737),
            .I(N__20734));
    Span4Mux_h I__2384 (
            .O(N__20734),
            .I(N__20731));
    Odrv4 I__2383 (
            .O(N__20731),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__2382 (
            .O(N__20728),
            .I(N__20725));
    InMux I__2381 (
            .O(N__20725),
            .I(N__20722));
    LocalMux I__2380 (
            .O(N__20722),
            .I(N__20719));
    Span4Mux_v I__2379 (
            .O(N__20719),
            .I(N__20716));
    Span4Mux_h I__2378 (
            .O(N__20716),
            .I(N__20713));
    Odrv4 I__2377 (
            .O(N__20713),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2376 (
            .O(N__20710),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2375 (
            .O(N__20707),
            .I(N__20703));
    CascadeMux I__2374 (
            .O(N__20706),
            .I(N__20700));
    LocalMux I__2373 (
            .O(N__20703),
            .I(N__20696));
    InMux I__2372 (
            .O(N__20700),
            .I(N__20693));
    InMux I__2371 (
            .O(N__20699),
            .I(N__20690));
    Span4Mux_h I__2370 (
            .O(N__20696),
            .I(N__20687));
    LocalMux I__2369 (
            .O(N__20693),
            .I(N__20682));
    LocalMux I__2368 (
            .O(N__20690),
            .I(N__20682));
    Span4Mux_v I__2367 (
            .O(N__20687),
            .I(N__20677));
    Span4Mux_h I__2366 (
            .O(N__20682),
            .I(N__20677));
    Odrv4 I__2365 (
            .O(N__20677),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2364 (
            .O(N__20674),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    CascadeMux I__2363 (
            .O(N__20671),
            .I(N__20668));
    InMux I__2362 (
            .O(N__20668),
            .I(N__20664));
    InMux I__2361 (
            .O(N__20667),
            .I(N__20661));
    LocalMux I__2360 (
            .O(N__20664),
            .I(N__20656));
    LocalMux I__2359 (
            .O(N__20661),
            .I(N__20653));
    InMux I__2358 (
            .O(N__20660),
            .I(N__20650));
    InMux I__2357 (
            .O(N__20659),
            .I(N__20647));
    Span4Mux_v I__2356 (
            .O(N__20656),
            .I(N__20638));
    Span4Mux_s2_h I__2355 (
            .O(N__20653),
            .I(N__20638));
    LocalMux I__2354 (
            .O(N__20650),
            .I(N__20638));
    LocalMux I__2353 (
            .O(N__20647),
            .I(N__20638));
    Span4Mux_v I__2352 (
            .O(N__20638),
            .I(N__20635));
    Odrv4 I__2351 (
            .O(N__20635),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2350 (
            .O(N__20632),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__2349 (
            .O(N__20629),
            .I(N__20625));
    InMux I__2348 (
            .O(N__20628),
            .I(N__20621));
    LocalMux I__2347 (
            .O(N__20625),
            .I(N__20618));
    InMux I__2346 (
            .O(N__20624),
            .I(N__20615));
    LocalMux I__2345 (
            .O(N__20621),
            .I(N__20612));
    Span12Mux_s4_h I__2344 (
            .O(N__20618),
            .I(N__20607));
    LocalMux I__2343 (
            .O(N__20615),
            .I(N__20607));
    Span4Mux_h I__2342 (
            .O(N__20612),
            .I(N__20604));
    Odrv12 I__2341 (
            .O(N__20607),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__2340 (
            .O(N__20604),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2339 (
            .O(N__20599),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    CascadeMux I__2338 (
            .O(N__20596),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ));
    CascadeMux I__2337 (
            .O(N__20593),
            .I(N__20590));
    InMux I__2336 (
            .O(N__20590),
            .I(N__20586));
    InMux I__2335 (
            .O(N__20589),
            .I(N__20583));
    LocalMux I__2334 (
            .O(N__20586),
            .I(N__20580));
    LocalMux I__2333 (
            .O(N__20583),
            .I(N__20577));
    Span4Mux_h I__2332 (
            .O(N__20580),
            .I(N__20574));
    Odrv4 I__2331 (
            .O(N__20577),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    Odrv4 I__2330 (
            .O(N__20574),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__2329 (
            .O(N__20569),
            .I(N__20566));
    LocalMux I__2328 (
            .O(N__20566),
            .I(N__20562));
    InMux I__2327 (
            .O(N__20565),
            .I(N__20559));
    Odrv4 I__2326 (
            .O(N__20562),
            .I(clk_10khz_RNIIENAZ0Z2));
    LocalMux I__2325 (
            .O(N__20559),
            .I(clk_10khz_RNIIENAZ0Z2));
    InMux I__2324 (
            .O(N__20554),
            .I(N__20551));
    LocalMux I__2323 (
            .O(N__20551),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ));
    InMux I__2322 (
            .O(N__20548),
            .I(N__20545));
    LocalMux I__2321 (
            .O(N__20545),
            .I(N__20542));
    Glb2LocalMux I__2320 (
            .O(N__20542),
            .I(N__20539));
    GlobalMux I__2319 (
            .O(N__20539),
            .I(clk_12mhz));
    IoInMux I__2318 (
            .O(N__20536),
            .I(N__20533));
    LocalMux I__2317 (
            .O(N__20533),
            .I(N__20530));
    Span4Mux_s0_v I__2316 (
            .O(N__20530),
            .I(N__20527));
    Span4Mux_h I__2315 (
            .O(N__20527),
            .I(N__20524));
    Odrv4 I__2314 (
            .O(N__20524),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__2313 (
            .O(N__20521),
            .I(N__20518));
    LocalMux I__2312 (
            .O(N__20518),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    CascadeMux I__2311 (
            .O(N__20515),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_ ));
    InMux I__2310 (
            .O(N__20512),
            .I(N__20509));
    LocalMux I__2309 (
            .O(N__20509),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    CascadeMux I__2308 (
            .O(N__20506),
            .I(N__20503));
    InMux I__2307 (
            .O(N__20503),
            .I(N__20500));
    LocalMux I__2306 (
            .O(N__20500),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__2305 (
            .O(N__20497),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__2304 (
            .O(N__20494),
            .I(N__20491));
    LocalMux I__2303 (
            .O(N__20491),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__2302 (
            .O(N__20488),
            .I(N__20485));
    LocalMux I__2301 (
            .O(N__20485),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__2300 (
            .O(N__20482),
            .I(N__20479));
    LocalMux I__2299 (
            .O(N__20479),
            .I(N__20476));
    Odrv4 I__2298 (
            .O(N__20476),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    CascadeMux I__2297 (
            .O(N__20473),
            .I(N__20470));
    InMux I__2296 (
            .O(N__20470),
            .I(N__20467));
    LocalMux I__2295 (
            .O(N__20467),
            .I(N__20464));
    Odrv4 I__2294 (
            .O(N__20464),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__2293 (
            .O(N__20461),
            .I(N__20458));
    LocalMux I__2292 (
            .O(N__20458),
            .I(N__20455));
    Odrv4 I__2291 (
            .O(N__20455),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__2290 (
            .O(N__20452),
            .I(N__20449));
    LocalMux I__2289 (
            .O(N__20449),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__2288 (
            .O(N__20446),
            .I(N__20443));
    LocalMux I__2287 (
            .O(N__20443),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__2286 (
            .O(N__20440),
            .I(N__20437));
    LocalMux I__2285 (
            .O(N__20437),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__2284 (
            .O(N__20434),
            .I(N__20431));
    LocalMux I__2283 (
            .O(N__20431),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__2282 (
            .O(N__20428),
            .I(N__20425));
    LocalMux I__2281 (
            .O(N__20425),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__2280 (
            .O(N__20422),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    InMux I__2279 (
            .O(N__20419),
            .I(N__20416));
    LocalMux I__2278 (
            .O(N__20416),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    InMux I__2277 (
            .O(N__20413),
            .I(N__20410));
    LocalMux I__2276 (
            .O(N__20410),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    InMux I__2275 (
            .O(N__20407),
            .I(N__20404));
    LocalMux I__2274 (
            .O(N__20404),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__2273 (
            .O(N__20401),
            .I(N__20398));
    LocalMux I__2272 (
            .O(N__20398),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    CascadeMux I__2271 (
            .O(N__20395),
            .I(N__20392));
    InMux I__2270 (
            .O(N__20392),
            .I(N__20388));
    InMux I__2269 (
            .O(N__20391),
            .I(N__20385));
    LocalMux I__2268 (
            .O(N__20388),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    LocalMux I__2267 (
            .O(N__20385),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    InMux I__2266 (
            .O(N__20380),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    InMux I__2265 (
            .O(N__20377),
            .I(N__20374));
    LocalMux I__2264 (
            .O(N__20374),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    CascadeMux I__2263 (
            .O(N__20371),
            .I(N__20368));
    InMux I__2262 (
            .O(N__20368),
            .I(N__20365));
    LocalMux I__2261 (
            .O(N__20365),
            .I(N__20362));
    Span4Mux_s3_h I__2260 (
            .O(N__20362),
            .I(N__20359));
    Odrv4 I__2259 (
            .O(N__20359),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    InMux I__2258 (
            .O(N__20356),
            .I(bfn_3_13_0_));
    InMux I__2257 (
            .O(N__20353),
            .I(N__20350));
    LocalMux I__2256 (
            .O(N__20350),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__2255 (
            .O(N__20347),
            .I(N__20344));
    LocalMux I__2254 (
            .O(N__20344),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__2253 (
            .O(N__20341),
            .I(N__20338));
    LocalMux I__2252 (
            .O(N__20338),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    InMux I__2251 (
            .O(N__20335),
            .I(N__20332));
    LocalMux I__2250 (
            .O(N__20332),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__2249 (
            .O(N__20329),
            .I(N__20326));
    LocalMux I__2248 (
            .O(N__20326),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__2247 (
            .O(N__20323),
            .I(N__20320));
    LocalMux I__2246 (
            .O(N__20320),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__2245 (
            .O(N__20317),
            .I(N__20312));
    CascadeMux I__2244 (
            .O(N__20316),
            .I(N__20309));
    InMux I__2243 (
            .O(N__20315),
            .I(N__20306));
    LocalMux I__2242 (
            .O(N__20312),
            .I(N__20303));
    InMux I__2241 (
            .O(N__20309),
            .I(N__20300));
    LocalMux I__2240 (
            .O(N__20306),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    Odrv4 I__2239 (
            .O(N__20303),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__2238 (
            .O(N__20300),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    InMux I__2237 (
            .O(N__20293),
            .I(N__20289));
    InMux I__2236 (
            .O(N__20292),
            .I(N__20286));
    LocalMux I__2235 (
            .O(N__20289),
            .I(N__20283));
    LocalMux I__2234 (
            .O(N__20286),
            .I(N__20280));
    Span4Mux_v I__2233 (
            .O(N__20283),
            .I(N__20275));
    Span4Mux_v I__2232 (
            .O(N__20280),
            .I(N__20275));
    Odrv4 I__2231 (
            .O(N__20275),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__2230 (
            .O(N__20272),
            .I(N__20269));
    LocalMux I__2229 (
            .O(N__20269),
            .I(N__20266));
    Span4Mux_v I__2228 (
            .O(N__20266),
            .I(N__20263));
    Odrv4 I__2227 (
            .O(N__20263),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__2226 (
            .O(N__20260),
            .I(N__20257));
    LocalMux I__2225 (
            .O(N__20257),
            .I(N__20253));
    InMux I__2224 (
            .O(N__20256),
            .I(N__20250));
    Odrv4 I__2223 (
            .O(N__20253),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    LocalMux I__2222 (
            .O(N__20250),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    InMux I__2221 (
            .O(N__20245),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    CascadeMux I__2220 (
            .O(N__20242),
            .I(N__20239));
    InMux I__2219 (
            .O(N__20239),
            .I(N__20236));
    LocalMux I__2218 (
            .O(N__20236),
            .I(N__20233));
    Span4Mux_v I__2217 (
            .O(N__20233),
            .I(N__20230));
    Odrv4 I__2216 (
            .O(N__20230),
            .I(\pwm_generator_inst.O_13 ));
    CascadeMux I__2215 (
            .O(N__20227),
            .I(N__20224));
    InMux I__2214 (
            .O(N__20224),
            .I(N__20220));
    InMux I__2213 (
            .O(N__20223),
            .I(N__20217));
    LocalMux I__2212 (
            .O(N__20220),
            .I(N__20212));
    LocalMux I__2211 (
            .O(N__20217),
            .I(N__20212));
    Odrv4 I__2210 (
            .O(N__20212),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    InMux I__2209 (
            .O(N__20209),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__2208 (
            .O(N__20206),
            .I(N__20203));
    LocalMux I__2207 (
            .O(N__20203),
            .I(N__20200));
    Span4Mux_v I__2206 (
            .O(N__20200),
            .I(N__20197));
    Odrv4 I__2205 (
            .O(N__20197),
            .I(\pwm_generator_inst.O_14 ));
    CascadeMux I__2204 (
            .O(N__20194),
            .I(N__20191));
    InMux I__2203 (
            .O(N__20191),
            .I(N__20187));
    InMux I__2202 (
            .O(N__20190),
            .I(N__20184));
    LocalMux I__2201 (
            .O(N__20187),
            .I(N__20179));
    LocalMux I__2200 (
            .O(N__20184),
            .I(N__20179));
    Odrv4 I__2199 (
            .O(N__20179),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    InMux I__2198 (
            .O(N__20176),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    InMux I__2197 (
            .O(N__20173),
            .I(N__20170));
    LocalMux I__2196 (
            .O(N__20170),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    CascadeMux I__2195 (
            .O(N__20167),
            .I(N__20164));
    InMux I__2194 (
            .O(N__20164),
            .I(N__20161));
    LocalMux I__2193 (
            .O(N__20161),
            .I(N__20157));
    InMux I__2192 (
            .O(N__20160),
            .I(N__20154));
    Odrv4 I__2191 (
            .O(N__20157),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    LocalMux I__2190 (
            .O(N__20154),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    InMux I__2189 (
            .O(N__20149),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    CascadeMux I__2188 (
            .O(N__20146),
            .I(N__20143));
    InMux I__2187 (
            .O(N__20143),
            .I(N__20140));
    LocalMux I__2186 (
            .O(N__20140),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__2185 (
            .O(N__20137),
            .I(N__20131));
    InMux I__2184 (
            .O(N__20136),
            .I(N__20131));
    LocalMux I__2183 (
            .O(N__20131),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    InMux I__2182 (
            .O(N__20128),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    InMux I__2181 (
            .O(N__20125),
            .I(N__20122));
    LocalMux I__2180 (
            .O(N__20122),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__2179 (
            .O(N__20119),
            .I(N__20115));
    InMux I__2178 (
            .O(N__20118),
            .I(N__20112));
    LocalMux I__2177 (
            .O(N__20115),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    LocalMux I__2176 (
            .O(N__20112),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    InMux I__2175 (
            .O(N__20107),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    InMux I__2174 (
            .O(N__20104),
            .I(N__20099));
    InMux I__2173 (
            .O(N__20103),
            .I(N__20096));
    InMux I__2172 (
            .O(N__20102),
            .I(N__20093));
    LocalMux I__2171 (
            .O(N__20099),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__2170 (
            .O(N__20096),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__2169 (
            .O(N__20093),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    InMux I__2168 (
            .O(N__20086),
            .I(N__20083));
    LocalMux I__2167 (
            .O(N__20083),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    InMux I__2166 (
            .O(N__20080),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    InMux I__2165 (
            .O(N__20077),
            .I(N__20074));
    LocalMux I__2164 (
            .O(N__20074),
            .I(N__20071));
    Span4Mux_v I__2163 (
            .O(N__20071),
            .I(N__20068));
    Odrv4 I__2162 (
            .O(N__20068),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    InMux I__2161 (
            .O(N__20065),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    InMux I__2160 (
            .O(N__20062),
            .I(N__20058));
    InMux I__2159 (
            .O(N__20061),
            .I(N__20055));
    LocalMux I__2158 (
            .O(N__20058),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__2157 (
            .O(N__20055),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    InMux I__2156 (
            .O(N__20050),
            .I(N__20047));
    LocalMux I__2155 (
            .O(N__20047),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    InMux I__2154 (
            .O(N__20044),
            .I(bfn_3_11_0_));
    CascadeMux I__2153 (
            .O(N__20041),
            .I(N__20038));
    InMux I__2152 (
            .O(N__20038),
            .I(N__20035));
    LocalMux I__2151 (
            .O(N__20035),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    InMux I__2150 (
            .O(N__20032),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__2149 (
            .O(N__20029),
            .I(N__20026));
    LocalMux I__2148 (
            .O(N__20026),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    InMux I__2147 (
            .O(N__20023),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__2146 (
            .O(N__20020),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__2145 (
            .O(N__20017),
            .I(N__20014));
    LocalMux I__2144 (
            .O(N__20014),
            .I(N__20011));
    Odrv4 I__2143 (
            .O(N__20011),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    InMux I__2142 (
            .O(N__20008),
            .I(N__20004));
    InMux I__2141 (
            .O(N__20007),
            .I(N__20000));
    LocalMux I__2140 (
            .O(N__20004),
            .I(N__19997));
    InMux I__2139 (
            .O(N__20003),
            .I(N__19994));
    LocalMux I__2138 (
            .O(N__20000),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    Odrv4 I__2137 (
            .O(N__19997),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__2136 (
            .O(N__19994),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    InMux I__2135 (
            .O(N__19987),
            .I(N__19982));
    InMux I__2134 (
            .O(N__19986),
            .I(N__19977));
    InMux I__2133 (
            .O(N__19985),
            .I(N__19977));
    LocalMux I__2132 (
            .O(N__19982),
            .I(N__19974));
    LocalMux I__2131 (
            .O(N__19977),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    Odrv4 I__2130 (
            .O(N__19974),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__2129 (
            .O(N__19969),
            .I(N__19964));
    InMux I__2128 (
            .O(N__19968),
            .I(N__19959));
    InMux I__2127 (
            .O(N__19967),
            .I(N__19959));
    LocalMux I__2126 (
            .O(N__19964),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__2125 (
            .O(N__19959),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    InMux I__2124 (
            .O(N__19954),
            .I(N__19951));
    LocalMux I__2123 (
            .O(N__19951),
            .I(N__19948));
    Span4Mux_h I__2122 (
            .O(N__19948),
            .I(N__19945));
    Odrv4 I__2121 (
            .O(N__19945),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__2120 (
            .O(N__19942),
            .I(N__19939));
    LocalMux I__2119 (
            .O(N__19939),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    InMux I__2118 (
            .O(N__19936),
            .I(N__19933));
    LocalMux I__2117 (
            .O(N__19933),
            .I(N__19930));
    Span4Mux_v I__2116 (
            .O(N__19930),
            .I(N__19927));
    Odrv4 I__2115 (
            .O(N__19927),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__2114 (
            .O(N__19924),
            .I(N__19921));
    LocalMux I__2113 (
            .O(N__19921),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    InMux I__2112 (
            .O(N__19918),
            .I(N__19915));
    LocalMux I__2111 (
            .O(N__19915),
            .I(N__19912));
    Span4Mux_v I__2110 (
            .O(N__19912),
            .I(N__19909));
    Odrv4 I__2109 (
            .O(N__19909),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__2108 (
            .O(N__19906),
            .I(N__19903));
    LocalMux I__2107 (
            .O(N__19903),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__2106 (
            .O(N__19900),
            .I(N__19897));
    LocalMux I__2105 (
            .O(N__19897),
            .I(N__19892));
    InMux I__2104 (
            .O(N__19896),
            .I(N__19889));
    InMux I__2103 (
            .O(N__19895),
            .I(N__19886));
    Span4Mux_h I__2102 (
            .O(N__19892),
            .I(N__19883));
    LocalMux I__2101 (
            .O(N__19889),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    LocalMux I__2100 (
            .O(N__19886),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    Odrv4 I__2099 (
            .O(N__19883),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    CascadeMux I__2098 (
            .O(N__19876),
            .I(N__19873));
    InMux I__2097 (
            .O(N__19873),
            .I(N__19870));
    LocalMux I__2096 (
            .O(N__19870),
            .I(N__19867));
    Span4Mux_v I__2095 (
            .O(N__19867),
            .I(N__19864));
    Odrv4 I__2094 (
            .O(N__19864),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    InMux I__2093 (
            .O(N__19861),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    CascadeMux I__2092 (
            .O(N__19858),
            .I(N__19854));
    InMux I__2091 (
            .O(N__19857),
            .I(N__19842));
    InMux I__2090 (
            .O(N__19854),
            .I(N__19839));
    InMux I__2089 (
            .O(N__19853),
            .I(N__19828));
    InMux I__2088 (
            .O(N__19852),
            .I(N__19828));
    InMux I__2087 (
            .O(N__19851),
            .I(N__19828));
    InMux I__2086 (
            .O(N__19850),
            .I(N__19828));
    InMux I__2085 (
            .O(N__19849),
            .I(N__19828));
    InMux I__2084 (
            .O(N__19848),
            .I(N__19825));
    InMux I__2083 (
            .O(N__19847),
            .I(N__19818));
    InMux I__2082 (
            .O(N__19846),
            .I(N__19818));
    InMux I__2081 (
            .O(N__19845),
            .I(N__19818));
    LocalMux I__2080 (
            .O(N__19842),
            .I(N__19811));
    LocalMux I__2079 (
            .O(N__19839),
            .I(N__19811));
    LocalMux I__2078 (
            .O(N__19828),
            .I(N__19811));
    LocalMux I__2077 (
            .O(N__19825),
            .I(N__19807));
    LocalMux I__2076 (
            .O(N__19818),
            .I(N__19802));
    Span4Mux_v I__2075 (
            .O(N__19811),
            .I(N__19802));
    InMux I__2074 (
            .O(N__19810),
            .I(N__19799));
    Span4Mux_v I__2073 (
            .O(N__19807),
            .I(N__19796));
    Odrv4 I__2072 (
            .O(N__19802),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2071 (
            .O(N__19799),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2070 (
            .O(N__19796),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    InMux I__2069 (
            .O(N__19789),
            .I(N__19786));
    LocalMux I__2068 (
            .O(N__19786),
            .I(N__19783));
    Odrv4 I__2067 (
            .O(N__19783),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    InMux I__2066 (
            .O(N__19780),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    CascadeMux I__2065 (
            .O(N__19777),
            .I(N__19774));
    InMux I__2064 (
            .O(N__19774),
            .I(N__19771));
    LocalMux I__2063 (
            .O(N__19771),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    InMux I__2062 (
            .O(N__19768),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    CascadeMux I__2061 (
            .O(N__19765),
            .I(N__19760));
    InMux I__2060 (
            .O(N__19764),
            .I(N__19757));
    InMux I__2059 (
            .O(N__19763),
            .I(N__19754));
    InMux I__2058 (
            .O(N__19760),
            .I(N__19751));
    LocalMux I__2057 (
            .O(N__19757),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    LocalMux I__2056 (
            .O(N__19754),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    LocalMux I__2055 (
            .O(N__19751),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    InMux I__2054 (
            .O(N__19744),
            .I(N__19741));
    LocalMux I__2053 (
            .O(N__19741),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    InMux I__2052 (
            .O(N__19738),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__2051 (
            .O(N__19735),
            .I(N__19722));
    InMux I__2050 (
            .O(N__19734),
            .I(N__19722));
    InMux I__2049 (
            .O(N__19733),
            .I(N__19717));
    InMux I__2048 (
            .O(N__19732),
            .I(N__19717));
    InMux I__2047 (
            .O(N__19731),
            .I(N__19706));
    InMux I__2046 (
            .O(N__19730),
            .I(N__19706));
    InMux I__2045 (
            .O(N__19729),
            .I(N__19706));
    InMux I__2044 (
            .O(N__19728),
            .I(N__19706));
    InMux I__2043 (
            .O(N__19727),
            .I(N__19706));
    LocalMux I__2042 (
            .O(N__19722),
            .I(N__19699));
    LocalMux I__2041 (
            .O(N__19717),
            .I(N__19699));
    LocalMux I__2040 (
            .O(N__19706),
            .I(N__19696));
    InMux I__2039 (
            .O(N__19705),
            .I(N__19693));
    InMux I__2038 (
            .O(N__19704),
            .I(N__19690));
    Span4Mux_h I__2037 (
            .O(N__19699),
            .I(N__19687));
    Span4Mux_h I__2036 (
            .O(N__19696),
            .I(N__19684));
    LocalMux I__2035 (
            .O(N__19693),
            .I(N__19681));
    LocalMux I__2034 (
            .O(N__19690),
            .I(pwm_duty_input_6));
    Odrv4 I__2033 (
            .O(N__19687),
            .I(pwm_duty_input_6));
    Odrv4 I__2032 (
            .O(N__19684),
            .I(pwm_duty_input_6));
    Odrv4 I__2031 (
            .O(N__19681),
            .I(pwm_duty_input_6));
    CascadeMux I__2030 (
            .O(N__19672),
            .I(N__19666));
    CascadeMux I__2029 (
            .O(N__19671),
            .I(N__19663));
    CascadeMux I__2028 (
            .O(N__19670),
            .I(N__19660));
    InMux I__2027 (
            .O(N__19669),
            .I(N__19649));
    InMux I__2026 (
            .O(N__19666),
            .I(N__19649));
    InMux I__2025 (
            .O(N__19663),
            .I(N__19644));
    InMux I__2024 (
            .O(N__19660),
            .I(N__19644));
    InMux I__2023 (
            .O(N__19659),
            .I(N__19641));
    InMux I__2022 (
            .O(N__19658),
            .I(N__19630));
    InMux I__2021 (
            .O(N__19657),
            .I(N__19630));
    InMux I__2020 (
            .O(N__19656),
            .I(N__19630));
    InMux I__2019 (
            .O(N__19655),
            .I(N__19630));
    InMux I__2018 (
            .O(N__19654),
            .I(N__19630));
    LocalMux I__2017 (
            .O(N__19649),
            .I(N__19627));
    LocalMux I__2016 (
            .O(N__19644),
            .I(N__19624));
    LocalMux I__2015 (
            .O(N__19641),
            .I(i8_mux));
    LocalMux I__2014 (
            .O(N__19630),
            .I(i8_mux));
    Odrv4 I__2013 (
            .O(N__19627),
            .I(i8_mux));
    Odrv4 I__2012 (
            .O(N__19624),
            .I(i8_mux));
    CascadeMux I__2011 (
            .O(N__19615),
            .I(N__19604));
    CascadeMux I__2010 (
            .O(N__19614),
            .I(N__19601));
    CascadeMux I__2009 (
            .O(N__19613),
            .I(N__19598));
    CascadeMux I__2008 (
            .O(N__19612),
            .I(N__19595));
    CascadeMux I__2007 (
            .O(N__19611),
            .I(N__19592));
    InMux I__2006 (
            .O(N__19610),
            .I(N__19587));
    InMux I__2005 (
            .O(N__19609),
            .I(N__19587));
    InMux I__2004 (
            .O(N__19608),
            .I(N__19582));
    InMux I__2003 (
            .O(N__19607),
            .I(N__19582));
    InMux I__2002 (
            .O(N__19604),
            .I(N__19574));
    InMux I__2001 (
            .O(N__19601),
            .I(N__19574));
    InMux I__2000 (
            .O(N__19598),
            .I(N__19574));
    InMux I__1999 (
            .O(N__19595),
            .I(N__19569));
    InMux I__1998 (
            .O(N__19592),
            .I(N__19569));
    LocalMux I__1997 (
            .O(N__19587),
            .I(N__19564));
    LocalMux I__1996 (
            .O(N__19582),
            .I(N__19564));
    InMux I__1995 (
            .O(N__19581),
            .I(N__19561));
    LocalMux I__1994 (
            .O(N__19574),
            .I(N__19556));
    LocalMux I__1993 (
            .O(N__19569),
            .I(N__19556));
    Span4Mux_h I__1992 (
            .O(N__19564),
            .I(N__19553));
    LocalMux I__1991 (
            .O(N__19561),
            .I(N__19548));
    Span4Mux_h I__1990 (
            .O(N__19556),
            .I(N__19548));
    Span4Mux_v I__1989 (
            .O(N__19553),
            .I(N__19545));
    Odrv4 I__1988 (
            .O(N__19548),
            .I(N_28_mux));
    Odrv4 I__1987 (
            .O(N__19545),
            .I(N_28_mux));
    InMux I__1986 (
            .O(N__19540),
            .I(N__19537));
    LocalMux I__1985 (
            .O(N__19537),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    InMux I__1984 (
            .O(N__19534),
            .I(N__19531));
    LocalMux I__1983 (
            .O(N__19531),
            .I(N__19528));
    Span4Mux_v I__1982 (
            .O(N__19528),
            .I(N__19525));
    Odrv4 I__1981 (
            .O(N__19525),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1980 (
            .O(N__19522),
            .I(N__19519));
    LocalMux I__1979 (
            .O(N__19519),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__1978 (
            .O(N__19516),
            .I(N__19513));
    LocalMux I__1977 (
            .O(N__19513),
            .I(N__19510));
    Span4Mux_v I__1976 (
            .O(N__19510),
            .I(N__19507));
    Odrv4 I__1975 (
            .O(N__19507),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1974 (
            .O(N__19504),
            .I(N__19501));
    LocalMux I__1973 (
            .O(N__19501),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__1972 (
            .O(N__19498),
            .I(N__19495));
    LocalMux I__1971 (
            .O(N__19495),
            .I(N__19492));
    Span4Mux_h I__1970 (
            .O(N__19492),
            .I(N__19489));
    Odrv4 I__1969 (
            .O(N__19489),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1968 (
            .O(N__19486),
            .I(N__19483));
    LocalMux I__1967 (
            .O(N__19483),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    InMux I__1966 (
            .O(N__19480),
            .I(N__19477));
    LocalMux I__1965 (
            .O(N__19477),
            .I(N__19474));
    Span4Mux_h I__1964 (
            .O(N__19474),
            .I(N__19471));
    Odrv4 I__1963 (
            .O(N__19471),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1962 (
            .O(N__19468),
            .I(N__19465));
    LocalMux I__1961 (
            .O(N__19465),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__1960 (
            .O(N__19462),
            .I(N__19459));
    LocalMux I__1959 (
            .O(N__19459),
            .I(N__19456));
    Span4Mux_h I__1958 (
            .O(N__19456),
            .I(N__19453));
    Odrv4 I__1957 (
            .O(N__19453),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1956 (
            .O(N__19450),
            .I(N__19447));
    LocalMux I__1955 (
            .O(N__19447),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__1954 (
            .O(N__19444),
            .I(N__19441));
    LocalMux I__1953 (
            .O(N__19441),
            .I(N__19438));
    Span4Mux_h I__1952 (
            .O(N__19438),
            .I(N__19435));
    Odrv4 I__1951 (
            .O(N__19435),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1950 (
            .O(N__19432),
            .I(N__19429));
    LocalMux I__1949 (
            .O(N__19429),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__1948 (
            .O(N__19426),
            .I(N__19423));
    LocalMux I__1947 (
            .O(N__19423),
            .I(N__19420));
    Span4Mux_h I__1946 (
            .O(N__19420),
            .I(N__19417));
    Odrv4 I__1945 (
            .O(N__19417),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1944 (
            .O(N__19414),
            .I(N__19411));
    LocalMux I__1943 (
            .O(N__19411),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    InMux I__1942 (
            .O(N__19408),
            .I(N__19405));
    LocalMux I__1941 (
            .O(N__19405),
            .I(N__19402));
    Span4Mux_s2_v I__1940 (
            .O(N__19402),
            .I(N__19399));
    Odrv4 I__1939 (
            .O(N__19399),
            .I(N_22_i_i));
    InMux I__1938 (
            .O(N__19396),
            .I(N__19393));
    LocalMux I__1937 (
            .O(N__19393),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    CascadeMux I__1936 (
            .O(N__19390),
            .I(N__19387));
    InMux I__1935 (
            .O(N__19387),
            .I(N__19384));
    LocalMux I__1934 (
            .O(N__19384),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__1933 (
            .O(N__19381),
            .I(N__19378));
    LocalMux I__1932 (
            .O(N__19378),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    InMux I__1931 (
            .O(N__19375),
            .I(N__19372));
    LocalMux I__1930 (
            .O(N__19372),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    InMux I__1929 (
            .O(N__19369),
            .I(N__19366));
    LocalMux I__1928 (
            .O(N__19366),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    InMux I__1927 (
            .O(N__19363),
            .I(N__19360));
    LocalMux I__1926 (
            .O(N__19360),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    InMux I__1925 (
            .O(N__19357),
            .I(N__19354));
    LocalMux I__1924 (
            .O(N__19354),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    InMux I__1923 (
            .O(N__19351),
            .I(N__19348));
    LocalMux I__1922 (
            .O(N__19348),
            .I(N__19344));
    InMux I__1921 (
            .O(N__19347),
            .I(N__19341));
    Span4Mux_h I__1920 (
            .O(N__19344),
            .I(N__19336));
    LocalMux I__1919 (
            .O(N__19341),
            .I(N__19336));
    Odrv4 I__1918 (
            .O(N__19336),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__1917 (
            .O(N__19333),
            .I(N__19330));
    LocalMux I__1916 (
            .O(N__19330),
            .I(N__19327));
    Odrv12 I__1915 (
            .O(N__19327),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    InMux I__1914 (
            .O(N__19324),
            .I(N__19321));
    LocalMux I__1913 (
            .O(N__19321),
            .I(N__19318));
    Span4Mux_v I__1912 (
            .O(N__19318),
            .I(N__19314));
    InMux I__1911 (
            .O(N__19317),
            .I(N__19311));
    Odrv4 I__1910 (
            .O(N__19314),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    LocalMux I__1909 (
            .O(N__19311),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    CascadeMux I__1908 (
            .O(N__19306),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__1907 (
            .O(N__19303),
            .I(N__19300));
    LocalMux I__1906 (
            .O(N__19300),
            .I(N__19295));
    InMux I__1905 (
            .O(N__19299),
            .I(N__19292));
    InMux I__1904 (
            .O(N__19298),
            .I(N__19289));
    Odrv4 I__1903 (
            .O(N__19295),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__1902 (
            .O(N__19292),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__1901 (
            .O(N__19289),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__1900 (
            .O(N__19282),
            .I(N__19278));
    InMux I__1899 (
            .O(N__19281),
            .I(N__19271));
    LocalMux I__1898 (
            .O(N__19278),
            .I(N__19268));
    InMux I__1897 (
            .O(N__19277),
            .I(N__19259));
    InMux I__1896 (
            .O(N__19276),
            .I(N__19259));
    InMux I__1895 (
            .O(N__19275),
            .I(N__19259));
    InMux I__1894 (
            .O(N__19274),
            .I(N__19259));
    LocalMux I__1893 (
            .O(N__19271),
            .I(N__19251));
    Span4Mux_s2_h I__1892 (
            .O(N__19268),
            .I(N__19251));
    LocalMux I__1891 (
            .O(N__19259),
            .I(N__19251));
    InMux I__1890 (
            .O(N__19258),
            .I(N__19248));
    Span4Mux_v I__1889 (
            .O(N__19251),
            .I(N__19243));
    LocalMux I__1888 (
            .O(N__19248),
            .I(N__19243));
    Odrv4 I__1887 (
            .O(N__19243),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    CascadeMux I__1886 (
            .O(N__19240),
            .I(N__19236));
    InMux I__1885 (
            .O(N__19239),
            .I(N__19229));
    InMux I__1884 (
            .O(N__19236),
            .I(N__19218));
    InMux I__1883 (
            .O(N__19235),
            .I(N__19218));
    InMux I__1882 (
            .O(N__19234),
            .I(N__19218));
    InMux I__1881 (
            .O(N__19233),
            .I(N__19218));
    InMux I__1880 (
            .O(N__19232),
            .I(N__19218));
    LocalMux I__1879 (
            .O(N__19229),
            .I(N__19213));
    LocalMux I__1878 (
            .O(N__19218),
            .I(N__19210));
    InMux I__1877 (
            .O(N__19217),
            .I(N__19207));
    InMux I__1876 (
            .O(N__19216),
            .I(N__19204));
    Span4Mux_v I__1875 (
            .O(N__19213),
            .I(N__19194));
    Span4Mux_s2_h I__1874 (
            .O(N__19210),
            .I(N__19194));
    LocalMux I__1873 (
            .O(N__19207),
            .I(N__19194));
    LocalMux I__1872 (
            .O(N__19204),
            .I(N__19194));
    InMux I__1871 (
            .O(N__19203),
            .I(N__19191));
    Span4Mux_v I__1870 (
            .O(N__19194),
            .I(N__19186));
    LocalMux I__1869 (
            .O(N__19191),
            .I(N__19186));
    Odrv4 I__1868 (
            .O(N__19186),
            .I(\current_shift_inst.PI_CTRL.N_178 ));
    CascadeMux I__1867 (
            .O(N__19183),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ));
    InMux I__1866 (
            .O(N__19180),
            .I(N__19177));
    LocalMux I__1865 (
            .O(N__19177),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__1864 (
            .O(N__19174),
            .I(N__19171));
    LocalMux I__1863 (
            .O(N__19171),
            .I(N__19168));
    Span4Mux_h I__1862 (
            .O(N__19168),
            .I(N__19165));
    Span4Mux_v I__1861 (
            .O(N__19165),
            .I(N__19162));
    Odrv4 I__1860 (
            .O(N__19162),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    InMux I__1859 (
            .O(N__19159),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    CascadeMux I__1858 (
            .O(N__19156),
            .I(N__19153));
    InMux I__1857 (
            .O(N__19153),
            .I(N__19150));
    LocalMux I__1856 (
            .O(N__19150),
            .I(N__19147));
    Span4Mux_h I__1855 (
            .O(N__19147),
            .I(N__19144));
    Span4Mux_v I__1854 (
            .O(N__19144),
            .I(N__19141));
    Odrv4 I__1853 (
            .O(N__19141),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1852 (
            .O(N__19138),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    InMux I__1851 (
            .O(N__19135),
            .I(N__19132));
    LocalMux I__1850 (
            .O(N__19132),
            .I(N__19129));
    Span4Mux_h I__1849 (
            .O(N__19129),
            .I(N__19126));
    Span4Mux_v I__1848 (
            .O(N__19126),
            .I(N__19123));
    Odrv4 I__1847 (
            .O(N__19123),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    InMux I__1846 (
            .O(N__19120),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    CascadeMux I__1845 (
            .O(N__19117),
            .I(N__19114));
    InMux I__1844 (
            .O(N__19114),
            .I(N__19111));
    LocalMux I__1843 (
            .O(N__19111),
            .I(N__19108));
    Span4Mux_h I__1842 (
            .O(N__19108),
            .I(N__19105));
    Span4Mux_v I__1841 (
            .O(N__19105),
            .I(N__19102));
    Odrv4 I__1840 (
            .O(N__19102),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__1839 (
            .O(N__19099),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    InMux I__1838 (
            .O(N__19096),
            .I(N__19093));
    LocalMux I__1837 (
            .O(N__19093),
            .I(N__19090));
    Span4Mux_v I__1836 (
            .O(N__19090),
            .I(N__19087));
    Span4Mux_v I__1835 (
            .O(N__19087),
            .I(N__19084));
    Odrv4 I__1834 (
            .O(N__19084),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    InMux I__1833 (
            .O(N__19081),
            .I(N__19078));
    LocalMux I__1832 (
            .O(N__19078),
            .I(N__19071));
    InMux I__1831 (
            .O(N__19077),
            .I(N__19068));
    CascadeMux I__1830 (
            .O(N__19076),
            .I(N__19065));
    CascadeMux I__1829 (
            .O(N__19075),
            .I(N__19061));
    CascadeMux I__1828 (
            .O(N__19074),
            .I(N__19057));
    Span4Mux_v I__1827 (
            .O(N__19071),
            .I(N__19051));
    LocalMux I__1826 (
            .O(N__19068),
            .I(N__19051));
    InMux I__1825 (
            .O(N__19065),
            .I(N__19038));
    InMux I__1824 (
            .O(N__19064),
            .I(N__19038));
    InMux I__1823 (
            .O(N__19061),
            .I(N__19038));
    InMux I__1822 (
            .O(N__19060),
            .I(N__19038));
    InMux I__1821 (
            .O(N__19057),
            .I(N__19038));
    InMux I__1820 (
            .O(N__19056),
            .I(N__19038));
    Span4Mux_v I__1819 (
            .O(N__19051),
            .I(N__19035));
    LocalMux I__1818 (
            .O(N__19038),
            .I(N__19032));
    Odrv4 I__1817 (
            .O(N__19035),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    Odrv4 I__1816 (
            .O(N__19032),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    InMux I__1815 (
            .O(N__19027),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__1814 (
            .O(N__19024),
            .I(N__19021));
    LocalMux I__1813 (
            .O(N__19021),
            .I(N__19018));
    Span4Mux_v I__1812 (
            .O(N__19018),
            .I(N__19015));
    Odrv4 I__1811 (
            .O(N__19015),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    InMux I__1810 (
            .O(N__19012),
            .I(bfn_2_14_0_));
    InMux I__1809 (
            .O(N__19009),
            .I(N__19006));
    LocalMux I__1808 (
            .O(N__19006),
            .I(N__19001));
    InMux I__1807 (
            .O(N__19005),
            .I(N__18996));
    InMux I__1806 (
            .O(N__19004),
            .I(N__18996));
    Span4Mux_s2_h I__1805 (
            .O(N__19001),
            .I(N__18991));
    LocalMux I__1804 (
            .O(N__18996),
            .I(N__18991));
    Odrv4 I__1803 (
            .O(N__18991),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1802 (
            .O(N__18988),
            .I(N__18985));
    LocalMux I__1801 (
            .O(N__18985),
            .I(\current_shift_inst.PI_CTRL.N_98 ));
    InMux I__1800 (
            .O(N__18982),
            .I(N__18976));
    InMux I__1799 (
            .O(N__18981),
            .I(N__18976));
    LocalMux I__1798 (
            .O(N__18976),
            .I(N__18971));
    InMux I__1797 (
            .O(N__18975),
            .I(N__18966));
    InMux I__1796 (
            .O(N__18974),
            .I(N__18966));
    Span4Mux_s2_h I__1795 (
            .O(N__18971),
            .I(N__18960));
    LocalMux I__1794 (
            .O(N__18966),
            .I(N__18960));
    InMux I__1793 (
            .O(N__18965),
            .I(N__18957));
    Odrv4 I__1792 (
            .O(N__18960),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    LocalMux I__1791 (
            .O(N__18957),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    InMux I__1790 (
            .O(N__18952),
            .I(N__18949));
    LocalMux I__1789 (
            .O(N__18949),
            .I(N__18946));
    Odrv4 I__1788 (
            .O(N__18946),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    CascadeMux I__1787 (
            .O(N__18943),
            .I(N__18940));
    InMux I__1786 (
            .O(N__18940),
            .I(N__18937));
    LocalMux I__1785 (
            .O(N__18937),
            .I(N__18934));
    Span4Mux_h I__1784 (
            .O(N__18934),
            .I(N__18931));
    Span4Mux_v I__1783 (
            .O(N__18931),
            .I(N__18928));
    Odrv4 I__1782 (
            .O(N__18928),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    InMux I__1781 (
            .O(N__18925),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1780 (
            .O(N__18922),
            .I(N__18919));
    LocalMux I__1779 (
            .O(N__18919),
            .I(N__18916));
    Odrv4 I__1778 (
            .O(N__18916),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    CascadeMux I__1777 (
            .O(N__18913),
            .I(N__18910));
    InMux I__1776 (
            .O(N__18910),
            .I(N__18907));
    LocalMux I__1775 (
            .O(N__18907),
            .I(N__18904));
    Span4Mux_h I__1774 (
            .O(N__18904),
            .I(N__18901));
    Span4Mux_v I__1773 (
            .O(N__18901),
            .I(N__18898));
    Odrv4 I__1772 (
            .O(N__18898),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    InMux I__1771 (
            .O(N__18895),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1770 (
            .O(N__18892),
            .I(N__18889));
    LocalMux I__1769 (
            .O(N__18889),
            .I(N__18886));
    Span4Mux_h I__1768 (
            .O(N__18886),
            .I(N__18883));
    Span4Mux_v I__1767 (
            .O(N__18883),
            .I(N__18880));
    Odrv4 I__1766 (
            .O(N__18880),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    CascadeMux I__1765 (
            .O(N__18877),
            .I(N__18874));
    InMux I__1764 (
            .O(N__18874),
            .I(N__18871));
    LocalMux I__1763 (
            .O(N__18871),
            .I(N__18868));
    Odrv4 I__1762 (
            .O(N__18868),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    InMux I__1761 (
            .O(N__18865),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__1760 (
            .O(N__18862),
            .I(N__18859));
    LocalMux I__1759 (
            .O(N__18859),
            .I(N__18856));
    Span4Mux_h I__1758 (
            .O(N__18856),
            .I(N__18853));
    Span4Mux_v I__1757 (
            .O(N__18853),
            .I(N__18850));
    Odrv4 I__1756 (
            .O(N__18850),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    CascadeMux I__1755 (
            .O(N__18847),
            .I(N__18844));
    InMux I__1754 (
            .O(N__18844),
            .I(N__18841));
    LocalMux I__1753 (
            .O(N__18841),
            .I(N__18838));
    Odrv4 I__1752 (
            .O(N__18838),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    InMux I__1751 (
            .O(N__18835),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__1750 (
            .O(N__18832),
            .I(N__18829));
    LocalMux I__1749 (
            .O(N__18829),
            .I(N__18826));
    Span4Mux_v I__1748 (
            .O(N__18826),
            .I(N__18823));
    Span4Mux_v I__1747 (
            .O(N__18823),
            .I(N__18820));
    Odrv4 I__1746 (
            .O(N__18820),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    CascadeMux I__1745 (
            .O(N__18817),
            .I(N__18814));
    InMux I__1744 (
            .O(N__18814),
            .I(N__18811));
    LocalMux I__1743 (
            .O(N__18811),
            .I(N__18808));
    Odrv4 I__1742 (
            .O(N__18808),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    InMux I__1741 (
            .O(N__18805),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__1740 (
            .O(N__18802),
            .I(N__18799));
    LocalMux I__1739 (
            .O(N__18799),
            .I(N__18796));
    Span4Mux_h I__1738 (
            .O(N__18796),
            .I(N__18793));
    Odrv4 I__1737 (
            .O(N__18793),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    CascadeMux I__1736 (
            .O(N__18790),
            .I(N__18787));
    InMux I__1735 (
            .O(N__18787),
            .I(N__18784));
    LocalMux I__1734 (
            .O(N__18784),
            .I(N__18781));
    Span4Mux_v I__1733 (
            .O(N__18781),
            .I(N__18778));
    Span4Mux_v I__1732 (
            .O(N__18778),
            .I(N__18775));
    Odrv4 I__1731 (
            .O(N__18775),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    InMux I__1730 (
            .O(N__18772),
            .I(bfn_2_13_0_));
    InMux I__1729 (
            .O(N__18769),
            .I(N__18766));
    LocalMux I__1728 (
            .O(N__18766),
            .I(N__18763));
    Odrv4 I__1727 (
            .O(N__18763),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    CascadeMux I__1726 (
            .O(N__18760),
            .I(N__18757));
    InMux I__1725 (
            .O(N__18757),
            .I(N__18754));
    LocalMux I__1724 (
            .O(N__18754),
            .I(N__18751));
    Span4Mux_v I__1723 (
            .O(N__18751),
            .I(N__18748));
    Span4Mux_v I__1722 (
            .O(N__18748),
            .I(N__18745));
    Odrv4 I__1721 (
            .O(N__18745),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    InMux I__1720 (
            .O(N__18742),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    CascadeMux I__1719 (
            .O(N__18739),
            .I(N__18736));
    InMux I__1718 (
            .O(N__18736),
            .I(N__18733));
    LocalMux I__1717 (
            .O(N__18733),
            .I(N__18730));
    Span4Mux_h I__1716 (
            .O(N__18730),
            .I(N__18727));
    Span4Mux_v I__1715 (
            .O(N__18727),
            .I(N__18724));
    Odrv4 I__1714 (
            .O(N__18724),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1713 (
            .O(N__18721),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    CascadeMux I__1712 (
            .O(N__18718),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ));
    InMux I__1711 (
            .O(N__18715),
            .I(N__18712));
    LocalMux I__1710 (
            .O(N__18712),
            .I(N__18709));
    Odrv4 I__1709 (
            .O(N__18709),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    InMux I__1708 (
            .O(N__18706),
            .I(N__18703));
    LocalMux I__1707 (
            .O(N__18703),
            .I(N__18700));
    Odrv4 I__1706 (
            .O(N__18700),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    CascadeMux I__1705 (
            .O(N__18697),
            .I(N__18694));
    InMux I__1704 (
            .O(N__18694),
            .I(N__18691));
    LocalMux I__1703 (
            .O(N__18691),
            .I(N__18688));
    Odrv4 I__1702 (
            .O(N__18688),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    InMux I__1701 (
            .O(N__18685),
            .I(N__18682));
    LocalMux I__1700 (
            .O(N__18682),
            .I(N__18679));
    Span4Mux_v I__1699 (
            .O(N__18679),
            .I(N__18676));
    Span4Mux_v I__1698 (
            .O(N__18676),
            .I(N__18673));
    Odrv4 I__1697 (
            .O(N__18673),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1696 (
            .O(N__18670),
            .I(N__18667));
    InMux I__1695 (
            .O(N__18667),
            .I(N__18664));
    LocalMux I__1694 (
            .O(N__18664),
            .I(N__18661));
    Span4Mux_h I__1693 (
            .O(N__18661),
            .I(N__18658));
    Odrv4 I__1692 (
            .O(N__18658),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    InMux I__1691 (
            .O(N__18655),
            .I(N__18652));
    LocalMux I__1690 (
            .O(N__18652),
            .I(N__18649));
    Odrv4 I__1689 (
            .O(N__18649),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    CascadeMux I__1688 (
            .O(N__18646),
            .I(N__18643));
    InMux I__1687 (
            .O(N__18643),
            .I(N__18640));
    LocalMux I__1686 (
            .O(N__18640),
            .I(N__18637));
    Span4Mux_v I__1685 (
            .O(N__18637),
            .I(N__18634));
    Span4Mux_v I__1684 (
            .O(N__18634),
            .I(N__18631));
    Odrv4 I__1683 (
            .O(N__18631),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    InMux I__1682 (
            .O(N__18628),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1681 (
            .O(N__18625),
            .I(N__18622));
    LocalMux I__1680 (
            .O(N__18622),
            .I(N__18619));
    Odrv4 I__1679 (
            .O(N__18619),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    CascadeMux I__1678 (
            .O(N__18616),
            .I(N__18613));
    InMux I__1677 (
            .O(N__18613),
            .I(N__18610));
    LocalMux I__1676 (
            .O(N__18610),
            .I(N__18607));
    Span4Mux_h I__1675 (
            .O(N__18607),
            .I(N__18604));
    Span4Mux_v I__1674 (
            .O(N__18604),
            .I(N__18601));
    Odrv4 I__1673 (
            .O(N__18601),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    InMux I__1672 (
            .O(N__18598),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1671 (
            .O(N__18595),
            .I(bfn_2_9_0_));
    InMux I__1670 (
            .O(N__18592),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    InMux I__1669 (
            .O(N__18589),
            .I(N__18586));
    LocalMux I__1668 (
            .O(N__18586),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    CascadeMux I__1667 (
            .O(N__18583),
            .I(N__18579));
    InMux I__1666 (
            .O(N__18582),
            .I(N__18576));
    InMux I__1665 (
            .O(N__18579),
            .I(N__18572));
    LocalMux I__1664 (
            .O(N__18576),
            .I(N__18569));
    InMux I__1663 (
            .O(N__18575),
            .I(N__18566));
    LocalMux I__1662 (
            .O(N__18572),
            .I(N__18563));
    Span4Mux_s1_h I__1661 (
            .O(N__18569),
            .I(N__18560));
    LocalMux I__1660 (
            .O(N__18566),
            .I(pwm_duty_input_8));
    Odrv4 I__1659 (
            .O(N__18563),
            .I(pwm_duty_input_8));
    Odrv4 I__1658 (
            .O(N__18560),
            .I(pwm_duty_input_8));
    InMux I__1657 (
            .O(N__18553),
            .I(N__18524));
    InMux I__1656 (
            .O(N__18552),
            .I(N__18524));
    InMux I__1655 (
            .O(N__18551),
            .I(N__18524));
    InMux I__1654 (
            .O(N__18550),
            .I(N__18524));
    InMux I__1653 (
            .O(N__18549),
            .I(N__18524));
    InMux I__1652 (
            .O(N__18548),
            .I(N__18524));
    InMux I__1651 (
            .O(N__18547),
            .I(N__18524));
    InMux I__1650 (
            .O(N__18546),
            .I(N__18524));
    InMux I__1649 (
            .O(N__18545),
            .I(N__18519));
    InMux I__1648 (
            .O(N__18544),
            .I(N__18519));
    InMux I__1647 (
            .O(N__18543),
            .I(N__18513));
    CascadeMux I__1646 (
            .O(N__18542),
            .I(N__18510));
    InMux I__1645 (
            .O(N__18541),
            .I(N__18507));
    LocalMux I__1644 (
            .O(N__18524),
            .I(N__18504));
    LocalMux I__1643 (
            .O(N__18519),
            .I(N__18501));
    InMux I__1642 (
            .O(N__18518),
            .I(N__18494));
    InMux I__1641 (
            .O(N__18517),
            .I(N__18494));
    InMux I__1640 (
            .O(N__18516),
            .I(N__18494));
    LocalMux I__1639 (
            .O(N__18513),
            .I(N__18491));
    InMux I__1638 (
            .O(N__18510),
            .I(N__18488));
    LocalMux I__1637 (
            .O(N__18507),
            .I(N__18471));
    Span4Mux_v I__1636 (
            .O(N__18504),
            .I(N__18471));
    Span4Mux_s1_h I__1635 (
            .O(N__18501),
            .I(N__18471));
    LocalMux I__1634 (
            .O(N__18494),
            .I(N__18471));
    Span4Mux_v I__1633 (
            .O(N__18491),
            .I(N__18466));
    LocalMux I__1632 (
            .O(N__18488),
            .I(N__18466));
    InMux I__1631 (
            .O(N__18487),
            .I(N__18463));
    InMux I__1630 (
            .O(N__18486),
            .I(N__18448));
    InMux I__1629 (
            .O(N__18485),
            .I(N__18448));
    InMux I__1628 (
            .O(N__18484),
            .I(N__18448));
    InMux I__1627 (
            .O(N__18483),
            .I(N__18448));
    InMux I__1626 (
            .O(N__18482),
            .I(N__18448));
    InMux I__1625 (
            .O(N__18481),
            .I(N__18448));
    InMux I__1624 (
            .O(N__18480),
            .I(N__18448));
    Span4Mux_v I__1623 (
            .O(N__18471),
            .I(N__18445));
    Odrv4 I__1622 (
            .O(N__18466),
            .I(pwm_duty_input_10));
    LocalMux I__1621 (
            .O(N__18463),
            .I(pwm_duty_input_10));
    LocalMux I__1620 (
            .O(N__18448),
            .I(pwm_duty_input_10));
    Odrv4 I__1619 (
            .O(N__18445),
            .I(pwm_duty_input_10));
    CascadeMux I__1618 (
            .O(N__18436),
            .I(N__18433));
    InMux I__1617 (
            .O(N__18433),
            .I(N__18430));
    LocalMux I__1616 (
            .O(N__18430),
            .I(N__18427));
    Odrv4 I__1615 (
            .O(N__18427),
            .I(\current_shift_inst.PI_CTRL.m7_2 ));
    InMux I__1614 (
            .O(N__18424),
            .I(N__18419));
    InMux I__1613 (
            .O(N__18423),
            .I(N__18416));
    InMux I__1612 (
            .O(N__18422),
            .I(N__18413));
    LocalMux I__1611 (
            .O(N__18419),
            .I(N__18410));
    LocalMux I__1610 (
            .O(N__18416),
            .I(N__18407));
    LocalMux I__1609 (
            .O(N__18413),
            .I(pwm_duty_input_7));
    Odrv4 I__1608 (
            .O(N__18410),
            .I(pwm_duty_input_7));
    Odrv4 I__1607 (
            .O(N__18407),
            .I(pwm_duty_input_7));
    InMux I__1606 (
            .O(N__18400),
            .I(N__18397));
    LocalMux I__1605 (
            .O(N__18397),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__1604 (
            .O(N__18394),
            .I(N__18391));
    LocalMux I__1603 (
            .O(N__18391),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    CascadeMux I__1602 (
            .O(N__18388),
            .I(N__18385));
    InMux I__1601 (
            .O(N__18385),
            .I(N__18382));
    LocalMux I__1600 (
            .O(N__18382),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    CascadeMux I__1599 (
            .O(N__18379),
            .I(N__18376));
    InMux I__1598 (
            .O(N__18376),
            .I(N__18373));
    LocalMux I__1597 (
            .O(N__18373),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    InMux I__1596 (
            .O(N__18370),
            .I(N__18367));
    LocalMux I__1595 (
            .O(N__18367),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    InMux I__1594 (
            .O(N__18364),
            .I(N__18361));
    LocalMux I__1593 (
            .O(N__18361),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__1592 (
            .O(N__18358),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__1591 (
            .O(N__18355),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    InMux I__1590 (
            .O(N__18352),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__1589 (
            .O(N__18349),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    InMux I__1588 (
            .O(N__18346),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__1587 (
            .O(N__18343),
            .I(N__18340));
    LocalMux I__1586 (
            .O(N__18340),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__1585 (
            .O(N__18337),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__1584 (
            .O(N__18334),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    InMux I__1583 (
            .O(N__18331),
            .I(N__18327));
    InMux I__1582 (
            .O(N__18330),
            .I(N__18324));
    LocalMux I__1581 (
            .O(N__18327),
            .I(pwm_duty_input_2));
    LocalMux I__1580 (
            .O(N__18324),
            .I(pwm_duty_input_2));
    InMux I__1579 (
            .O(N__18319),
            .I(N__18314));
    InMux I__1578 (
            .O(N__18318),
            .I(N__18311));
    InMux I__1577 (
            .O(N__18317),
            .I(N__18308));
    LocalMux I__1576 (
            .O(N__18314),
            .I(N__18305));
    LocalMux I__1575 (
            .O(N__18311),
            .I(N__18302));
    LocalMux I__1574 (
            .O(N__18308),
            .I(N__18297));
    Span4Mux_s1_h I__1573 (
            .O(N__18305),
            .I(N__18297));
    Odrv4 I__1572 (
            .O(N__18302),
            .I(pwm_duty_input_3));
    Odrv4 I__1571 (
            .O(N__18297),
            .I(pwm_duty_input_3));
    CascadeMux I__1570 (
            .O(N__18292),
            .I(N__18289));
    InMux I__1569 (
            .O(N__18289),
            .I(N__18285));
    InMux I__1568 (
            .O(N__18288),
            .I(N__18282));
    LocalMux I__1567 (
            .O(N__18285),
            .I(pwm_duty_input_0));
    LocalMux I__1566 (
            .O(N__18282),
            .I(pwm_duty_input_0));
    InMux I__1565 (
            .O(N__18277),
            .I(N__18273));
    InMux I__1564 (
            .O(N__18276),
            .I(N__18270));
    LocalMux I__1563 (
            .O(N__18273),
            .I(N__18267));
    LocalMux I__1562 (
            .O(N__18270),
            .I(N__18264));
    Span4Mux_v I__1561 (
            .O(N__18267),
            .I(N__18261));
    Odrv4 I__1560 (
            .O(N__18264),
            .I(pwm_duty_input_1));
    Odrv4 I__1559 (
            .O(N__18261),
            .I(pwm_duty_input_1));
    InMux I__1558 (
            .O(N__18256),
            .I(N__18253));
    LocalMux I__1557 (
            .O(N__18253),
            .I(N__18250));
    Odrv12 I__1556 (
            .O(N__18250),
            .I(\current_shift_inst.PI_CTRL.m14_2 ));
    CascadeMux I__1555 (
            .O(N__18247),
            .I(\current_shift_inst.PI_CTRL.N_19_cascade_ ));
    InMux I__1554 (
            .O(N__18244),
            .I(N__18240));
    InMux I__1553 (
            .O(N__18243),
            .I(N__18236));
    LocalMux I__1552 (
            .O(N__18240),
            .I(N__18233));
    InMux I__1551 (
            .O(N__18239),
            .I(N__18230));
    LocalMux I__1550 (
            .O(N__18236),
            .I(pwm_duty_input_4));
    Odrv12 I__1549 (
            .O(N__18233),
            .I(pwm_duty_input_4));
    LocalMux I__1548 (
            .O(N__18230),
            .I(pwm_duty_input_4));
    InMux I__1547 (
            .O(N__18223),
            .I(N__18220));
    LocalMux I__1546 (
            .O(N__18220),
            .I(N__18217));
    Odrv4 I__1545 (
            .O(N__18217),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    InMux I__1544 (
            .O(N__18214),
            .I(N__18209));
    InMux I__1543 (
            .O(N__18213),
            .I(N__18204));
    InMux I__1542 (
            .O(N__18212),
            .I(N__18204));
    LocalMux I__1541 (
            .O(N__18209),
            .I(N__18199));
    LocalMux I__1540 (
            .O(N__18204),
            .I(N__18199));
    Odrv12 I__1539 (
            .O(N__18199),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    InMux I__1538 (
            .O(N__18196),
            .I(N__18193));
    LocalMux I__1537 (
            .O(N__18193),
            .I(N__18189));
    InMux I__1536 (
            .O(N__18192),
            .I(N__18186));
    Odrv4 I__1535 (
            .O(N__18189),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    LocalMux I__1534 (
            .O(N__18186),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    InMux I__1533 (
            .O(N__18181),
            .I(N__18178));
    LocalMux I__1532 (
            .O(N__18178),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    CascadeMux I__1531 (
            .O(N__18175),
            .I(N__18171));
    InMux I__1530 (
            .O(N__18174),
            .I(N__18167));
    InMux I__1529 (
            .O(N__18171),
            .I(N__18162));
    InMux I__1528 (
            .O(N__18170),
            .I(N__18162));
    LocalMux I__1527 (
            .O(N__18167),
            .I(N__18159));
    LocalMux I__1526 (
            .O(N__18162),
            .I(pwm_duty_input_9));
    Odrv4 I__1525 (
            .O(N__18159),
            .I(pwm_duty_input_9));
    InMux I__1524 (
            .O(N__18154),
            .I(N__18147));
    InMux I__1523 (
            .O(N__18153),
            .I(N__18147));
    InMux I__1522 (
            .O(N__18152),
            .I(N__18144));
    LocalMux I__1521 (
            .O(N__18147),
            .I(N__18141));
    LocalMux I__1520 (
            .O(N__18144),
            .I(N__18138));
    Odrv4 I__1519 (
            .O(N__18141),
            .I(pwm_duty_input_5));
    Odrv4 I__1518 (
            .O(N__18138),
            .I(pwm_duty_input_5));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_6 ),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_14 ),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_22 ),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_10_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_25_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_30 ),
            .carryinitout(bfn_10_25_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(un5_counter_cry_8),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_3_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_12_0_));
    defparam IN_MUX_bfv_3_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_13_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_3_13_0_));
    defparam IN_MUX_bfv_3_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_14_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_3_14_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_18_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_8_0_));
    defparam IN_MUX_bfv_18_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_9_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_18_9_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_12_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_24_0_));
    defparam IN_MUX_bfv_12_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_25_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_12_25_0_));
    defparam IN_MUX_bfv_12_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_26_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_12_26_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_8 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_16 ),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_24 ),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_3_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_10_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_3_10_0_));
    defparam IN_MUX_bfv_3_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_11_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_3_11_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_18_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_23_0_));
    defparam IN_MUX_bfv_18_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_24_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_18_24_0_));
    defparam IN_MUX_bfv_18_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_25_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_18_25_0_));
    defparam IN_MUX_bfv_18_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_26_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_18_26_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_17_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_24_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_17_24_0_));
    defparam IN_MUX_bfv_17_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_25_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_17_25_0_));
    defparam IN_MUX_bfv_17_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_26_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_17_26_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\current_shift_inst.z_cry_7 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\current_shift_inst.z_cry_15 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(\current_shift_inst.z_cry_23 ),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_8 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_16 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_24 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_16_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_25_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_16_25_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_7 ),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_15 ),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_23 ),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_7 ),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_15 ),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_23 ),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_4_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_17_0_));
    defparam IN_MUX_bfv_4_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_4_18_0_));
    defparam IN_MUX_bfv_4_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_4_19_0_));
    defparam IN_MUX_bfv_4_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_4_20_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryinitout(bfn_8_20_0_));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__27256),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_336_i_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__23056),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_187_i_g ));
    ICE_GB \current_shift_inst.timer_phase.running_RNIC90O_0  (
            .USERSIGNALTOGLOBALBUFFER(N__30070),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_phase.N_188_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__43350),
            .CLKHFEN(N__43449),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__43493),
            .RGB2PWM(N__19408),
            .RGB1(rgb_g),
            .CURREN(N__43334),
            .RGB2(rgb_b),
            .RGB1PWM(N__21415),
            .RGB0PWM(N__48279),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_5  (
            .in0(N__19081),
            .in1(N__18192),
            .in2(_gnd_net_),
            .in3(N__18487),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21528),
            .lcout(pwm_duty_input_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48874),
            .ce(N__25133),
            .sr(N__48174));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_1_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_1_8_3 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_1_8_3  (
            .in0(N__18318),
            .in1(N__18244),
            .in2(N__18175),
            .in3(N__18154),
            .lcout(\current_shift_inst.PI_CTRL.m7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_1_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_1_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_1_8_5  (
            .in0(N__18170),
            .in1(N__18424),
            .in2(N__18583),
            .in3(N__18153),
            .lcout(\current_shift_inst.PI_CTRL.m14_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_8_7 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_8_7  (
            .in0(N__18196),
            .in1(N__19077),
            .in2(N__18542),
            .in3(N__18181),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_9_2 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_9_2  (
            .in0(N__20917),
            .in1(N__19239),
            .in2(N__21527),
            .in3(N__19282),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48871),
            .ce(N__25081),
            .sr(N__48202));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_0 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_0  (
            .in0(N__19235),
            .in1(N__21514),
            .in2(N__20959),
            .in3(N__19277),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48868),
            .ce(N__25132),
            .sr(N__48209));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_1 .LUT_INIT=16'b1000111110001100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_1  (
            .in0(N__19274),
            .in1(N__20629),
            .in2(N__21526),
            .in3(N__19232),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48868),
            .ce(N__25132),
            .sr(N__48209));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_2 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_2  (
            .in0(N__19234),
            .in1(N__21513),
            .in2(N__20998),
            .in3(N__19276),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48868),
            .ce(N__25132),
            .sr(N__48209));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_4 .LUT_INIT=16'b1101110011011101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_4  (
            .in0(N__18982),
            .in1(N__20707),
            .in2(N__19240),
            .in3(N__19324),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48868),
            .ce(N__25132),
            .sr(N__48209));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_6 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_6  (
            .in0(N__19233),
            .in1(N__21512),
            .in2(N__21037),
            .in3(N__19275),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48868),
            .ce(N__25132),
            .sr(N__48209));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_7 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_7  (
            .in0(N__18214),
            .in1(N__18981),
            .in2(N__20764),
            .in3(N__19009),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48868),
            .ce(N__25132),
            .sr(N__48209));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_11_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_11_0  (
            .in0(N__18975),
            .in1(N__18213),
            .in2(N__20728),
            .in3(N__19005),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48864),
            .ce(N__25077),
            .sr(N__48213));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_11_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_11_4  (
            .in0(N__18974),
            .in1(N__18212),
            .in2(N__20782),
            .in3(N__19004),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48864),
            .ce(N__25077),
            .sr(N__48213));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_11_7 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_11_7  (
            .in0(N__20589),
            .in1(N__18223),
            .in2(N__20671),
            .in3(N__19281),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48864),
            .ce(N__25077),
            .sr(N__48213));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_1_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_1_12_1 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_1_12_1  (
            .in0(N__18331),
            .in1(N__18317),
            .in2(N__18292),
            .in3(N__18276),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_1_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_1_12_2 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_1_12_2  (
            .in0(N__18256),
            .in1(N__18541),
            .in2(N__18247),
            .in3(N__18243),
            .lcout(N_28_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_13_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_13_1  (
            .in0(N__19896),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19347),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_13_4 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_13_4  (
            .in0(N__20667),
            .in1(N__19303),
            .in2(N__21529),
            .in3(N__19216),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__20659),
            .in2(_gnd_net_),
            .in3(N__20699),
            .lcout(\current_shift_inst.PI_CTRL.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_15_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_15_4  (
            .in0(N__21505),
            .in1(N__19299),
            .in2(_gnd_net_),
            .in3(N__19203),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_2_7_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_2_7_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_2_7_4 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_2_7_4  (
            .in0(N__19610),
            .in1(N__19734),
            .in2(N__19671),
            .in3(N__18343),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48873),
            .ce(),
            .sr(N__48175));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_2_7_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_2_7_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_2_7_6 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_2_7_6  (
            .in0(N__19609),
            .in1(N__18364),
            .in2(N__19670),
            .in3(N__19735),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48873),
            .ce(),
            .sr(N__48175));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(N__19333),
            .in2(N__19858),
            .in3(N__19857),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__19789),
            .in2(_gnd_net_),
            .in3(N__18358),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__18394),
            .in2(_gnd_net_),
            .in3(N__18355),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_8_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18388),
            .in3(N__18352),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__18589),
            .in2(_gnd_net_),
            .in3(N__18349),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__18400),
            .in2(_gnd_net_),
            .in3(N__18346),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__18715),
            .in2(_gnd_net_),
            .in3(N__18337),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(N__18706),
            .in2(_gnd_net_),
            .in3(N__18334),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_9_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18697),
            .in3(N__18595),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_9_1 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_9_1  (
            .in0(N__20017),
            .in1(N__19853),
            .in2(N__20371),
            .in3(N__18592),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_2 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_2  (
            .in0(N__19851),
            .in1(N__20086),
            .in2(N__20194),
            .in3(N__20103),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_2_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_2_9_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_2_9_3  (
            .in0(N__18575),
            .in1(N__18543),
            .in2(N__18436),
            .in3(N__18422),
            .lcout(i8_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_4 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_4  (
            .in0(N__19852),
            .in1(N__20077),
            .in2(N__20167),
            .in3(N__20008),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_5 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_5  (
            .in0(N__20260),
            .in1(N__20317),
            .in2(N__19777),
            .in3(N__19850),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_6 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_6  (
            .in0(N__19849),
            .in1(N__19744),
            .in2(N__20227),
            .in3(N__19763),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_2_10_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_2_10_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_2_10_0 .LUT_INIT=16'b0101000000110000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_2_10_0  (
            .in0(N__19581),
            .in1(N__19659),
            .in2(N__18379),
            .in3(N__19704),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48865),
            .ce(),
            .sr(N__48203));
    defparam \pwm_generator_inst.threshold_9_LC_2_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_2_10_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_2_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18370),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48865),
            .ce(),
            .sr(N__48203));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_10_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_10_5  (
            .in0(N__19764),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20223),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_10_7  (
            .in0(N__20104),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20190),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_11_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_11_1  (
            .in0(N__20062),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20136),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_11_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_11_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_11_2  (
            .in0(N__20137),
            .in1(N__20050),
            .in2(N__18718),
            .in3(N__19845),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_11_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_11_4 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_11_4  (
            .in0(N__20119),
            .in1(N__19969),
            .in2(N__20041),
            .in3(N__19846),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_11_6 .LUT_INIT=16'b1011100001110100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_11_6  (
            .in0(N__19987),
            .in1(N__19847),
            .in2(N__20395),
            .in3(N__20029),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_12_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__18685),
            .in2(N__18670),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__18655),
            .in2(N__18646),
            .in3(N__18628),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__18625),
            .in2(N__18616),
            .in3(N__18598),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__18952),
            .in2(N__18943),
            .in3(N__18925),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__18922),
            .in2(N__18913),
            .in3(N__18895),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__18892),
            .in2(N__18877),
            .in3(N__18865),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__18862),
            .in2(N__18847),
            .in3(N__18835),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__18832),
            .in2(N__18817),
            .in3(N__18805),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__18802),
            .in2(N__18790),
            .in3(N__18772),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__18769),
            .in2(N__18760),
            .in3(N__18742),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__19056),
            .in2(N__18739),
            .in3(N__18721),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__19174),
            .in2(N__19074),
            .in3(N__19159),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__19060),
            .in2(N__19156),
            .in3(N__19138),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__19135),
            .in2(N__19075),
            .in3(N__19120),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__19064),
            .in2(N__19117),
            .in3(N__19099),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__19096),
            .in2(N__19076),
            .in3(N__19027),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_14_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_14_0  (
            .in0(N__20419),
            .in1(N__19024),
            .in2(_gnd_net_),
            .in3(N__19012),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_14_1 .LUT_INIT=16'b0000111100000010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_14_1  (
            .in0(N__19317),
            .in1(N__19217),
            .in2(N__20706),
            .in3(N__18965),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_14_2 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_14_2  (
            .in0(N__18988),
            .in1(N__21522),
            .in2(N__20593),
            .in3(N__19258),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_14_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_14_4 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_14_4  (
            .in0(N__19895),
            .in1(N__19351),
            .in2(N__19876),
            .in3(N__19810),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_14_6 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_14_6  (
            .in0(N__20660),
            .in1(N__21521),
            .in2(_gnd_net_),
            .in3(N__19298),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_2_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_2_15_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__20628),
            .in2(_gnd_net_),
            .in3(N__20994),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_15_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_15_4  (
            .in0(N__20952),
            .in1(N__21033),
            .in2(N__19306),
            .in3(N__20910),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_17_1  (
            .in0(N__20461),
            .in1(N__20512),
            .in2(N__20506),
            .in3(N__20488),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_2_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_2_17_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_2_17_3  (
            .in0(N__20407),
            .in1(N__20482),
            .in2(N__20473),
            .in3(N__19180),
            .lcout(\current_shift_inst.PI_CTRL.N_178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_2_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_2_18_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(N__20824),
            .in2(_gnd_net_),
            .in3(N__21169),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISHP8_10_LC_2_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISHP8_10_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISHP8_10_LC_2_18_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISHP8_10_LC_2_18_5  (
            .in0(N__20413),
            .in1(N__20854),
            .in2(N__19183),
            .in3(N__20874),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_2_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_2_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_2_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28105),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48801),
            .ce(N__25152),
            .sr(N__48238));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_2_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_2_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_2_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28762),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48801),
            .ce(N__25152),
            .sr(N__48238));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_2_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_2_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_2_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_2_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28684),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48801),
            .ce(N__25152),
            .sr(N__48238));
    defparam \current_shift_inst.N_22_i_i_LC_2_28_4 .C_ON=1'b0;
    defparam \current_shift_inst.N_22_i_i_LC_2_28_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.N_22_i_i_LC_2_28_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.N_22_i_i_LC_2_28_4  (
            .in0(N__48278),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31032),
            .lcout(N_22_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_7_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_7_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_7_0 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_3_7_0  (
            .in0(N__19732),
            .in1(N__19608),
            .in2(N__19672),
            .in3(N__19396),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48872),
            .ce(),
            .sr(N__48163));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_7_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_7_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_7_1 .LUT_INIT=16'b0100000001110000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_3_7_1  (
            .in0(N__19607),
            .in1(N__19733),
            .in2(N__19390),
            .in3(N__19669),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48872),
            .ce(),
            .sr(N__48163));
    defparam \pwm_generator_inst.threshold_6_LC_3_7_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_3_7_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_3_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_3_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19381),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48872),
            .ce(),
            .sr(N__48163));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_8_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_3_8_1 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_3_8_1  (
            .in0(N__19728),
            .in1(N__19657),
            .in2(N__19614),
            .in3(N__19375),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48869),
            .ce(),
            .sr(N__48176));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_8_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_8_2 .LUT_INIT=16'b0001110100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_3_8_2  (
            .in0(N__19654),
            .in1(N__19730),
            .in2(N__19611),
            .in3(N__19369),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48869),
            .ce(),
            .sr(N__48176));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_8_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_8_5 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_3_8_5  (
            .in0(N__19727),
            .in1(N__19656),
            .in2(N__19613),
            .in3(N__19363),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48869),
            .ce(),
            .sr(N__48176));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_8_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_8_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_8_6 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_3_8_6  (
            .in0(N__19655),
            .in1(N__19731),
            .in2(N__19612),
            .in3(N__19357),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48869),
            .ce(),
            .sr(N__48176));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_8_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_8_7 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_3_8_7  (
            .in0(N__19729),
            .in1(N__19658),
            .in2(N__19615),
            .in3(N__19540),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48869),
            .ce(),
            .sr(N__48176));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(N__19522),
            .in2(_gnd_net_),
            .in3(N__19534),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1  (
            .in0(_gnd_net_),
            .in1(N__19504),
            .in2(_gnd_net_),
            .in3(N__19516),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(N__19486),
            .in2(_gnd_net_),
            .in3(N__19498),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3  (
            .in0(_gnd_net_),
            .in1(N__19468),
            .in2(_gnd_net_),
            .in3(N__19480),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4  (
            .in0(_gnd_net_),
            .in1(N__19450),
            .in2(_gnd_net_),
            .in3(N__19462),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5  (
            .in0(_gnd_net_),
            .in1(N__19432),
            .in2(_gnd_net_),
            .in3(N__19444),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(N__19414),
            .in2(_gnd_net_),
            .in3(N__19426),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7  (
            .in0(_gnd_net_),
            .in1(N__19942),
            .in2(_gnd_net_),
            .in3(N__19954),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(N__19924),
            .in2(_gnd_net_),
            .in3(N__19936),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_3_10_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1  (
            .in0(_gnd_net_),
            .in1(N__19906),
            .in2(_gnd_net_),
            .in3(N__19918),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(N__19900),
            .in2(_gnd_net_),
            .in3(N__19861),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3  (
            .in0(N__19848),
            .in1(N__20293),
            .in2(_gnd_net_),
            .in3(N__19780),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20316),
            .in3(N__19768),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19765),
            .in3(N__19738),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6  (
            .in0(_gnd_net_),
            .in1(N__20102),
            .in2(_gnd_net_),
            .in3(N__20080),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7  (
            .in0(_gnd_net_),
            .in1(N__20003),
            .in2(_gnd_net_),
            .in3(N__20065),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0  (
            .in0(_gnd_net_),
            .in1(N__20061),
            .in2(_gnd_net_),
            .in3(N__20044),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_3_11_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1  (
            .in0(_gnd_net_),
            .in1(N__19967),
            .in2(_gnd_net_),
            .in3(N__20032),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__19985),
            .in2(_gnd_net_),
            .in3(N__20023),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20020),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_3_11_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_3_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_3_11_4  (
            .in0(N__20007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20160),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_3_11_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_3_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_3_11_5  (
            .in0(N__19986),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20391),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_3_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_3_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_3_11_6  (
            .in0(N__19968),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20118),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_3_11_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_3_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_3_11_7  (
            .in0(N__20315),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20256),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_3_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_3_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(N__20292),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_12_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_3_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_3_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_3_12_1  (
            .in0(_gnd_net_),
            .in1(N__20272),
            .in2(_gnd_net_),
            .in3(N__20245),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_3_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_3_12_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20242),
            .in3(N__20209),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_3_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_3_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_3_12_3  (
            .in0(_gnd_net_),
            .in1(N__20206),
            .in2(_gnd_net_),
            .in3(N__20176),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_3_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_3_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_3_12_4  (
            .in0(_gnd_net_),
            .in1(N__20173),
            .in2(_gnd_net_),
            .in3(N__20149),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_3_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_3_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_3_12_5  (
            .in0(_gnd_net_),
            .in1(N__43430),
            .in2(N__20146),
            .in3(N__20128),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_3_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_3_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_3_12_6  (
            .in0(_gnd_net_),
            .in1(N__20125),
            .in2(N__43472),
            .in3(N__20107),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_3_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_3_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_3_12_7  (
            .in0(_gnd_net_),
            .in1(N__20401),
            .in2(N__43434),
            .in3(N__20380),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_3_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_3_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(N__20377),
            .in2(_gnd_net_),
            .in3(N__20356),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_3_13_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_3_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_3_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(N__20353),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_3_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_3_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(N__20347),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_3_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_3_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_3_13_3  (
            .in0(_gnd_net_),
            .in1(N__20341),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_3_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_3_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_3_13_4  (
            .in0(_gnd_net_),
            .in1(N__20335),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_3_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_3_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_3_13_5  (
            .in0(_gnd_net_),
            .in1(N__20329),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_3_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_3_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_3_13_6  (
            .in0(_gnd_net_),
            .in1(N__20323),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_3_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_3_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_3_13_7  (
            .in0(_gnd_net_),
            .in1(N__20452),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_3_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_3_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_3_14_0  (
            .in0(_gnd_net_),
            .in1(N__20446),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_14_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_3_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_3_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(N__20440),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_3_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_3_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(N__20434),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_3_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_3_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__20428),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_3_14_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_3_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20422),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIEE4_12_LC_3_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIEE4_12_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIEE4_12_LC_3_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIEE4_12_LC_3_17_0  (
            .in0(N__21247),
            .in1(N__20806),
            .in2(N__21229),
            .in3(N__20836),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_3_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_3_17_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_3_17_3  (
            .in0(N__26376),
            .in1(N__26338),
            .in2(N__26301),
            .in3(N__26257),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRMD4_17_LC_3_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRMD4_17_LC_3_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRMD4_17_LC_3_17_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRMD4_17_LC_3_17_5  (
            .in0(N__21337),
            .in1(N__21115),
            .in2(N__21136),
            .in3(N__21298),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMJ62_12_LC_3_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMJ62_12_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMJ62_12_LC_3_17_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMJ62_12_LC_3_17_6  (
            .in0(N__21355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20835),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU8H5_14_LC_3_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU8H5_14_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU8H5_14_LC_3_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIU8H5_14_LC_3_17_7  (
            .in0(N__20805),
            .in1(N__21297),
            .in2(N__20515),
            .in3(N__21336),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_10_LC_3_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_10_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_10_LC_3_18_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_10_LC_3_18_1  (
            .in0(N__21246),
            .in1(N__20850),
            .in2(N__20875),
            .in3(N__21225),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_3_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_3_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_3_18_2  (
            .in0(N__21129),
            .in1(N__21162),
            .in2(N__21114),
            .in3(N__21183),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPM62_13_LC_3_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPM62_13_LC_3_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPM62_13_LC_3_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPM62_13_LC_3_18_3  (
            .in0(_gnd_net_),
            .in1(N__21316),
            .in2(_gnd_net_),
            .in3(N__20820),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKAQ8_27_LC_3_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKAQ8_27_LC_3_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKAQ8_27_LC_3_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIKAQ8_27_LC_3_18_4  (
            .in0(N__21265),
            .in1(N__21283),
            .in2(N__20497),
            .in3(N__20494),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI9LI5_19_LC_3_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI9LI5_19_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI9LI5_19_LC_3_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI9LI5_19_LC_3_19_0  (
            .in0(N__21094),
            .in1(N__20554),
            .in2(N__21082),
            .in3(N__21315),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIEAE4_15_LC_3_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIEAE4_15_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIEAE4_15_LC_3_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIEAE4_15_LC_3_19_2  (
            .in0(N__21067),
            .in1(N__21354),
            .in2(N__21187),
            .in3(N__21051),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_3_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_3_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_3_19_3  (
            .in0(N__21066),
            .in1(N__21078),
            .in2(N__21052),
            .in3(N__21093),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1082_27_LC_3_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1082_27_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1082_27_LC_3_20_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1082_27_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__21261),
            .in2(_gnd_net_),
            .in3(N__21279),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_0.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_0.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20548),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNII76D_3_LC_4_7_7.C_ON=1'b0;
    defparam counter_RNII76D_3_LC_4_7_7.SEQ_MODE=4'b0000;
    defparam counter_RNII76D_3_LC_4_7_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 counter_RNII76D_3_LC_4_7_7 (
            .in0(N__21369),
            .in1(N__21384),
            .in2(N__21658),
            .in3(N__21399),
            .lcout(un2_counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_7_LC_4_8_0.C_ON=1'b0;
    defparam counter_7_LC_4_8_0.SEQ_MODE=4'b1010;
    defparam counter_7_LC_4_8_0.LUT_INIT=16'b0111000011110000;
    LogicCell40 counter_7_LC_4_8_0 (
            .in0(N__21721),
            .in1(N__21751),
            .in2(N__21640),
            .in3(N__21786),
            .lcout(counterZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48866),
            .ce(),
            .sr(N__48164));
    defparam counter_12_LC_4_8_5.C_ON=1'b0;
    defparam counter_12_LC_4_8_5.SEQ_MODE=4'b1010;
    defparam counter_12_LC_4_8_5.LUT_INIT=16'b0111000011110000;
    LogicCell40 counter_12_LC_4_8_5 (
            .in0(N__21750),
            .in1(N__21785),
            .in2(N__21604),
            .in3(N__21720),
            .lcout(counterZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48866),
            .ce(),
            .sr(N__48164));
    defparam counter_1_LC_4_9_2.C_ON=1'b0;
    defparam counter_1_LC_4_9_2.SEQ_MODE=4'b1010;
    defparam counter_1_LC_4_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_1_LC_4_9_2 (
            .in0(_gnd_net_),
            .in1(N__21552),
            .in2(_gnd_net_),
            .in3(N__21872),
            .lcout(counterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48860),
            .ce(),
            .sr(N__48177));
    defparam \pwm_generator_inst.threshold_8_LC_4_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_4_9_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_4_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20521),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48860),
            .ce(),
            .sr(N__48177));
    defparam counter_10_LC_4_9_6.C_ON=1'b0;
    defparam counter_10_LC_4_9_6.SEQ_MODE=4'b1010;
    defparam counter_10_LC_4_9_6.LUT_INIT=16'b0111000011110000;
    LogicCell40 counter_10_LC_4_9_6 (
            .in0(N__21719),
            .in1(N__21749),
            .in2(N__21622),
            .in3(N__21792),
            .lcout(counterZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48860),
            .ce(),
            .sr(N__48177));
    defparam counter_0_LC_4_9_7.C_ON=1'b0;
    defparam counter_0_LC_4_9_7.SEQ_MODE=4'b1010;
    defparam counter_0_LC_4_9_7.LUT_INIT=16'b0000011100001111;
    LogicCell40 counter_0_LC_4_9_7 (
            .in0(N__21748),
            .in1(N__21791),
            .in2(N__21874),
            .in3(N__21718),
            .lcout(counterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48860),
            .ce(),
            .sr(N__48177));
    defparam clk_10khz_RNIIENA2_LC_4_10_1.C_ON=1'b0;
    defparam clk_10khz_RNIIENA2_LC_4_10_1.SEQ_MODE=4'b0000;
    defparam clk_10khz_RNIIENA2_LC_4_10_1.LUT_INIT=16'b0111100011110000;
    LogicCell40 clk_10khz_RNIIENA2_LC_4_10_1 (
            .in0(N__21746),
            .in1(N__21790),
            .in2(N__21689),
            .in3(N__21716),
            .lcout(clk_10khz_RNIIENAZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_4_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_4_11_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_4_11_1  (
            .in0(N__30988),
            .in1(N__21682),
            .in2(_gnd_net_),
            .in3(N__20565),
            .lcout(N_717_g),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU1LD_7_LC_4_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU1LD_7_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU1LD_7_LC_4_11_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIU1LD_7_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(N__20903),
            .in2(_gnd_net_),
            .in3(N__20990),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_4_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_4_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_4_11_5  (
            .in0(N__20945),
            .in1(N__21029),
            .in2(N__20596),
            .in3(N__20624),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_4_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_4_12_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \current_shift_inst.phase_valid_RNISLOR2_LC_4_12_7  (
            .in0(N__21690),
            .in1(N__24277),
            .in2(N__31033),
            .in3(N__20569),
            .lcout(\current_shift_inst.phase_valid_RNISLORZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_4_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_4_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_4_14_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_4_14_0  (
            .in0(N__23368),
            .in1(N__23492),
            .in2(N__23632),
            .in3(N__22507),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48829),
            .ce(),
            .sr(N__48214));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_4_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_4_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_4_14_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_4_14_2  (
            .in0(N__23365),
            .in1(N__23483),
            .in2(N__23629),
            .in3(N__22753),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48829),
            .ce(),
            .sr(N__48214));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_4_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_4_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_4_14_3 .LUT_INIT=16'b1010100010001010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_4_14_3  (
            .in0(N__22726),
            .in1(N__23493),
            .in2(N__23391),
            .in3(N__23613),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48829),
            .ce(),
            .sr(N__48214));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_4_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_4_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_4_14_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_4_14_4  (
            .in0(N__23366),
            .in1(N__23484),
            .in2(N__23630),
            .in3(N__22699),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48829),
            .ce(),
            .sr(N__48214));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_4_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_4_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_4_14_5 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_4_14_5  (
            .in0(N__23369),
            .in1(N__23617),
            .in2(N__23502),
            .in3(N__22669),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48829),
            .ce(),
            .sr(N__48214));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_4_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_4_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_4_14_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_4_14_6  (
            .in0(N__23367),
            .in1(N__23488),
            .in2(N__23631),
            .in3(N__22642),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48829),
            .ce(),
            .sr(N__48214));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_4_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_4_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_4_14_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_4_14_7  (
            .in0(N__23370),
            .in1(N__23621),
            .in2(N__23503),
            .in3(N__22612),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48829),
            .ce(),
            .sr(N__48214));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28183),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48819),
            .ce(N__25054),
            .sr(N__48218));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_17_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_17_0  (
            .in0(_gnd_net_),
            .in1(N__23938),
            .in2(N__20797),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__48802),
            .ce(N__25106),
            .sr(N__48225));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_17_1  (
            .in0(_gnd_net_),
            .in1(N__23914),
            .in2(N__22138),
            .in3(N__20746),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__48802),
            .ce(N__25106),
            .sr(N__48225));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_17_2  (
            .in0(_gnd_net_),
            .in1(N__23889),
            .in2(N__20743),
            .in3(N__20710),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__48802),
            .ce(N__25106),
            .sr(N__48225));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_17_3  (
            .in0(_gnd_net_),
            .in1(N__23845),
            .in2(N__22123),
            .in3(N__20674),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__48802),
            .ce(N__25106),
            .sr(N__48225));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(N__22144),
            .in2(N__23818),
            .in3(N__20632),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__48802),
            .ce(N__25106),
            .sr(N__48225));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_17_5  (
            .in0(_gnd_net_),
            .in1(N__23769),
            .in2(N__22081),
            .in3(N__20599),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__48802),
            .ce(N__25106),
            .sr(N__48225));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_17_6  (
            .in0(_gnd_net_),
            .in1(N__23731),
            .in2(N__23002),
            .in3(N__21001),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__48802),
            .ce(N__25106),
            .sr(N__48225));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_17_7  (
            .in0(_gnd_net_),
            .in1(N__23695),
            .in2(N__22153),
            .in3(N__20962),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__48802),
            .ce(N__25106),
            .sr(N__48225));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__24079),
            .in2(N__22969),
            .in3(N__20920),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_4_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__48792),
            .ce(N__25154),
            .sr(N__48230));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_18_1  (
            .in0(_gnd_net_),
            .in1(N__24034),
            .in2(N__22114),
            .in3(N__20878),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__48792),
            .ce(N__25154),
            .sr(N__48230));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_18_2  (
            .in0(_gnd_net_),
            .in1(N__26256),
            .in2(N__22252),
            .in3(N__20857),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__48792),
            .ce(N__25154),
            .sr(N__48230));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(N__26574),
            .in2(N__22225),
            .in3(N__20839),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__48792),
            .ce(N__25154),
            .sr(N__48230));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(N__26784),
            .in2(N__22939),
            .in3(N__20827),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__48792),
            .ce(N__25154),
            .sr(N__48230));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_18_5  (
            .in0(_gnd_net_),
            .in1(N__26653),
            .in2(N__21439),
            .in3(N__20809),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__48792),
            .ce(N__25154),
            .sr(N__48230));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_18_6  (
            .in0(_gnd_net_),
            .in1(N__22129),
            .in2(N__26695),
            .in3(N__21205),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__48792),
            .ce(N__25154),
            .sr(N__48230));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_18_7  (
            .in0(_gnd_net_),
            .in1(N__26337),
            .in2(N__21202),
            .in3(N__21172),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__48792),
            .ce(N__25154),
            .sr(N__48230));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_19_0  (
            .in0(_gnd_net_),
            .in1(N__26612),
            .in2(N__22270),
            .in3(N__21151),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_4_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__48784),
            .ce(N__25064),
            .sr(N__48233));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_19_1  (
            .in0(_gnd_net_),
            .in1(N__24826),
            .in2(N__21148),
            .in3(N__21118),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__48784),
            .ce(N__25064),
            .sr(N__48233));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_19_2  (
            .in0(_gnd_net_),
            .in1(N__24184),
            .in2(N__21427),
            .in3(N__21097),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__48784),
            .ce(N__25064),
            .sr(N__48233));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_19_3  (
            .in0(_gnd_net_),
            .in1(N__24937),
            .in2(N__22261),
            .in3(N__21085),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__48784),
            .ce(N__25064),
            .sr(N__48233));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(N__24972),
            .in2(N__22984),
            .in3(N__21070),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__48784),
            .ce(N__25064),
            .sr(N__48233));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_19_5  (
            .in0(_gnd_net_),
            .in1(N__26407),
            .in2(N__22243),
            .in3(N__21055),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__48784),
            .ce(N__25064),
            .sr(N__48233));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(N__24883),
            .in2(N__22234),
            .in3(N__21040),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__48784),
            .ce(N__25064),
            .sr(N__48233));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_19_7  (
            .in0(_gnd_net_),
            .in1(N__26375),
            .in2(N__22213),
            .in3(N__21340),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__48784),
            .ce(N__25064),
            .sr(N__48233));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_20_0  (
            .in0(_gnd_net_),
            .in1(N__26490),
            .in2(N__22954),
            .in3(N__21319),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_4_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__48775),
            .ce(N__25155),
            .sr(N__48236));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(N__26530),
            .in2(N__22199),
            .in3(N__21301),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__48775),
            .ce(N__25155),
            .sr(N__48236));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_20_2  (
            .in0(_gnd_net_),
            .in1(N__22189),
            .in2(N__26455),
            .in3(N__21286),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__48775),
            .ce(N__25155),
            .sr(N__48236));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_20_3  (
            .in0(_gnd_net_),
            .in1(N__26819),
            .in2(N__22200),
            .in3(N__21268),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__48775),
            .ce(N__25155),
            .sr(N__48236));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(N__22193),
            .in2(N__26749),
            .in3(N__21250),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__48775),
            .ce(N__25155),
            .sr(N__48236));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_20_5  (
            .in0(_gnd_net_),
            .in1(N__26294),
            .in2(N__22201),
            .in3(N__21232),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__48775),
            .ce(N__25155),
            .sr(N__48236));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_20_6  (
            .in0(_gnd_net_),
            .in1(N__22197),
            .in2(N__26191),
            .in3(N__21208),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__48775),
            .ce(N__25155),
            .sr(N__48236));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_20_7  (
            .in0(N__22198),
            .in1(N__25520),
            .in2(_gnd_net_),
            .in3(N__21532),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48775),
            .ce(N__25155),
            .sr(N__48236));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_4_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28212),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48766),
            .ce(N__25172),
            .sr(N__48239));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_4_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_4_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_4_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_4_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28647),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48757),
            .ce(N__25153),
            .sr(N__48241));
    defparam \current_shift_inst.un7_start_stop_0_a3_LC_4_28_4 .C_ON=1'b0;
    defparam \current_shift_inst.un7_start_stop_0_a3_LC_4_28_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un7_start_stop_0_a3_LC_4_28_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \current_shift_inst.un7_start_stop_0_a3_LC_4_28_4  (
            .in0(N__48277),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31028),
            .lcout(un7_start_stop_0_a3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_counter_cry_1_c_LC_5_7_0.C_ON=1'b1;
    defparam un5_counter_cry_1_c_LC_5_7_0.SEQ_MODE=4'b0000;
    defparam un5_counter_cry_1_c_LC_5_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_counter_cry_1_c_LC_5_7_0 (
            .in0(_gnd_net_),
            .in1(N__21873),
            .in2(N__21556),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(un5_counter_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_2_LC_5_7_1.C_ON=1'b1;
    defparam counter_2_LC_5_7_1.SEQ_MODE=4'b1010;
    defparam counter_2_LC_5_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_2_LC_5_7_1 (
            .in0(_gnd_net_),
            .in1(N__21570),
            .in2(_gnd_net_),
            .in3(N__21403),
            .lcout(counterZ0Z_2),
            .ltout(),
            .carryin(un5_counter_cry_1),
            .carryout(un5_counter_cry_2),
            .clk(N__48867),
            .ce(),
            .sr(N__48149));
    defparam counter_3_LC_5_7_2.C_ON=1'b1;
    defparam counter_3_LC_5_7_2.SEQ_MODE=4'b1010;
    defparam counter_3_LC_5_7_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_3_LC_5_7_2 (
            .in0(_gnd_net_),
            .in1(N__21400),
            .in2(_gnd_net_),
            .in3(N__21388),
            .lcout(counterZ0Z_3),
            .ltout(),
            .carryin(un5_counter_cry_2),
            .carryout(un5_counter_cry_3),
            .clk(N__48867),
            .ce(),
            .sr(N__48149));
    defparam counter_4_LC_5_7_3.C_ON=1'b1;
    defparam counter_4_LC_5_7_3.SEQ_MODE=4'b1010;
    defparam counter_4_LC_5_7_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_4_LC_5_7_3 (
            .in0(_gnd_net_),
            .in1(N__21385),
            .in2(_gnd_net_),
            .in3(N__21373),
            .lcout(counterZ0Z_4),
            .ltout(),
            .carryin(un5_counter_cry_3),
            .carryout(un5_counter_cry_4),
            .clk(N__48867),
            .ce(),
            .sr(N__48149));
    defparam counter_5_LC_5_7_4.C_ON=1'b1;
    defparam counter_5_LC_5_7_4.SEQ_MODE=4'b1010;
    defparam counter_5_LC_5_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_5_LC_5_7_4 (
            .in0(_gnd_net_),
            .in1(N__21370),
            .in2(_gnd_net_),
            .in3(N__21358),
            .lcout(counterZ0Z_5),
            .ltout(),
            .carryin(un5_counter_cry_4),
            .carryout(un5_counter_cry_5),
            .clk(N__48867),
            .ce(),
            .sr(N__48149));
    defparam counter_6_LC_5_7_5.C_ON=1'b1;
    defparam counter_6_LC_5_7_5.SEQ_MODE=4'b1010;
    defparam counter_6_LC_5_7_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_6_LC_5_7_5 (
            .in0(_gnd_net_),
            .in1(N__21657),
            .in2(_gnd_net_),
            .in3(N__21643),
            .lcout(counterZ0Z_6),
            .ltout(),
            .carryin(un5_counter_cry_5),
            .carryout(un5_counter_cry_6),
            .clk(N__48867),
            .ce(),
            .sr(N__48149));
    defparam counter_RNO_0_7_LC_5_7_6.C_ON=1'b1;
    defparam counter_RNO_0_7_LC_5_7_6.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_7_LC_5_7_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_7_LC_5_7_6 (
            .in0(_gnd_net_),
            .in1(N__21583),
            .in2(_gnd_net_),
            .in3(N__21631),
            .lcout(counter_RNO_0Z0Z_7),
            .ltout(),
            .carryin(un5_counter_cry_6),
            .carryout(un5_counter_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_8_LC_5_7_7.C_ON=1'b1;
    defparam counter_8_LC_5_7_7.SEQ_MODE=4'b1010;
    defparam counter_8_LC_5_7_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_8_LC_5_7_7 (
            .in0(_gnd_net_),
            .in1(N__21807),
            .in2(_gnd_net_),
            .in3(N__21628),
            .lcout(counterZ0Z_8),
            .ltout(),
            .carryin(un5_counter_cry_7),
            .carryout(un5_counter_cry_8),
            .clk(N__48867),
            .ce(),
            .sr(N__48149));
    defparam counter_9_LC_5_8_0.C_ON=1'b1;
    defparam counter_9_LC_5_8_0.SEQ_MODE=4'b1010;
    defparam counter_9_LC_5_8_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_9_LC_5_8_0 (
            .in0(_gnd_net_),
            .in1(N__21835),
            .in2(_gnd_net_),
            .in3(N__21625),
            .lcout(counterZ0Z_9),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(un5_counter_cry_9),
            .clk(N__48861),
            .ce(),
            .sr(N__48155));
    defparam counter_RNO_0_10_LC_5_8_1.C_ON=1'b1;
    defparam counter_RNO_0_10_LC_5_8_1.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_10_LC_5_8_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_10_LC_5_8_1 (
            .in0(_gnd_net_),
            .in1(N__21595),
            .in2(_gnd_net_),
            .in3(N__21613),
            .lcout(counter_RNO_0Z0Z_10),
            .ltout(),
            .carryin(un5_counter_cry_9),
            .carryout(un5_counter_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_11_LC_5_8_2.C_ON=1'b1;
    defparam counter_11_LC_5_8_2.SEQ_MODE=4'b1010;
    defparam counter_11_LC_5_8_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_11_LC_5_8_2 (
            .in0(_gnd_net_),
            .in1(N__21847),
            .in2(_gnd_net_),
            .in3(N__21610),
            .lcout(counterZ0Z_11),
            .ltout(),
            .carryin(un5_counter_cry_10),
            .carryout(un5_counter_cry_11),
            .clk(N__48861),
            .ce(),
            .sr(N__48155));
    defparam counter_RNO_0_12_LC_5_8_3.C_ON=1'b0;
    defparam counter_RNO_0_12_LC_5_8_3.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_12_LC_5_8_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 counter_RNO_0_12_LC_5_8_3 (
            .in0(_gnd_net_),
            .in1(N__21822),
            .in2(_gnd_net_),
            .in3(N__21607),
            .lcout(counter_RNO_0Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI800G_7_LC_5_9_1.C_ON=1'b0;
    defparam counter_RNI800G_7_LC_5_9_1.SEQ_MODE=4'b0000;
    defparam counter_RNI800G_7_LC_5_9_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 counter_RNI800G_7_LC_5_9_1 (
            .in0(_gnd_net_),
            .in1(N__21594),
            .in2(_gnd_net_),
            .in3(N__21582),
            .lcout(),
            .ltout(un2_counter_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI3BSP_1_LC_5_9_2.C_ON=1'b0;
    defparam counter_RNI3BSP_1_LC_5_9_2.SEQ_MODE=4'b0000;
    defparam counter_RNI3BSP_1_LC_5_9_2.LUT_INIT=16'b0000000000010000;
    LogicCell40 counter_RNI3BSP_1_LC_5_9_2 (
            .in0(N__21571),
            .in1(N__21548),
            .in2(N__21877),
            .in3(N__21865),
            .lcout(un2_counter_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIM6001_12_LC_5_9_4.C_ON=1'b0;
    defparam counter_RNIM6001_12_LC_5_9_4.SEQ_MODE=4'b0000;
    defparam counter_RNIM6001_12_LC_5_9_4.LUT_INIT=16'b0000000000010000;
    LogicCell40 counter_RNIM6001_12_LC_5_9_4 (
            .in0(N__21846),
            .in1(N__21834),
            .in2(N__21823),
            .in3(N__21808),
            .lcout(un2_counter_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_10khz_LC_5_10_6.C_ON=1'b0;
    defparam clk_10khz_LC_5_10_6.SEQ_MODE=4'b1010;
    defparam clk_10khz_LC_5_10_6.LUT_INIT=16'b0111100011110000;
    LogicCell40 clk_10khz_LC_5_10_6 (
            .in0(N__21793),
            .in1(N__21747),
            .in2(N__21691),
            .in3(N__21717),
            .lcout(clk_10khz_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48848),
            .ce(),
            .sr(N__48178));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_5_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_5_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_5_11_0 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_5_11_0  (
            .in0(N__35774),
            .in1(N__35713),
            .in2(N__36450),
            .in3(N__36655),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48842),
            .ce(N__24637),
            .sr(N__48187));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_5_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_5_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_5_11_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_5_11_1  (
            .in0(N__36658),
            .in1(N__36439),
            .in2(N__35266),
            .in3(N__35777),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48842),
            .ce(N__24637),
            .sr(N__48187));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_5_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_5_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_5_11_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_5_11_3  (
            .in0(N__36660),
            .in1(N__36441),
            .in2(_gnd_net_),
            .in3(N__36496),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48842),
            .ce(N__24637),
            .sr(N__48187));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_5_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_5_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_5_11_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_5_11_4  (
            .in0(N__36440),
            .in1(N__36150),
            .in2(_gnd_net_),
            .in3(N__36659),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48842),
            .ce(N__24637),
            .sr(N__48187));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_5_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_5_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_5_11_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_5_11_5  (
            .in0(N__36656),
            .in1(N__35775),
            .in2(N__35380),
            .in3(N__36437),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48842),
            .ce(N__24637),
            .sr(N__48187));
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_5_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_5_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_5_11_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_0_LC_5_11_6  (
            .in0(N__35773),
            .in1(N__35841),
            .in2(N__36449),
            .in3(N__36654),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48842),
            .ce(N__24637),
            .sr(N__48187));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_5_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_5_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_5_11_7 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_5_11_7  (
            .in0(N__36657),
            .in1(N__35776),
            .in2(N__36094),
            .in3(N__36438),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48842),
            .ce(N__24637),
            .sr(N__48187));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_5_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_5_12_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_5_12_0  (
            .in0(N__23375),
            .in1(N__23498),
            .in2(N__23625),
            .in3(N__22576),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48838),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_5_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_5_12_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_5_12_1  (
            .in0(N__23494),
            .in1(N__23597),
            .in2(N__23392),
            .in3(N__22858),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48838),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_5_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_5_12_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_5_12_2  (
            .in0(N__23376),
            .in1(N__23499),
            .in2(N__23626),
            .in3(N__22822),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48838),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_5_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_5_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_5_12_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_5_12_3  (
            .in0(N__23495),
            .in1(N__23604),
            .in2(N__23393),
            .in3(N__22543),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48838),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_5_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_5_12_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_5_12_4  (
            .in0(N__23377),
            .in1(N__23500),
            .in2(N__23627),
            .in3(N__22090),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48838),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_5_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_5_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_5_12_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_5_12_5  (
            .in0(N__23496),
            .in1(N__23605),
            .in2(N__23394),
            .in3(N__22474),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48838),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_5_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_5_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_5_12_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_5_12_6  (
            .in0(N__23378),
            .in1(N__23501),
            .in2(N__23628),
            .in3(N__22441),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48838),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_5_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_5_12_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_5_12_7  (
            .in0(N__23497),
            .in1(N__23609),
            .in2(N__23395),
            .in3(N__22408),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48838),
            .ce(),
            .sr(N__48195));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_5_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_5_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__21886),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_5_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_5_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__22000),
            .in2(N__22012),
            .in3(N__22286),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_5_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_5_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__21982),
            .in2(N__21994),
            .in3(N__22554),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_5_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_5_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__21964),
            .in2(N__21976),
            .in3(N__22518),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_5_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_5_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__21946),
            .in2(N__21958),
            .in3(N__22485),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_5_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_5_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__21925),
            .in2(N__21940),
            .in3(N__22452),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_5_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_5_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__21919),
            .in2(N__24679),
            .in3(N__22419),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_5_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_5_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(N__21913),
            .in2(N__24667),
            .in3(N__23254),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_5_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_5_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__21892),
            .in2(N__21907),
            .in3(N__23230),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_5_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_5_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__22069),
            .in2(N__22363),
            .in3(N__23203),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_5_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_5_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__22063),
            .in2(N__23104),
            .in3(N__22764),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_5_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_5_14_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_5_14_3  (
            .in0(N__22737),
            .in1(N__22057),
            .in2(N__22348),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_5_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_5_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__22051),
            .in2(N__24652),
            .in3(N__22710),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_5_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_5_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__22045),
            .in2(N__23089),
            .in3(N__22686),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_5_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_5_14_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_5_14_6  (
            .in0(N__22653),
            .in1(N__22039),
            .in2(N__23119),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_5_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_5_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_5_14_7  (
            .in0(N__22623),
            .in1(N__23149),
            .in2(N__22033),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_5_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_5_15_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_5_15_0  (
            .in0(N__23647),
            .in1(N__22024),
            .in2(N__23071),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_5_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_5_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__22018),
            .in2(N__22330),
            .in3(N__22593),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_5_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_5_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__22105),
            .in2(N__22315),
            .in3(N__22875),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_5_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_5_15_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_5_15_3  (
            .in0(N__22839),
            .in1(N__22099),
            .in2(N__23134),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_5_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_5_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22093),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_5_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_5_15_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_5_15_6  (
            .in0(N__24594),
            .in1(N__22296),
            .in2(_gnd_net_),
            .in3(N__24541),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_5_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27967),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48803),
            .ce(N__25134),
            .sr(N__48219));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_5_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_5_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_5_16_3 .LUT_INIT=16'b1000101010001111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_5_16_3  (
            .in0(N__23746),
            .in1(N__25677),
            .in2(N__25558),
            .in3(N__25294),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48803),
            .ce(N__25134),
            .sr(N__48219));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_5_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_5_17_0 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_5_17_0  (
            .in0(N__23913),
            .in1(_gnd_net_),
            .in2(N__23890),
            .in3(N__23937),
            .lcout(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_5_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_5_17_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(N__24032),
            .in2(_gnd_net_),
            .in3(N__24077),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_5_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_5_17_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_5_17_2  (
            .in0(N__23690),
            .in1(N__23730),
            .in2(N__22072),
            .in3(N__23765),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_5_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_5_17_3 .LUT_INIT=16'b1111010111110001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_5_17_3  (
            .in0(N__23816),
            .in1(N__23844),
            .in2(N__22165),
            .in3(N__22162),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_5_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_5_17_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_5_17_4  (
            .in0(N__24033),
            .in1(N__23729),
            .in2(N__23694),
            .in3(N__23764),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_5_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_5_17_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_5_17_5  (
            .in0(N__23817),
            .in1(N__23843),
            .in2(N__22156),
            .in3(N__24078),
            .lcout(\current_shift_inst.PI_CTRL.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28450),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48785),
            .ce(N__25135),
            .sr(N__48226));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28012),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48785),
            .ce(N__25135),
            .sr(N__48226));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28147),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48785),
            .ce(N__25135),
            .sr(N__48226));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28801),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48785),
            .ce(N__25135),
            .sr(N__48226));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_5_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28060),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48785),
            .ce(N__25135),
            .sr(N__48226));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_5_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28369),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48785),
            .ce(N__25135),
            .sr(N__48226));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28723),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48776),
            .ce(N__25145),
            .sr(N__48231));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_5_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_5_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_5_19_2 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_5_19_2  (
            .in0(N__24103),
            .in1(N__25696),
            .in2(N__25550),
            .in3(N__25336),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48776),
            .ce(N__25145),
            .sr(N__48231));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_5_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28612),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48776),
            .ce(N__25145),
            .sr(N__48231));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_5_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28332),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48776),
            .ce(N__25145),
            .sr(N__48231));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_5_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_5_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_5_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28537),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48776),
            .ce(N__25145),
            .sr(N__48231));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_5_19_7  (
            .in0(N__29074),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48776),
            .ce(N__25145),
            .sr(N__48231));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_5_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28293),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48767),
            .ce(N__25178),
            .sr(N__48234));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_5_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29032),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48758),
            .ce(N__25194),
            .sr(N__48237));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_5_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27343),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48751),
            .ce(N__25179),
            .sr(N__48240));
    defparam \pwm_generator_inst.threshold_0_LC_7_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_7_7_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_7_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22384),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48855),
            .ce(),
            .sr(N__48139));
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_7_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_7_8_2 .LUT_INIT=16'b1011101111110011;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_6_LC_7_8_2  (
            .in0(N__29122),
            .in1(N__33456),
            .in2(N__35313),
            .in3(N__33633),
            .lcout(measured_delay_hc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48849),
            .ce(),
            .sr(N__48145));
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_7_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_7_9_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_21_LC_7_9_0  (
            .in0(N__24369),
            .in1(N__33650),
            .in2(_gnd_net_),
            .in3(N__30480),
            .lcout(measured_delay_hc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48843),
            .ce(),
            .sr(N__48150));
    defparam \pwm_generator_inst.threshold_5_LC_7_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_7_9_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_7_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22375),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48843),
            .ce(),
            .sr(N__48150));
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_7_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_7_9_3 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_2_LC_7_9_3  (
            .in0(N__33649),
            .in1(N__29209),
            .in2(N__35378),
            .in3(N__33460),
            .lcout(measured_delay_hc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48843),
            .ce(),
            .sr(N__48150));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_7_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_7_12_0 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_7_12_0  (
            .in0(N__35986),
            .in1(N__35790),
            .in2(N__36451),
            .in3(N__36614),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48820),
            .ce(N__24626),
            .sr(N__48179));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_7_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_7_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_7_12_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_7_12_2  (
            .in0(N__36443),
            .in1(N__35889),
            .in2(_gnd_net_),
            .in3(N__36611),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48820),
            .ce(N__24626),
            .sr(N__48179));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_7_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_7_12_6 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_7_12_6  (
            .in0(N__36444),
            .in1(N__33258),
            .in2(_gnd_net_),
            .in3(N__36612),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48820),
            .ce(N__24626),
            .sr(N__48179));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_7_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_7_12_7 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_7_12_7  (
            .in0(N__36613),
            .in1(N__36445),
            .in2(_gnd_net_),
            .in3(N__33210),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48820),
            .ce(N__24626),
            .sr(N__48179));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_7_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_7_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__22810),
            .in2(N__22300),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_7_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_7_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__22561),
            .in2(_gnd_net_),
            .in3(N__22531),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_7_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_7_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__23185),
            .in2(N__22528),
            .in3(N__22495),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_7_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_7_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__22492),
            .in2(_gnd_net_),
            .in3(N__22462),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_7_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_7_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__22459),
            .in2(_gnd_net_),
            .in3(N__22429),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_7_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_7_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__22426),
            .in2(_gnd_net_),
            .in3(N__22396),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_7_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_7_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__23250),
            .in2(_gnd_net_),
            .in3(N__22393),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_7_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_7_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__23229),
            .in2(_gnd_net_),
            .in3(N__22390),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_7_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_7_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__23199),
            .in2(_gnd_net_),
            .in3(N__22387),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_7_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_7_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__22768),
            .in2(_gnd_net_),
            .in3(N__22744),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_7_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_7_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__22741),
            .in2(_gnd_net_),
            .in3(N__22717),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_7_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_7_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__22714),
            .in2(_gnd_net_),
            .in3(N__22690),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_7_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_7_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__22687),
            .in2(_gnd_net_),
            .in3(N__22660),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_7_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_7_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__22657),
            .in2(_gnd_net_),
            .in3(N__22633),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_7_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_7_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__22630),
            .in2(_gnd_net_),
            .in3(N__22603),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_7_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_7_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__23646),
            .in2(_gnd_net_),
            .in3(N__22600),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_7_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_7_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__22597),
            .in2(_gnd_net_),
            .in3(N__22564),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_7_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_7_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__22879),
            .in2(_gnd_net_),
            .in3(N__22846),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_7_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_7_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__22843),
            .in2(_gnd_net_),
            .in3(N__22825),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__24586),
            .in2(_gnd_net_),
            .in3(N__24542),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_7_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_7_15_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__23438),
            .in2(_gnd_net_),
            .in3(N__23306),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_7_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_7_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_7_16_0  (
            .in0(N__24968),
            .in1(N__24922),
            .in2(N__24901),
            .in3(N__24821),
            .lcout(\current_shift_inst.PI_CTRL.N_47_16 ),
            .ltout(\current_shift_inst.PI_CTRL.N_47_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_7_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_7_16_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_7_16_1  (
            .in0(N__22912),
            .in1(N__22789),
            .in2(N__22801),
            .in3(N__24183),
            .lcout(\current_shift_inst.PI_CTRL.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_7_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_7_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_7_17_0  (
            .in0(N__22924),
            .in1(N__22774),
            .in2(N__26542),
            .in3(N__22798),
            .lcout(\current_shift_inst.PI_CTRL.N_47_21 ),
            .ltout(\current_shift_inst.PI_CTRL.N_47_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_17_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_17_1  (
            .in0(N__25478),
            .in1(N__22783),
            .in2(N__22777),
            .in3(N__24168),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_7_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_7_17_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_7_17_3  (
            .in0(N__26646),
            .in1(N__26677),
            .in2(N__26613),
            .in3(N__26563),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_7_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_7_17_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_7_17_4  (
            .in0(N__26742),
            .in1(N__26820),
            .in2(N__26190),
            .in3(N__26783),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_17_5  (
            .in0(N__24169),
            .in1(N__24858),
            .in2(N__25526),
            .in3(N__22890),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_17_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_17_6  (
            .in0(N__22918),
            .in1(N__22908),
            .in2(N__22894),
            .in3(N__26206),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_17_7  (
            .in0(N__26205),
            .in1(N__24859),
            .in2(N__24179),
            .in3(N__22891),
            .lcout(\current_shift_inst.PI_CTRL.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_7_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_7_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_7_18_1 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_7_18_1  (
            .in0(N__24139),
            .in1(N__25622),
            .in2(N__25549),
            .in3(N__25293),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48768),
            .ce(N__25208),
            .sr(N__48220));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_7_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_7_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_7_18_3 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_7_18_3  (
            .in0(N__23992),
            .in1(N__25614),
            .in2(N__25547),
            .in3(N__25289),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48768),
            .ce(N__25208),
            .sr(N__48220));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_7_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_7_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_7_18_4 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_7_18_4  (
            .in0(N__25290),
            .in1(N__25509),
            .in2(N__25655),
            .in3(N__23980),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48768),
            .ce(N__25208),
            .sr(N__48220));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_7_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_7_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_7_18_5 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_7_18_5  (
            .in0(N__23947),
            .in1(N__25621),
            .in2(N__25548),
            .in3(N__25292),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48768),
            .ce(N__25208),
            .sr(N__48220));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_7_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_7_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_7_18_6 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_7_18_6  (
            .in0(N__25291),
            .in1(N__25510),
            .in2(N__25656),
            .in3(N__23971),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48768),
            .ce(N__25208),
            .sr(N__48220));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_7_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_7_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_7_19_2 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_7_19_2  (
            .in0(N__24115),
            .in1(N__25671),
            .in2(N__25545),
            .in3(N__25322),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48759),
            .ce(N__25173),
            .sr(N__48223));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_19_4 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_7_19_4  (
            .in0(N__24091),
            .in1(N__25672),
            .in2(N__25546),
            .in3(N__25323),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48759),
            .ce(N__25173),
            .sr(N__48223));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_7_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_7_19_5 .LUT_INIT=16'b1111001100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_7_19_5  (
            .in0(N__25324),
            .in1(N__25499),
            .in2(N__25697),
            .in3(N__24001),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48759),
            .ce(N__25173),
            .sr(N__48223));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_7_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_7_19_6 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_7_19_6  (
            .in0(N__24196),
            .in1(N__25670),
            .in2(N__25544),
            .in3(N__25321),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48759),
            .ce(N__25173),
            .sr(N__48223));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28485),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48752),
            .ce(N__25209),
            .sr(N__48227));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_7_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_7_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_7_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28572),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48752),
            .ce(N__25209),
            .sr(N__48227));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_20_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_7_20_5  (
            .in0(N__28407),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48752),
            .ce(N__25209),
            .sr(N__48227));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_7_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_7_20_6 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_7_20_6  (
            .in0(N__24211),
            .in1(N__25676),
            .in2(N__25521),
            .in3(N__25325),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48752),
            .ce(N__25209),
            .sr(N__48227));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_7_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_7_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28996),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48752),
            .ce(N__25209),
            .sr(N__48227));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_21_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_7_21_0  (
            .in0(N__28254),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48746),
            .ce(N__25195),
            .sr(N__48232));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_7_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_7_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__33781),
            .in2(_gnd_net_),
            .in3(N__29815),
            .lcout(\current_shift_inst.timer_s1.N_187_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_3_1 (
            .in0(N__23038),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48870),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_8_6_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_8_6_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_8_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_8_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23029),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48856),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_8_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_8_7_0 .LUT_INIT=16'b1111111010101110;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_17_LC_8_7_0  (
            .in0(N__30482),
            .in1(N__33249),
            .in2(N__33645),
            .in3(N__29671),
            .lcout(measured_delay_hc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48850),
            .ce(),
            .sr(N__48133));
    defparam \pwm_generator_inst.threshold_7_LC_8_7_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_8_7_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_8_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23020),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48850),
            .ce(),
            .sr(N__48133));
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_8_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_8_7_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_4_LC_8_7_6  (
            .in0(N__30483),
            .in1(N__35244),
            .in2(N__33646),
            .in3(N__29178),
            .lcout(measured_delay_hc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48850),
            .ce(),
            .sr(N__48133));
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_8_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_8_7_7 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_15_LC_8_7_7  (
            .in0(N__29275),
            .in1(N__33613),
            .in2(N__35663),
            .in3(N__30481),
            .lcout(measured_delay_hc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48850),
            .ce(),
            .sr(N__48133));
    defparam \pwm_generator_inst.threshold_2_LC_8_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_8_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_8_8_5  (
            .in0(N__23011),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48844),
            .ce(),
            .sr(N__48140));
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_8_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_8_8_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_20_LC_8_8_6  (
            .in0(N__24349),
            .in1(N__33651),
            .in2(_gnd_net_),
            .in3(N__30455),
            .lcout(measured_delay_hc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48844),
            .ce(),
            .sr(N__48140));
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_8_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_8_8_7 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_22_LC_8_8_7  (
            .in0(N__30456),
            .in1(_gnd_net_),
            .in2(N__33655),
            .in3(N__24329),
            .lcout(measured_delay_hc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48844),
            .ce(),
            .sr(N__48140));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_8_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_8_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_8_9_4  (
            .in0(N__24365),
            .in1(N__24347),
            .in2(N__24331),
            .in3(N__26066),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_3_LC_8_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_8_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23179),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48830),
            .ce(),
            .sr(N__48151));
    defparam \pwm_generator_inst.threshold_1_LC_8_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_8_10_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_8_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23164),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48830),
            .ce(),
            .sr(N__48151));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_8_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_8_11_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_8_11_2  (
            .in0(N__35662),
            .in1(N__36398),
            .in2(_gnd_net_),
            .in3(N__36526),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48821),
            .ce(N__24636),
            .sr(N__48156));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_8_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_8_11_5 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_8_11_5  (
            .in0(N__36396),
            .in1(N__33155),
            .in2(_gnd_net_),
            .in3(N__33130),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48821),
            .ce(N__24636),
            .sr(N__48156));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_8_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_8_11_6 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_8_11_6  (
            .in0(N__33370),
            .in1(N__36397),
            .in2(_gnd_net_),
            .in3(N__36525),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48821),
            .ce(N__24636),
            .sr(N__48156));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_8_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_8_12_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_8_12_0  (
            .in0(N__36419),
            .in1(N__35931),
            .in2(_gnd_net_),
            .in3(N__36564),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48811),
            .ce(N__24621),
            .sr(N__48165));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_8_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_8_12_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_8_12_1  (
            .in0(N__36565),
            .in1(N__36420),
            .in2(_gnd_net_),
            .in3(N__36027),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48811),
            .ce(N__24621),
            .sr(N__48165));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_8_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_8_12_5 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_8_12_5  (
            .in0(N__36566),
            .in1(N__36421),
            .in2(_gnd_net_),
            .in3(N__33310),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48811),
            .ce(N__24621),
            .sr(N__48165));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_13_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_13_0  (
            .in0(N__23440),
            .in1(N__23552),
            .in2(N__23344),
            .in3(N__23260),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48804),
            .ce(),
            .sr(N__48180));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_13_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_13_1  (
            .in0(N__23339),
            .in1(N__23442),
            .in2(N__23578),
            .in3(N__23236),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48804),
            .ce(),
            .sr(N__48180));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_13_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_13_2  (
            .in0(N__23441),
            .in1(N__23556),
            .in2(N__23345),
            .in3(N__23209),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48804),
            .ce(),
            .sr(N__48180));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_13_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_13_3  (
            .in0(N__23551),
            .in1(N__23439),
            .in2(_gnd_net_),
            .in3(N__23307),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_8_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_8_13_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_0_LC_8_13_7  (
            .in0(N__35827),
            .in1(N__33634),
            .in2(_gnd_net_),
            .in3(N__30490),
            .lcout(measured_delay_hc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48804),
            .ce(),
            .sr(N__48180));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_8_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_8_14_0 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_8_14_0  (
            .in0(N__24554),
            .in1(N__23340),
            .in2(N__23577),
            .in3(N__23465),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48793),
            .ce(N__31454),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_8_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_8_14_1 .LUT_INIT=16'b0100000001001010;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_8_14_1  (
            .in0(N__23464),
            .in1(N__23550),
            .in2(N__23374),
            .in3(N__24555),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48793),
            .ce(N__31454),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_8_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_8_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__24587),
            .in2(_gnd_net_),
            .in3(N__24553),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_8_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_8_14_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_8_14_4  (
            .in0(N__32896),
            .in1(N__32472),
            .in2(N__32733),
            .in3(N__32367),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48793),
            .ce(N__31454),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_8_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_8_15_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_8_15_0  (
            .in0(N__29926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29968),
            .lcout(),
            .ltout(\phase_controller_inst1.N_228_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_8_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_8_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_8_15_1 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_8_15_1  (
            .in0(N__23531),
            .in1(N__27532),
            .in2(N__23656),
            .in3(N__26110),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48786),
            .ce(),
            .sr(N__48196));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_15_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_15_6  (
            .in0(N__23444),
            .in1(N__23530),
            .in2(N__23346),
            .in3(N__23653),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48786),
            .ce(),
            .sr(N__48196));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_15_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_15_7  (
            .in0(N__23529),
            .in1(N__23443),
            .in2(_gnd_net_),
            .in3(N__23314),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_16_0 .LUT_INIT=16'b1010101100001011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_8_16_0  (
            .in0(N__24046),
            .in1(N__25252),
            .in2(N__25553),
            .in3(N__25651),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48777),
            .ce(N__25197),
            .sr(N__48204));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_16_1 .LUT_INIT=16'b1110000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_8_16_1  (
            .in0(N__25248),
            .in1(N__25527),
            .in2(N__24130),
            .in3(N__25652),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48777),
            .ce(N__25197),
            .sr(N__48204));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_8_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_8_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_8_16_2 .LUT_INIT=16'b1010101100001011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_8_16_2  (
            .in0(N__23704),
            .in1(N__25250),
            .in2(N__25552),
            .in3(N__25650),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48777),
            .ce(N__25197),
            .sr(N__48204));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_16_3 .LUT_INIT=16'b1100110100001101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_8_16_3  (
            .in0(N__25251),
            .in1(N__23662),
            .in2(N__25554),
            .in3(N__25654),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48777),
            .ce(N__25197),
            .sr(N__48204));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_8_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_8_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_8_16_6 .LUT_INIT=16'b1010100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_8_16_6  (
            .in0(N__23959),
            .in1(N__25247),
            .in2(N__25551),
            .in3(N__25649),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48777),
            .ce(N__25197),
            .sr(N__48204));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_8_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_8_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_8_16_7 .LUT_INIT=16'b1110000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_8_16_7  (
            .in0(N__25249),
            .in1(N__25528),
            .in2(N__23785),
            .in3(N__25653),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48777),
            .ce(N__25197),
            .sr(N__48204));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_8_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_8_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_8_17_0 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__23930),
            .in2(N__28179),
            .in3(N__23862),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ),
            .clk(N__48769),
            .ce(N__25207),
            .sr(N__48210));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_8_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_8_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_8_17_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_8_17_1  (
            .in0(N__23860),
            .in1(N__23912),
            .in2(N__28146),
            .in3(N__23893),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(N__48769),
            .ce(N__25207),
            .sr(N__48210));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_8_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_8_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_8_17_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_8_17_2  (
            .in0(N__23863),
            .in1(N__23885),
            .in2(N__28101),
            .in3(N__23866),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(N__48769),
            .ce(N__25207),
            .sr(N__48210));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_8_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_8_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_8_17_3 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_8_17_3  (
            .in0(N__23861),
            .in1(N__23842),
            .in2(N__28056),
            .in3(N__23821),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(N__48769),
            .ce(N__25207),
            .sr(N__48210));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_8_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_8_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__23796),
            .in2(N__28011),
            .in3(N__23776),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_8_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_8_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__23773),
            .in2(N__27963),
            .in3(N__23734),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_8_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_8_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__23720),
            .in2(N__28492),
            .in3(N__23698),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_8_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_8_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__23678),
            .in2(N__28449),
            .in3(N__24082),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_8_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_8_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__24073),
            .in2(N__28408),
            .in3(N__24037),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_8_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_8_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__24020),
            .in2(N__28368),
            .in3(N__23995),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_8_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_8_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__26248),
            .in2(N__28333),
            .in3(N__23983),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_8_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_8_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__26567),
            .in2(N__28294),
            .in3(N__23974),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_8_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_8_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__26776),
            .in2(N__28255),
            .in3(N__23965),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_8_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_8_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__26642),
            .in2(N__28219),
            .in3(N__23962),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_8_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_8_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__26687),
            .in2(N__28800),
            .in3(N__23950),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_8_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_8_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__26329),
            .in2(N__28761),
            .in3(N__23941),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_8_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_8_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__26602),
            .in2(N__28722),
            .in3(N__24190),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_8_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_8_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__28683),
            .in2(N__24825),
            .in3(N__24187),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_8_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_8_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__24167),
            .in2(N__28648),
            .in3(N__24133),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_8_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_8_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__24930),
            .in2(N__28611),
            .in3(N__24118),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_8_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_8_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__24964),
            .in2(N__28573),
            .in3(N__24109),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_8_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_8_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__26402),
            .in2(N__28536),
            .in3(N__24106),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_8_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_8_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__24899),
            .in2(N__29073),
            .in3(N__24094),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_8_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_8_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__26365),
            .in2(N__29031),
            .in3(N__24085),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_8_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_8_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__26482),
            .in2(N__28995),
            .in3(N__24226),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_8_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_8_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(N__26518),
            .in2(N__27344),
            .in3(N__24223),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_8_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_8_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__27333),
            .in2(N__26440),
            .in3(N__24220),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_8_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_8_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__26809),
            .in2(N__27345),
            .in3(N__24217),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_8_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_8_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__27337),
            .in2(N__26738),
            .in3(N__24214),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_8_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_8_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_8_20_5  (
            .in0(_gnd_net_),
            .in1(N__26284),
            .in2(N__27346),
            .in3(N__24205),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_8_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_8_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(N__27341),
            .in2(N__26180),
            .in3(N__24202),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_8_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_8_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_8_20_7  (
            .in0(N__27342),
            .in1(N__25401),
            .in2(_gnd_net_),
            .in3(N__24199),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.start_timer_s1_LC_8_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_8_21_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.start_timer_s1_LC_8_21_4 .LUT_INIT=16'b0111001111110000;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_8_21_4  (
            .in0(N__24269),
            .in1(N__25805),
            .in2(N__29877),
            .in3(N__27928),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48740),
            .ce(N__31432),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_LC_8_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_8_21_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.stop_timer_s1_LC_8_21_5 .LUT_INIT=16'b1111110111001100;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_8_21_5  (
            .in0(N__27929),
            .in1(N__24283),
            .in2(N__25812),
            .in3(N__29822),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48740),
            .ce(N__31432),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_8_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_8_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_8_22_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.stop_timer_s1_RNO_0_LC_8_22_3  (
            .in0(N__24255),
            .in1(N__25793),
            .in2(N__29878),
            .in3(N__27927),
            .lcout(\current_shift_inst.N_199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.meas_state_0_LC_8_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.meas_state_0_LC_8_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.meas_state_0_LC_8_23_3 .LUT_INIT=16'b0111111110101010;
    LogicCell40 \current_shift_inst.meas_state_0_LC_8_23_3  (
            .in0(N__27937),
            .in1(N__24262),
            .in2(N__29879),
            .in3(N__25794),
            .lcout(\current_shift_inst.meas_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48728),
            .ce(),
            .sr(N__48235));
    defparam \current_shift_inst.phase_valid_LC_8_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.phase_valid_LC_8_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.phase_valid_LC_8_23_4 .LUT_INIT=16'b1010100011111000;
    LogicCell40 \current_shift_inst.phase_valid_LC_8_23_4  (
            .in0(N__25795),
            .in1(N__25757),
            .in2(N__24270),
            .in3(N__27936),
            .lcout(\current_shift_inst.phase_validZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48728),
            .ce(),
            .sr(N__48235));
    defparam \delay_measurement_inst.hc_state_0_LC_9_5_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_0_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_state_0_LC_9_5_6 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.hc_state_0_LC_9_5_6  (
            .in0(N__26006),
            .in1(N__25988),
            .in2(_gnd_net_),
            .in3(N__25969),
            .lcout(\delay_measurement_inst.hc_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48857),
            .ce(N__31465),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_9_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_hc_LC_9_6_7 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_9_6_7  (
            .in0(N__25972),
            .in1(N__26008),
            .in2(_gnd_net_),
            .in3(N__25989),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48851),
            .ce(),
            .sr(N__48124));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_7_0 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_7_0  (
            .in0(N__25893),
            .in1(N__27273),
            .in2(_gnd_net_),
            .in3(N__30172),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_337_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_9_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_9_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_9_7_5  (
            .in0(N__30358),
            .in1(N__29204),
            .in2(N__29149),
            .in3(N__29226),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_9_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_9_8_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_9_8_1  (
            .in0(N__29528),
            .in1(N__29179),
            .in2(N__29497),
            .in3(N__29269),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_9_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_9_8_2 .LUT_INIT=16'b0000111011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_9_8_2  (
            .in0(N__29270),
            .in1(N__29456),
            .in2(N__24235),
            .in3(N__24232),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_9_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_9_8_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_9_8_7  (
            .in0(N__24373),
            .in1(N__24348),
            .in2(N__24330),
            .in3(N__33115),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto30_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_9_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_9_9_0 .LUT_INIT=16'b1101100011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_9_LC_9_9_0  (
            .in0(N__33621),
            .in1(N__29461),
            .in2(N__35984),
            .in3(N__33445),
            .lcout(measured_delay_hc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48831),
            .ce(),
            .sr(N__48141));
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_9_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_9_9_2 .LUT_INIT=16'b1010110011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_19_LC_9_9_2  (
            .in0(N__29617),
            .in1(N__26068),
            .in2(N__33647),
            .in3(N__33442),
            .lcout(measured_delay_hc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48831),
            .ce(),
            .sr(N__48141));
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_9_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_9_9_3 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_12_LC_9_9_3  (
            .in0(N__33411),
            .in1(N__33622),
            .in2(N__29353),
            .in3(N__30437),
            .lcout(measured_delay_hc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48831),
            .ce(),
            .sr(N__48141));
    defparam \pwm_generator_inst.threshold_4_LC_9_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_9_9_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_9_9_4  (
            .in0(N__24307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48831),
            .ce(),
            .sr(N__48141));
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_9_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_9_9_6 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_8_LC_9_9_6  (
            .in0(N__33620),
            .in1(N__29496),
            .in2(N__36495),
            .in3(N__33444),
            .lcout(measured_delay_hc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48831),
            .ce(),
            .sr(N__48141));
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_9_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_9_9_7 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_7_LC_9_9_7  (
            .in0(N__33443),
            .in1(N__29530),
            .in2(N__35423),
            .in3(N__33626),
            .lcout(measured_delay_hc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48831),
            .ce(),
            .sr(N__48141));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_9_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_9_10_4 .LUT_INIT=16'b0000110001001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_9_10_4  (
            .in0(N__35658),
            .in1(N__24295),
            .in2(N__26050),
            .in3(N__24517),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_9_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_9_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_9_10_5  (
            .in0(N__35370),
            .in1(N__35691),
            .in2(N__36086),
            .in3(N__35837),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_9_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_9_10_6 .LUT_INIT=16'b1100110010001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto6_LC_9_10_6  (
            .in0(N__36129),
            .in1(N__35315),
            .in2(N__24286),
            .in3(N__35254),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlt8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_9_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_9_10_7 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_9_10_7  (
            .in0(N__33365),
            .in1(N__35967),
            .in2(N__24520),
            .in3(N__26074),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__24493),
            .in2(N__24511),
            .in3(N__27660),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_11_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_11_1  (
            .in0(N__27605),
            .in1(N__24478),
            .in2(N__24487),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__24457),
            .in2(N__24472),
            .in3(N__27642),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__24442),
            .in2(N__24451),
            .in3(N__27584),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__24424),
            .in2(N__24436),
            .in3(N__27623),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__24403),
            .in2(N__24418),
            .in3(N__27719),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__24379),
            .in2(N__24397),
            .in3(N__27737),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__24754),
            .in2(N__24772),
            .in3(N__27755),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__24730),
            .in2(N__24748),
            .in3(N__27774),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__24706),
            .in2(N__24724),
            .in3(N__27792),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_9_12_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_9_12_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_9_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24700),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48805),
            .ce(),
            .sr(N__48157));
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_9_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_9_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_9_13_4 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_9_13_4  (
            .in0(N__35323),
            .in1(N__35769),
            .in2(N__36442),
            .in3(N__36561),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48794),
            .ce(N__24622),
            .sr(N__48166));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_9_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_9_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_9_13_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_9_13_5  (
            .in0(N__36563),
            .in1(N__36418),
            .in2(_gnd_net_),
            .in3(N__35424),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48794),
            .ce(N__24622),
            .sr(N__48166));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_13_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_9_13_7  (
            .in0(N__36562),
            .in1(N__36417),
            .in2(_gnd_net_),
            .in3(N__33407),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48794),
            .ce(N__24622),
            .sr(N__48166));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_9_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_9_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_9_15_6 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_9_15_6  (
            .in0(N__29970),
            .in1(N__24595),
            .in2(N__24565),
            .in3(N__24556),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48778),
            .ce(),
            .sr(N__48188));
    defparam \phase_controller_inst1.state_2_LC_9_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_9_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_9_15_7 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst1.state_2_LC_9_15_7  (
            .in0(N__29969),
            .in1(N__39583),
            .in2(N__29936),
            .in3(N__26139),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48778),
            .ce(),
            .sr(N__48188));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_9_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_9_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_9_16_0  (
            .in0(N__24973),
            .in1(N__24923),
            .in2(N__24900),
            .in3(N__24811),
            .lcout(\current_shift_inst.PI_CTRL.N_46_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_9_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_9_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__39643),
            .in2(_gnd_net_),
            .in3(N__39549),
            .lcout(\phase_controller_inst1.N_231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_17_2 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_9_17_2  (
            .in0(N__25657),
            .in1(N__24844),
            .in2(N__25522),
            .in3(N__25326),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48760),
            .ce(N__25210),
            .sr(N__48205));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_17_5 .LUT_INIT=16'b1110000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_9_17_5  (
            .in0(N__25327),
            .in1(N__25466),
            .in2(N__24838),
            .in3(N__25658),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48760),
            .ce(N__25210),
            .sr(N__48205));
    defparam \current_shift_inst.start_timer_phase_LC_9_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_phase_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.start_timer_phase_LC_9_18_5 .LUT_INIT=16'b0011101100101010;
    LogicCell40 \current_shift_inst.start_timer_phase_LC_9_18_5  (
            .in0(N__31784),
            .in1(N__25813),
            .in2(N__25765),
            .in3(N__27915),
            .lcout(\current_shift_inst.start_timer_phaseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48753),
            .ce(N__31444),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_9_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_9_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_9_19_1 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_9_19_1  (
            .in0(N__24790),
            .in1(N__25698),
            .in2(N__25476),
            .in3(N__25328),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48747),
            .ce(N__25174),
            .sr(N__48215));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_9_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_9_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_9_19_4 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_9_19_4  (
            .in0(N__25330),
            .in1(N__25421),
            .in2(N__25708),
            .in3(N__24784),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48747),
            .ce(N__25174),
            .sr(N__48215));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_9_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_9_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_9_19_5 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_9_19_5  (
            .in0(N__24778),
            .in1(N__25699),
            .in2(N__25477),
            .in3(N__25329),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48747),
            .ce(N__25174),
            .sr(N__48215));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_9_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_9_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_9_20_1 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_9_20_1  (
            .in0(N__25706),
            .in1(N__25738),
            .in2(N__25474),
            .in3(N__25334),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48741),
            .ce(N__25196),
            .sr(N__48221));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_9_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_9_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_9_20_2 .LUT_INIT=16'b1110000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_9_20_2  (
            .in0(N__25332),
            .in1(N__25410),
            .in2(N__25732),
            .in3(N__25704),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48741),
            .ce(N__25196),
            .sr(N__48221));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_9_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_9_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_9_20_4 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_9_20_4  (
            .in0(N__25335),
            .in1(N__25723),
            .in2(N__25475),
            .in3(N__25707),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48741),
            .ce(N__25196),
            .sr(N__48221));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_9_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_9_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_9_20_5 .LUT_INIT=16'b1111010011000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_9_20_5  (
            .in0(N__25705),
            .in1(N__25417),
            .in2(N__25717),
            .in3(N__25333),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48741),
            .ce(N__25196),
            .sr(N__48221));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_9_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_9_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_9_20_7 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_9_20_7  (
            .in0(N__25703),
            .in1(N__25564),
            .in2(N__25473),
            .in3(N__25331),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48741),
            .ce(N__25196),
            .sr(N__48221));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_9_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_9_21_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__40419),
            .in2(_gnd_net_),
            .in3(N__34357),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNILORI_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_9_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_9_21_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_9_21_3  (
            .in0(N__40564),
            .in1(N__40503),
            .in2(N__34444),
            .in3(N__34401),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_9_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_9_21_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__40563),
            .in2(_gnd_net_),
            .in3(N__34440),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_9_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_9_21_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__40265),
            .in2(_gnd_net_),
            .in3(N__34275),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_9_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_9_22_0 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_9_22_0  (
            .in0(N__33916),
            .in1(N__39930),
            .in2(N__40701),
            .in3(N__34522),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_9_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_9_22_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_9_22_1  (
            .in0(N__39929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33915),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_9_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_9_22_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_9_22_2  (
            .in0(N__40697),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34521),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_9_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_9_22_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__39990),
            .in2(_gnd_net_),
            .in3(N__33960),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_9_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_9_22_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_9_22_4  (
            .in0(N__34600),
            .in1(N__40764),
            .in2(N__34642),
            .in3(N__41721),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync0_LC_9_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync0_LC_9_22_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync0_LC_9_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S3_sync0_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45684),
            .lcout(\current_shift_inst.S3_syncZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48729),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_9_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_9_22_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_9_22_7  (
            .in0(N__32810),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32509),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_phase_LC_9_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_phase_LC_9_23_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.stop_timer_phase_LC_9_23_4 .LUT_INIT=16'b1101110111000000;
    LogicCell40 \current_shift_inst.stop_timer_phase_LC_9_23_4  (
            .in0(N__27930),
            .in1(N__25801),
            .in2(N__25761),
            .in3(N__31750),
            .lcout(\current_shift_inst.stop_timer_phaseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48721),
            .ce(N__31412),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_9_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_9_23_5 .LUT_INIT=16'b0000100001011000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_9_23_5  (
            .in0(N__32851),
            .in1(N__32731),
            .in2(N__32596),
            .in3(N__32360),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48721),
            .ce(N__31412),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_rise_LC_9_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.S3_rise_LC_9_24_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_rise_LC_9_24_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \current_shift_inst.S3_rise_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__25840),
            .in2(_gnd_net_),
            .in3(N__25848),
            .lcout(\current_shift_inst.S3_riseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48714),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync1_LC_9_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync1_LC_9_24_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync1_LC_9_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S3_sync1_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25858),
            .lcout(\current_shift_inst.S3_syncZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48714),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync_prev_LC_9_24_6 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync_prev_LC_9_24_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync_prev_LC_9_24_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.S3_sync_prev_LC_9_24_6  (
            .in0(N__25849),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.S3_sync_prevZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48714),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_ibuf_gb_io_RNI79U7_LC_9_29_3.C_ON=1'b0;
    defparam reset_ibuf_gb_io_RNI79U7_LC_9_29_3.SEQ_MODE=4'b0000;
    defparam reset_ibuf_gb_io_RNI79U7_LC_9_29_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 reset_ibuf_gb_io_RNI79U7_LC_9_29_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48276),
            .lcout(red_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_10_3_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_10_3_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_10_3_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_10_3_2 (
            .in0(N__25834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48858),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC2_LC_10_4_4.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC2_LC_10_4_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC2_LC_10_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC2_LC_10_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37966),
            .lcout(delay_hc_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48852),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.prev_hc_sig_LC_10_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_hc_sig_LC_10_5_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_hc_sig_LC_10_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_hc_sig_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25970),
            .lcout(\delay_measurement_inst.prev_hc_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48845),
            .ce(),
            .sr(N__48101));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_10_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_10_6_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__25944),
            .in2(_gnd_net_),
            .in3(N__25917),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_10_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_10_6_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_10_6_2  (
            .in0(N__25881),
            .in1(N__25905),
            .in2(N__25822),
            .in3(N__25819),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_10_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_10_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_10_6_3  (
            .in0(N__25869),
            .in1(N__27231),
            .in2(N__25933),
            .in3(N__27243),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_10_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_hc_LC_10_6_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_10_6_4  (
            .in0(N__26007),
            .in1(N__25990),
            .in2(N__48280),
            .in3(N__25971),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48839),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_10_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_10_7_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_10_7_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_26_LC_10_7_0  (
            .in0(N__25945),
            .in1(N__33558),
            .in2(_gnd_net_),
            .in3(N__30425),
            .lcout(measured_delay_hc_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48832),
            .ce(),
            .sr(N__48117));
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_10_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_10_7_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_30_LC_10_7_1  (
            .in0(N__30427),
            .in1(N__25932),
            .in2(_gnd_net_),
            .in3(N__33561),
            .lcout(measured_delay_hc_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48832),
            .ce(),
            .sr(N__48117));
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_10_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_10_7_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_25_LC_10_7_2  (
            .in0(N__25918),
            .in1(N__33557),
            .in2(_gnd_net_),
            .in3(N__30424),
            .lcout(measured_delay_hc_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48832),
            .ce(),
            .sr(N__48117));
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_10_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_10_7_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_5_LC_10_7_3  (
            .in0(N__30428),
            .in1(N__33559),
            .in2(N__36139),
            .in3(N__29148),
            .lcout(measured_delay_hc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48832),
            .ce(),
            .sr(N__48117));
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_10_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_10_7_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_23_LC_10_7_4  (
            .in0(N__25906),
            .in1(N__33555),
            .in2(_gnd_net_),
            .in3(N__30422),
            .lcout(measured_delay_hc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48832),
            .ce(),
            .sr(N__48117));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_7_5 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_10_7_5  (
            .in0(N__27274),
            .in1(N__25894),
            .in2(_gnd_net_),
            .in3(N__30173),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48832),
            .ce(),
            .sr(N__48117));
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_10_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_10_7_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_10_7_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_24_LC_10_7_6  (
            .in0(N__25882),
            .in1(N__33556),
            .in2(_gnd_net_),
            .in3(N__30423),
            .lcout(measured_delay_hc_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48832),
            .ce(),
            .sr(N__48117));
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_10_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_10_7_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_29_LC_10_7_7  (
            .in0(N__30426),
            .in1(N__25870),
            .in2(_gnd_net_),
            .in3(N__33560),
            .lcout(measured_delay_hc_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48832),
            .ce(),
            .sr(N__48117));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_10_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_10_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_10_8_0  (
            .in0(N__29495),
            .in1(N__29529),
            .in2(N__29121),
            .in3(N__29271),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_10_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_10_8_1 .LUT_INIT=16'b0100110001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_10_8_1  (
            .in0(N__26017),
            .in1(N__27481),
            .in2(N__26035),
            .in3(N__26032),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_10_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_10_8_2 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_10_8_2  (
            .in0(N__27378),
            .in1(N__27452),
            .in2(N__26026),
            .in3(N__29721),
            .lcout(\delay_measurement_inst.delay_hc_reg3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_10_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_10_8_3 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_10_8_3  (
            .in0(N__27453),
            .in1(N__27379),
            .in2(N__29725),
            .in3(N__26023),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_10_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_10_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_10_8_4  (
            .in0(N__29379),
            .in1(N__29415),
            .in2(N__29352),
            .in3(N__29307),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOHNN2_6_LC_10_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOHNN2_6_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOHNN2_6_LC_10_8_5 .LUT_INIT=16'b0011000010110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOHNN2_6_LC_10_8_5  (
            .in0(N__27409),
            .in1(N__29457),
            .in2(N__26011),
            .in3(N__29117),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_10_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_10_9_1 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_10_9_1 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_1_LC_10_9_1  (
            .in0(N__33544),
            .in1(N__29227),
            .in2(N__35709),
            .in3(N__33441),
            .lcout(measured_delay_hc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48813),
            .ce(),
            .sr(N__48128));
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_10_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_10_9_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_11_LC_10_9_3  (
            .in0(N__30419),
            .in1(N__29383),
            .in2(N__33602),
            .in3(N__35888),
            .lcout(measured_delay_hc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48813),
            .ce(),
            .sr(N__48128));
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_10_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_10_9_5 .LUT_INIT=16'b1111111010101110;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_18_LC_10_9_5  (
            .in0(N__30421),
            .in1(N__33208),
            .in2(N__33604),
            .in3(N__29644),
            .lcout(measured_delay_hc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48813),
            .ce(),
            .sr(N__48128));
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_10_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_10_9_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_10_9_6 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_10_LC_10_9_6  (
            .in0(N__35930),
            .in1(N__33545),
            .in2(N__29419),
            .in3(N__30418),
            .lcout(measured_delay_hc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48813),
            .ce(),
            .sr(N__48128));
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_10_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_10_9_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_10_9_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_13_LC_10_9_7  (
            .in0(N__30420),
            .in1(N__36018),
            .in2(N__33603),
            .in3(N__29311),
            .lcout(measured_delay_hc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48813),
            .ce(),
            .sr(N__48128));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_10_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_10_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_10_10_0  (
            .in0(N__33393),
            .in1(N__35868),
            .in2(N__36019),
            .in3(N__35910),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_10_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_10_10_1 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_10_10_1  (
            .in0(N__36477),
            .in1(N__35403),
            .in2(N__26077),
            .in3(N__35966),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_10_10_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_10_10_7  (
            .in0(N__33254),
            .in1(N__26067),
            .in2(N__33204),
            .in3(N__33307),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_10_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_10_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_10_11_0  (
            .in0(N__36020),
            .in1(N__35664),
            .in2(N__33308),
            .in3(N__33369),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_10_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_10_11_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_10_11_1  (
            .in0(N__36490),
            .in1(N__35416),
            .in2(N__36149),
            .in3(N__35923),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_10_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_10_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_10_11_2  (
            .in0(N__33253),
            .in1(N__33406),
            .in2(N__33209),
            .in3(N__35881),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_10_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_10_12_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_10_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_10_12_0  (
            .in0(N__27697),
            .in1(N__27661),
            .in2(_gnd_net_),
            .in3(N__26041),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__48788),
            .ce(),
            .sr(N__48146));
    defparam \pwm_generator_inst.counter_1_LC_10_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_10_12_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_10_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_10_12_1  (
            .in0(N__27691),
            .in1(N__27607),
            .in2(_gnd_net_),
            .in3(N__26038),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__48788),
            .ce(),
            .sr(N__48146));
    defparam \pwm_generator_inst.counter_2_LC_10_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_10_12_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_10_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_10_12_2  (
            .in0(N__27698),
            .in1(N__27643),
            .in2(_gnd_net_),
            .in3(N__26101),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__48788),
            .ce(),
            .sr(N__48146));
    defparam \pwm_generator_inst.counter_3_LC_10_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_10_12_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_10_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_10_12_3  (
            .in0(N__27692),
            .in1(N__27586),
            .in2(_gnd_net_),
            .in3(N__26098),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__48788),
            .ce(),
            .sr(N__48146));
    defparam \pwm_generator_inst.counter_4_LC_10_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_10_12_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_10_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_10_12_4  (
            .in0(N__27699),
            .in1(N__27625),
            .in2(_gnd_net_),
            .in3(N__26095),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__48788),
            .ce(),
            .sr(N__48146));
    defparam \pwm_generator_inst.counter_5_LC_10_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_10_12_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_10_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_10_12_5  (
            .in0(N__27693),
            .in1(N__27720),
            .in2(_gnd_net_),
            .in3(N__26092),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__48788),
            .ce(),
            .sr(N__48146));
    defparam \pwm_generator_inst.counter_6_LC_10_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_10_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_10_12_6  (
            .in0(N__27700),
            .in1(N__27738),
            .in2(_gnd_net_),
            .in3(N__26089),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__48788),
            .ce(),
            .sr(N__48146));
    defparam \pwm_generator_inst.counter_7_LC_10_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_10_12_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_10_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_10_12_7  (
            .in0(N__27694),
            .in1(N__27757),
            .in2(_gnd_net_),
            .in3(N__26086),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__48788),
            .ce(),
            .sr(N__48146));
    defparam \pwm_generator_inst.counter_8_LC_10_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_10_13_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_10_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_10_13_0  (
            .in0(N__27696),
            .in1(N__27775),
            .in2(_gnd_net_),
            .in3(N__26083),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__48780),
            .ce(),
            .sr(N__48152));
    defparam \pwm_generator_inst.counter_9_LC_10_13_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_10_13_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_10_13_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_10_13_1  (
            .in0(N__27793),
            .in1(N__27695),
            .in2(_gnd_net_),
            .in3(N__26080),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48780),
            .ce(),
            .sr(N__48152));
    defparam \phase_controller_inst1.state_RNO_0_3_LC_10_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_10_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNO_0_3_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__31021),
            .in2(_gnd_net_),
            .in3(N__27526),
            .lcout(),
            .ltout(\phase_controller_inst1.N_232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_10_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_10_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_10_14_3 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst1.state_3_LC_10_14_3  (
            .in0(N__39584),
            .in1(N__26143),
            .in2(N__26146),
            .in3(N__27552),
            .lcout(\phase_controller_inst1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48771),
            .ce(),
            .sr(N__48158));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_15_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_15_3  (
            .in0(N__41190),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34866),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI190J_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_15_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__39579),
            .in2(_gnd_net_),
            .in3(N__26138),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_10_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_10_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__40504),
            .in2(_gnd_net_),
            .in3(N__34400),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_10_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_10_16_0 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_10_16_0  (
            .in0(N__34554),
            .in1(N__41728),
            .in2(N__41661),
            .in3(N__34596),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_10_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_10_16_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_10_16_1  (
            .in0(N__40843),
            .in1(N__40770),
            .in2(N__34686),
            .in3(N__34628),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_10_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_10_16_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_10_16_2  (
            .in0(N__41047),
            .in1(N__34749),
            .in2(N__34801),
            .in3(N__40984),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_10_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_10_16_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__40771),
            .in2(_gnd_net_),
            .in3(N__34627),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_16_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_16_4  (
            .in0(N__41191),
            .in1(N__34834),
            .in2(N__34873),
            .in3(N__41111),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_10_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_10_16_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_10_16_5  (
            .in0(N__32626),
            .in1(N__32852),
            .in2(_gnd_net_),
            .in3(N__32499),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_10_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_10_16_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__41727),
            .in2(_gnd_net_),
            .in3(N__34595),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_10_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_10_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_10_17_0  (
            .in0(N__26691),
            .in1(N__26641),
            .in2(N__26617),
            .in3(N__26575),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_10_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_10_17_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_10_17_2  (
            .in0(N__34276),
            .in1(N__40194),
            .in2(N__40276),
            .in3(N__34232),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_10_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_10_17_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_10_17_3  (
            .in0(N__26526),
            .in1(N__26491),
            .in2(N__26454),
            .in3(N__26406),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_10_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_10_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(N__41247),
            .in2(_gnd_net_),
            .in3(N__34959),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_10_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_10_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_10_18_2  (
            .in0(N__26525),
            .in1(N__26489),
            .in2(N__26453),
            .in3(N__26401),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_10_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_10_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_10_18_3  (
            .in0(N__26377),
            .in1(N__26336),
            .in2(N__26302),
            .in3(N__26255),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_10_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_10_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_10_18_4  (
            .in0(N__26221),
            .in1(N__26215),
            .in2(N__26209),
            .in3(N__26704),
            .lcout(\current_shift_inst.PI_CTRL.N_46_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_10_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_10_18_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_10_18_5  (
            .in0(N__26176),
            .in1(N__26821),
            .in2(N__26785),
            .in3(N__26728),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_10_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_10_18_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__40842),
            .in2(_gnd_net_),
            .in3(N__34685),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_18_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_18_7  (
            .in0(N__37362),
            .in1(N__40058),
            .in2(_gnd_net_),
            .in3(N__34001),
            .lcout(\current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_19_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__40342),
            .in2(_gnd_net_),
            .in3(N__34312),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_10_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_10_19_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__38884),
            .in2(_gnd_net_),
            .in3(N__36822),
            .lcout(\phase_controller_inst1.stoper_tr.N_21 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_10_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_10_19_3 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26698),
            .in3(N__45154),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_19_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__40195),
            .in2(_gnd_net_),
            .in3(N__34234),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_10_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_10_19_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_10_19_5  (
            .in0(N__40983),
            .in1(N__40905),
            .in2(N__34759),
            .in3(N__34723),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_10_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_10_19_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__40982),
            .in2(_gnd_net_),
            .in3(N__34755),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_10_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_10_19_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_10_19_7  (
            .in0(N__34486),
            .in1(N__40562),
            .in2(N__40636),
            .in3(N__34439),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_10_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_10_20_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_10_20_1  (
            .in0(N__34108),
            .in1(N__37444),
            .in2(_gnd_net_),
            .in3(N__37329),
            .lcout(\current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_20_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__40059),
            .in2(_gnd_net_),
            .in3(N__34002),
            .lcout(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_20_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_20_3  (
            .in0(N__40060),
            .in1(N__39989),
            .in2(N__34006),
            .in3(N__33953),
            .lcout(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_10_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_10_20_6 .LUT_INIT=16'b1001110010011100;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_10_20_6  (
            .in0(N__37330),
            .in1(N__37294),
            .in2(N__37450),
            .in3(N__34069),
            .lcout(\current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_10_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_10_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__37448),
            .in2(N__37449),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_10_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_10_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__26857),
            .in2(N__34171),
            .in3(N__34893),
            .lcout(\current_shift_inst.z_i_0_31 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_10_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_10_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_1_c_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__34107),
            .in2(N__26851),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_0 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_10_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_10_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_2_c_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__34065),
            .in2(N__26839),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_1 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_10_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_10_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__34033),
            .in2(N__26830),
            .in3(N__37465),
            .lcout(\current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_2 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_10_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_10_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_4_c_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__26977),
            .in2(N__37363),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_3 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_10_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_10_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__26968),
            .in2(N__26959),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_4 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_10_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_10_21_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__30079),
            .in2(N__26947),
            .in3(N__26938),
            .lcout(\current_shift_inst.control_input_1_axb_0 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_5 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_10_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_10_22_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__26935),
            .in2(N__26929),
            .in3(N__26917),
            .lcout(\current_shift_inst.control_input_1_axb_1 ),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_10_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_10_22_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__31621),
            .in2(N__26914),
            .in3(N__26905),
            .lcout(\current_shift_inst.control_input_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_7 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_10_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_10_22_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__26902),
            .in2(N__31375),
            .in3(N__26893),
            .lcout(\current_shift_inst.control_input_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_8 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_10_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_10_22_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__26890),
            .in2(N__26884),
            .in3(N__26875),
            .lcout(\current_shift_inst.control_input_1_axb_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_9 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_10_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_10_22_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__27817),
            .in2(N__26872),
            .in3(N__26860),
            .lcout(\current_shift_inst.control_input_1_axb_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_10 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_10_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_10_22_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(N__31588),
            .in2(N__27112),
            .in3(N__27103),
            .lcout(\current_shift_inst.control_input_1_axb_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_11 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_10_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_10_22_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(N__31555),
            .in2(N__27100),
            .in3(N__27088),
            .lcout(\current_shift_inst.control_input_1_axb_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_12 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_10_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_10_22_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(N__27085),
            .in2(N__27079),
            .in3(N__27067),
            .lcout(\current_shift_inst.control_input_1_axb_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_13 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_10_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_10_23_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__31540),
            .in2(N__27064),
            .in3(N__27052),
            .lcout(\current_shift_inst.control_input_1_axb_9 ),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_10_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_10_23_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(N__27049),
            .in2(N__27037),
            .in3(N__27025),
            .lcout(\current_shift_inst.control_input_1_axb_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_15 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_10_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_10_23_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__31510),
            .in2(N__31483),
            .in3(N__27022),
            .lcout(\current_shift_inst.control_input_1_axb_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_16 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_10_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_10_23_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(N__27019),
            .in2(N__34189),
            .in3(N__27010),
            .lcout(\current_shift_inst.control_input_1_axb_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_17 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_10_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_10_23_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__27007),
            .in2(N__26998),
            .in3(N__26983),
            .lcout(\current_shift_inst.control_input_1_axb_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_18 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_10_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_10_23_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(N__31525),
            .in2(N__31609),
            .in3(N__26980),
            .lcout(\current_shift_inst.control_input_1_axb_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_19 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_10_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_10_23_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_10_23_6  (
            .in0(_gnd_net_),
            .in1(N__27208),
            .in2(N__27199),
            .in3(N__27187),
            .lcout(\current_shift_inst.control_input_1_axb_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_20 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_10_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_10_23_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(N__27184),
            .in2(N__27178),
            .in3(N__27166),
            .lcout(\current_shift_inst.control_input_1_axb_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_21 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_10_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_10_24_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_10_24_0  (
            .in0(_gnd_net_),
            .in1(N__27163),
            .in2(N__27148),
            .in3(N__27130),
            .lcout(\current_shift_inst.control_input_1_axb_17 ),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_10_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_10_24_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_10_24_1  (
            .in0(_gnd_net_),
            .in1(N__28837),
            .in2(N__31573),
            .in3(N__27127),
            .lcout(\current_shift_inst.control_input_1_axb_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_23 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_10_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_10_24_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_10_24_2  (
            .in0(_gnd_net_),
            .in1(N__31666),
            .in2(N__28831),
            .in3(N__27124),
            .lcout(\current_shift_inst.control_input_1_axb_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_24 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_10_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_10_24_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_10_24_3  (
            .in0(_gnd_net_),
            .in1(N__31651),
            .in2(N__28822),
            .in3(N__27121),
            .lcout(\current_shift_inst.control_input_1_axb_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_25 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_10_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_10_24_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(N__31807),
            .in2(N__31720),
            .in3(N__27118),
            .lcout(\current_shift_inst.control_input_1_axb_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_26 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_10_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_10_24_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_10_24_5  (
            .in0(_gnd_net_),
            .in1(N__31636),
            .in2(N__31699),
            .in3(N__27115),
            .lcout(\current_shift_inst.control_input_1_axb_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_27 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_10_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_10_24_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_10_24_6  (
            .in0(_gnd_net_),
            .in1(N__31681),
            .in2(N__27832),
            .in3(N__27355),
            .lcout(\current_shift_inst.control_input_1_axb_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_28 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_10_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_10_24_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_10_24_7  (
            .in0(_gnd_net_),
            .in1(N__28843),
            .in2(N__28866),
            .in3(N__27352),
            .lcout(\current_shift_inst.control_input_1_axb_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_29 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_25_LC_10_25_0 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_25_LC_10_25_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_25_LC_10_25_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.control_input_25_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(N__31495),
            .in2(N__28879),
            .in3(N__27349),
            .lcout(\current_shift_inst.control_inputZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48704),
            .ce(N__28963),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_11_3_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_11_3_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_11_3_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_11_3_1 (
            .in0(N__27289),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48853),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_11_5_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_11_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__27272),
            .in2(_gnd_net_),
            .in3(N__30174),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_336_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_11_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_11_6_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_27_LC_11_6_1  (
            .in0(N__27244),
            .in1(N__33586),
            .in2(_gnd_net_),
            .in3(N__30467),
            .lcout(measured_delay_hc_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48833),
            .ce(),
            .sr(N__48102));
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_11_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_11_6_2 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_28_LC_11_6_2  (
            .in0(N__30468),
            .in1(_gnd_net_),
            .in2(N__33627),
            .in3(N__27232),
            .lcout(measured_delay_hc_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48833),
            .ce(),
            .sr(N__48102));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_11_7_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_11_7_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_11_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_11_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27220),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48823),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_11_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_11_7_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_11_7_1  (
            .in0(N__29348),
            .in1(N__29372),
            .in2(N__30519),
            .in3(N__29268),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_11_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_11_7_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__29475),
            .in2(_gnd_net_),
            .in3(N__29511),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_10_LC_11_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_10_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_10_LC_11_7_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_10_LC_11_7_3  (
            .in0(N__27403),
            .in1(N__27394),
            .in2(N__27397),
            .in3(N__27385),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_11_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_11_7_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_11_7_4  (
            .in0(N__29616),
            .in1(N__30356),
            .in2(N__29208),
            .in3(N__29405),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_11_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_11_7_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__29637),
            .in2(_gnd_net_),
            .in3(N__29664),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_4_LC_11_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_4_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_4_LC_11_7_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_4_LC_11_7_6  (
            .in0(N__27475),
            .in1(N__29171),
            .in2(N__27388),
            .in3(N__29144),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP8VO1_20_LC_11_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP8VO1_20_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP8VO1_20_LC_11_8_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP8VO1_20_LC_11_8_0  (
            .in0(N__29569),
            .in1(N__27468),
            .in2(N__29557),
            .in3(N__29587),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_11_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_11_8_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__29553),
            .in2(_gnd_net_),
            .in3(N__29568),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1LC84_14_LC_11_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1LC84_14_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1LC84_14_LC_11_8_2 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1LC84_14_LC_11_8_2  (
            .in0(N__30515),
            .in1(N__27370),
            .in2(N__27493),
            .in3(N__29267),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_11_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_11_8_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_11_8_3  (
            .in0(N__27364),
            .in1(N__27457),
            .in2(N__27358),
            .in3(N__27499),
            .lcout(\delay_measurement_inst.un1_elapsed_time_hc ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINN412_20_LC_11_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINN412_20_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINN412_20_LC_11_8_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINN412_20_LC_11_8_4  (
            .in0(N__29586),
            .in1(N__27469),
            .in2(N__29720),
            .in3(N__27505),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_11_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_11_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_11_8_5  (
            .in0(N__29636),
            .in1(N__29663),
            .in2(N__29615),
            .in3(N__29990),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_11_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_11_8_6 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__30511),
            .in2(N__27484),
            .in3(N__29266),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_11_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_11_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_11_8_7  (
            .in0(N__29438),
            .in1(N__29100),
            .in2(N__29306),
            .in3(N__29991),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_11_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_11_9_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_11_9_3  (
            .in0(N__29788),
            .in1(N__29797),
            .in2(N__29779),
            .in3(N__29539),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_11_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_11_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_11_10_5  (
            .in0(N__29749),
            .in1(N__29758),
            .in2(N__29740),
            .in3(N__29767),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_11_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_11_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_11_11_0  (
            .in0(N__27433),
            .in1(N__27427),
            .in2(N__27421),
            .in3(N__27799),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_11_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_11_11_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__33159),
            .in2(N__27412),
            .in3(N__33125),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlt31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_11_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_11_4  (
            .in0(N__35314),
            .in1(N__35985),
            .in2(_gnd_net_),
            .in3(N__35255),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_11_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_11_11_5 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_11_11_5  (
            .in0(N__36087),
            .in1(N__35379),
            .in2(N__27802),
            .in3(N__35704),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_11_12_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_11_12_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_11_12_1  (
            .in0(N__27791),
            .in1(N__27773),
            .in2(_gnd_net_),
            .in3(N__27756),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto9_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_11_12_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_11_12_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_11_12_2  (
            .in0(N__27739),
            .in1(N__27721),
            .in2(N__27703),
            .in3(N__27568),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_11_12_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_11_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__27659),
            .in2(_gnd_net_),
            .in3(N__27641),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_11_12_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_11_12_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_11_12_4  (
            .in0(N__27624),
            .in1(N__27606),
            .in2(N__27589),
            .in3(N__27585),
            .lcout(\pwm_generator_inst.un1_counterlt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_14_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_14_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_11_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27562),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48761),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.running_LC_11_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_LC_11_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.running_LC_11_15_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_phase.running_LC_11_15_2  (
            .in0(N__31792),
            .in1(N__31831),
            .in2(_gnd_net_),
            .in3(N__31762),
            .lcout(\current_shift_inst.timer_phase.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48755),
            .ce(),
            .sr(N__48159));
    defparam \phase_controller_inst1.start_timer_tr_LC_11_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_11_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_11_15_3 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_11_15_3  (
            .in0(N__27528),
            .in1(N__27853),
            .in2(N__32684),
            .in3(N__27553),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48755),
            .ce(),
            .sr(N__48159));
    defparam \phase_controller_inst1.state_4_LC_11_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_11_15_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_11_15_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__30984),
            .in2(_gnd_net_),
            .in3(N__27527),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48755),
            .ce(),
            .sr(N__48159));
    defparam \current_shift_inst.S1_rise_LC_11_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.S1_rise_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_rise_LC_11_16_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \current_shift_inst.S1_rise_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__27838),
            .in2(_gnd_net_),
            .in3(N__27846),
            .lcout(\current_shift_inst.S1_riseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48749),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync0_LC_11_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync0_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync0_LC_11_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S1_sync0_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30030),
            .lcout(\current_shift_inst.S1_syncZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48749),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync1_LC_11_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync1_LC_11_16_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync1_LC_11_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S1_sync1_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27859),
            .lcout(\current_shift_inst.S1_syncZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48749),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__39666),
            .in2(_gnd_net_),
            .in3(N__29903),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync_prev_LC_11_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync_prev_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync_prev_LC_11_16_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.S1_sync_prev_LC_11_16_7  (
            .in0(N__27847),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.S1_sync_prevZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48749),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_0_LC_11_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_11_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_11_17_0 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst1.state_0_LC_11_17_0  (
            .in0(N__29904),
            .in1(N__39635),
            .in2(N__39683),
            .in3(N__39545),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48743),
            .ce(),
            .sr(N__48181));
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_11_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_11_18_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_18_LC_11_18_3  (
            .in0(N__49126),
            .in1(N__47179),
            .in2(_gnd_net_),
            .in3(N__46240),
            .lcout(measured_delay_tr_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48736),
            .ce(N__46354),
            .sr(N__48189));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_11_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_11_19_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_11_19_0  (
            .in0(N__41336),
            .in1(N__34960),
            .in2(N__35002),
            .in3(N__41248),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_11_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_11_19_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_11_19_1  (
            .in0(N__40502),
            .in1(N__34355),
            .in2(N__34402),
            .in3(N__40412),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_11_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_11_19_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_11_19_6  (
            .in0(N__39814),
            .in1(N__39763),
            .in2(N__39736),
            .in3(N__45253),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_11_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_11_19_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_11_19_7  (
            .in0(N__45153),
            .in1(N__45057),
            .in2(_gnd_net_),
            .in3(N__44994),
            .lcout(\phase_controller_inst1.stoper_tr.N_20_li ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_0_LC_11_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_0_LC_11_20_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_0_LC_11_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_0_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__28189),
            .in2(N__30094),
            .in3(N__30093),
            .lcout(\current_shift_inst.control_inputZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\current_shift_inst.control_input_1_cry_0 ),
            .clk(N__48723),
            .ce(N__28950),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_LC_11_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_1_LC_11_20_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_1_LC_11_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_1_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__28156),
            .in2(_gnd_net_),
            .in3(N__28117),
            .lcout(\current_shift_inst.control_inputZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_0 ),
            .carryout(\current_shift_inst.control_input_1_cry_1 ),
            .clk(N__48723),
            .ce(N__28950),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_2_LC_11_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_2_LC_11_20_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_2_LC_11_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_2_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__28114),
            .in2(_gnd_net_),
            .in3(N__28072),
            .lcout(\current_shift_inst.control_inputZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_1 ),
            .carryout(\current_shift_inst.control_input_1_cry_2 ),
            .clk(N__48723),
            .ce(N__28950),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_3_LC_11_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_3_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_3_LC_11_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_3_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__28069),
            .in2(_gnd_net_),
            .in3(N__28027),
            .lcout(\current_shift_inst.control_inputZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_2 ),
            .carryout(\current_shift_inst.control_input_1_cry_3 ),
            .clk(N__48723),
            .ce(N__28950),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_4_LC_11_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_4_LC_11_20_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_4_LC_11_20_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_4_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28024),
            .in3(N__27982),
            .lcout(\current_shift_inst.control_inputZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_3 ),
            .carryout(\current_shift_inst.control_input_1_cry_4 ),
            .clk(N__48723),
            .ce(N__28950),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_5_LC_11_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_5_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_5_LC_11_20_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_5_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27979),
            .in3(N__27940),
            .lcout(\current_shift_inst.control_inputZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_4 ),
            .carryout(\current_shift_inst.control_input_1_cry_5 ),
            .clk(N__48723),
            .ce(N__28950),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_6_LC_11_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_6_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_6_LC_11_20_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_6_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28504),
            .in3(N__28465),
            .lcout(\current_shift_inst.control_inputZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_5 ),
            .carryout(\current_shift_inst.control_input_1_cry_6 ),
            .clk(N__48723),
            .ce(N__28950),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_7_LC_11_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_7_LC_11_20_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_7_LC_11_20_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_7_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28462),
            .in3(N__28420),
            .lcout(\current_shift_inst.control_inputZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_6 ),
            .carryout(\current_shift_inst.control_input_1_cry_7 ),
            .clk(N__48723),
            .ce(N__28950),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_8_LC_11_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_8_LC_11_21_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_8_LC_11_21_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_8_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28417),
            .in3(N__28381),
            .lcout(\current_shift_inst.control_inputZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\current_shift_inst.control_input_1_cry_8 ),
            .clk(N__48716),
            .ce(N__28964),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_9_LC_11_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_9_LC_11_21_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_9_LC_11_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_9_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__28378),
            .in2(_gnd_net_),
            .in3(N__28345),
            .lcout(\current_shift_inst.control_inputZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_8 ),
            .carryout(\current_shift_inst.control_input_1_cry_9 ),
            .clk(N__48716),
            .ce(N__28964),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_10_LC_11_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_10_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_10_LC_11_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_10_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(N__28342),
            .in2(_gnd_net_),
            .in3(N__28306),
            .lcout(\current_shift_inst.control_inputZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_9 ),
            .carryout(\current_shift_inst.control_input_1_cry_10 ),
            .clk(N__48716),
            .ce(N__28964),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_11_LC_11_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_11_LC_11_21_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_11_LC_11_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_11_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__28303),
            .in2(_gnd_net_),
            .in3(N__28267),
            .lcout(\current_shift_inst.control_inputZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_10 ),
            .carryout(\current_shift_inst.control_input_1_cry_11 ),
            .clk(N__48716),
            .ce(N__28964),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_12_LC_11_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_12_LC_11_21_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_12_LC_11_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_12_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__28264),
            .in2(_gnd_net_),
            .in3(N__28234),
            .lcout(\current_shift_inst.control_inputZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_11 ),
            .carryout(\current_shift_inst.control_input_1_cry_12 ),
            .clk(N__48716),
            .ce(N__28964),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_13_LC_11_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_13_LC_11_21_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_13_LC_11_21_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_13_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28231),
            .in3(N__28192),
            .lcout(\current_shift_inst.control_inputZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_12 ),
            .carryout(\current_shift_inst.control_input_1_cry_13 ),
            .clk(N__48716),
            .ce(N__28964),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_14_LC_11_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_14_LC_11_21_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_14_LC_11_21_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_14_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28813),
            .in3(N__28777),
            .lcout(\current_shift_inst.control_inputZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_13 ),
            .carryout(\current_shift_inst.control_input_1_cry_14 ),
            .clk(N__48716),
            .ce(N__28964),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_15_LC_11_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_15_LC_11_21_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_15_LC_11_21_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_15_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28774),
            .in3(N__28732),
            .lcout(\current_shift_inst.control_inputZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_14 ),
            .carryout(\current_shift_inst.control_input_1_cry_15 ),
            .clk(N__48716),
            .ce(N__28964),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_16_LC_11_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_16_LC_11_22_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_16_LC_11_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_16_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__28729),
            .in2(_gnd_net_),
            .in3(N__28696),
            .lcout(\current_shift_inst.control_inputZ0Z_16 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\current_shift_inst.control_input_1_cry_16 ),
            .clk(N__48710),
            .ce(N__28965),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_17_LC_11_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_17_LC_11_22_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_17_LC_11_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_17_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__28693),
            .in2(_gnd_net_),
            .in3(N__28660),
            .lcout(\current_shift_inst.control_inputZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_16 ),
            .carryout(\current_shift_inst.control_input_1_cry_17 ),
            .clk(N__48710),
            .ce(N__28965),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_18_LC_11_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_18_LC_11_22_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_18_LC_11_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_18_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__28657),
            .in2(_gnd_net_),
            .in3(N__28624),
            .lcout(\current_shift_inst.control_inputZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_17 ),
            .carryout(\current_shift_inst.control_input_1_cry_18 ),
            .clk(N__48710),
            .ce(N__28965),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_19_LC_11_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_19_LC_11_22_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_19_LC_11_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_19_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__28621),
            .in2(_gnd_net_),
            .in3(N__28588),
            .lcout(\current_shift_inst.control_inputZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_18 ),
            .carryout(\current_shift_inst.control_input_1_cry_19 ),
            .clk(N__48710),
            .ce(N__28965),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_20_LC_11_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_20_LC_11_22_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_20_LC_11_22_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_20_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28585),
            .in3(N__28552),
            .lcout(\current_shift_inst.control_inputZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_19 ),
            .carryout(\current_shift_inst.control_input_1_cry_20 ),
            .clk(N__48710),
            .ce(N__28965),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_21_LC_11_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_21_LC_11_22_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_21_LC_11_22_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_21_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28549),
            .in3(N__28507),
            .lcout(\current_shift_inst.control_inputZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_20 ),
            .carryout(\current_shift_inst.control_input_1_cry_21 ),
            .clk(N__48710),
            .ce(N__28965),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_22_LC_11_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_22_LC_11_22_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_22_LC_11_22_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_22_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29086),
            .in3(N__29047),
            .lcout(\current_shift_inst.control_inputZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_21 ),
            .carryout(\current_shift_inst.control_input_1_cry_22 ),
            .clk(N__48710),
            .ce(N__28965),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_23_LC_11_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_23_LC_11_22_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_23_LC_11_22_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_23_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29044),
            .in3(N__29005),
            .lcout(\current_shift_inst.control_inputZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_22 ),
            .carryout(\current_shift_inst.control_input_1_cry_23 ),
            .clk(N__48710),
            .ce(N__28965),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_24_LC_11_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_24_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_24_LC_11_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_24_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__29002),
            .in2(_gnd_net_),
            .in3(N__28972),
            .lcout(\current_shift_inst.control_inputZ0Z_24 ),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\current_shift_inst.control_input_1_cry_24 ),
            .clk(N__48707),
            .ce(N__28969),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_11_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_11_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28882),
            .lcout(\current_shift_inst.control_input_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_11_24_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_11_24_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_11_24_0  (
            .in0(N__28867),
            .in1(N__41886),
            .in2(_gnd_net_),
            .in3(N__34927),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_11_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_11_24_1 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_11_24_1  (
            .in0(N__34558),
            .in1(N__41579),
            .in2(N__35131),
            .in3(N__41654),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_11_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_11_24_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_11_24_2  (
            .in0(N__41580),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35130),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_11_24_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_11_24_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_11_24_7  (
            .in0(_gnd_net_),
            .in1(N__41520),
            .in2(_gnd_net_),
            .in3(N__35095),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_25_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_25_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_25_0  (
            .in0(N__32686),
            .in1(N__32895),
            .in2(N__30199),
            .in3(N__32569),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48702),
            .ce(),
            .sr(N__48228));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_11_25_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_11_25_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_11_25_2  (
            .in0(N__32685),
            .in1(N__32894),
            .in2(_gnd_net_),
            .in3(N__32568),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_11_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_11_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_11_25_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_11_25_3  (
            .in0(N__39631),
            .in1(N__32406),
            .in2(N__29230),
            .in3(N__32368),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48702),
            .ce(),
            .sr(N__48228));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_12_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_12_6_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_12_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30337),
            .lcout(\delay_measurement_inst.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48822),
            .ce(N__29691),
            .sr(N__48095));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_12_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_12_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_12_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30316),
            .lcout(\delay_measurement_inst.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48822),
            .ce(N__29691),
            .sr(N__48095));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_12_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_12_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_12_7_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__30336),
            .in2(N__30294),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__48812),
            .ce(N__29692),
            .sr(N__48103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_12_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_12_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_12_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__30315),
            .in2(N__30270),
            .in3(N__29152),
            .lcout(\delay_measurement_inst.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__48812),
            .ce(N__29692),
            .sr(N__48103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_12_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_12_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_12_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(N__30245),
            .in2(N__30295),
            .in3(N__29125),
            .lcout(\delay_measurement_inst.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__48812),
            .ce(N__29692),
            .sr(N__48103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_12_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_12_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_12_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__30227),
            .in2(N__30271),
            .in3(N__29089),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__48812),
            .ce(N__29692),
            .sr(N__48103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_12_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_12_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_12_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__30246),
            .in2(N__30726),
            .in3(N__29500),
            .lcout(\delay_measurement_inst.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__48812),
            .ce(N__29692),
            .sr(N__48103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_12_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_12_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_12_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__30228),
            .in2(N__30702),
            .in3(N__29464),
            .lcout(\delay_measurement_inst.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__48812),
            .ce(N__29692),
            .sr(N__48103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_12_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_12_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_12_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(N__30679),
            .in2(N__30727),
            .in3(N__29422),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__48812),
            .ce(N__29692),
            .sr(N__48103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_12_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_12_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_12_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(N__30655),
            .in2(N__30703),
            .in3(N__29386),
            .lcout(\delay_measurement_inst.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__48812),
            .ce(N__29692),
            .sr(N__48103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_12_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_12_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_12_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__30678),
            .in2(N__30630),
            .in3(N__29356),
            .lcout(\delay_measurement_inst.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__48806),
            .ce(N__29693),
            .sr(N__48109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_12_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_12_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_12_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__30654),
            .in2(N__30606),
            .in3(N__29314),
            .lcout(\delay_measurement_inst.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__48806),
            .ce(N__29693),
            .sr(N__48109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_12_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_12_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__30581),
            .in2(N__30631),
            .in3(N__29281),
            .lcout(\delay_measurement_inst.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__48806),
            .ce(N__29693),
            .sr(N__48109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_12_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_12_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__30563),
            .in2(N__30607),
            .in3(N__29278),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__48806),
            .ce(N__29693),
            .sr(N__48109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_12_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_12_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__30582),
            .in2(N__30546),
            .in3(N__29233),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__48806),
            .ce(N__29693),
            .sr(N__48109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_12_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_12_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_12_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__30564),
            .in2(N__30906),
            .in3(N__29674),
            .lcout(\delay_measurement_inst.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__48806),
            .ce(N__29693),
            .sr(N__48109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_12_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_12_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_12_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(N__30883),
            .in2(N__30547),
            .in3(N__29647),
            .lcout(\delay_measurement_inst.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__48806),
            .ce(N__29693),
            .sr(N__48109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_12_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_12_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_12_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__30859),
            .in2(N__30907),
            .in3(N__29620),
            .lcout(\delay_measurement_inst.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__48806),
            .ce(N__29693),
            .sr(N__48109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_12_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_12_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_12_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__30882),
            .in2(N__30834),
            .in3(N__29590),
            .lcout(\delay_measurement_inst.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__48795),
            .ce(N__29694),
            .sr(N__48118));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_12_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_12_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_12_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__30858),
            .in2(N__30810),
            .in3(N__29572),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__48795),
            .ce(N__29694),
            .sr(N__48118));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_12_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_12_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_12_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__30785),
            .in2(N__30835),
            .in3(N__29560),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__48795),
            .ce(N__29694),
            .sr(N__48118));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_12_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_12_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__30767),
            .in2(N__30811),
            .in3(N__29542),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__48795),
            .ce(N__29694),
            .sr(N__48118));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_12_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_12_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_12_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__30786),
            .in2(N__30750),
            .in3(N__29533),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__48795),
            .ce(N__29694),
            .sr(N__48118));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_12_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_12_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_12_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__30768),
            .in2(N__31356),
            .in3(N__29791),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__48795),
            .ce(N__29694),
            .sr(N__48118));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_12_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_12_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_12_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__31333),
            .in2(N__30751),
            .in3(N__29782),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__48795),
            .ce(N__29694),
            .sr(N__48118));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_12_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_12_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_12_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__31309),
            .in2(N__31357),
            .in3(N__29770),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__48795),
            .ce(N__29694),
            .sr(N__48118));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_12_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_12_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_12_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__31332),
            .in2(N__31284),
            .in3(N__29761),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__48787),
            .ce(N__29695),
            .sr(N__48125));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_12_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_12_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__31308),
            .in2(N__31260),
            .in3(N__29752),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__48787),
            .ce(N__29695),
            .sr(N__48125));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_12_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_12_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__31236),
            .in2(N__31285),
            .in3(N__29743),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__48787),
            .ce(N__29695),
            .sr(N__48125));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_12_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_12_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__31095),
            .in2(N__31261),
            .in3(N__29731),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__48787),
            .ce(N__29695),
            .sr(N__48125));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_12_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_12_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_12_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29728),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48787),
            .ce(N__29695),
            .sr(N__48125));
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_12_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_12_11_0 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_16_LC_12_11_0  (
            .in0(N__33574),
            .in1(N__29995),
            .in2(N__33306),
            .in3(N__30486),
            .lcout(measured_delay_hc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48779),
            .ce(),
            .sr(N__48129));
    defparam \phase_controller_slave.state_4_LC_12_12_5 .C_ON=1'b0;
    defparam \phase_controller_slave.state_4_LC_12_12_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.state_4_LC_12_12_5 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_slave.state_4_LC_12_12_5  (
            .in0(N__31008),
            .in1(N__45714),
            .in2(_gnd_net_),
            .in3(N__45923),
            .lcout(\phase_controller_slave.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48770),
            .ce(),
            .sr(N__48134));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_13_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_13_1  (
            .in0(N__29880),
            .in1(N__33780),
            .in2(_gnd_net_),
            .in3(N__29833),
            .lcout(\current_shift_inst.timer_s1.N_191_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.T01_er_LC_12_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_er_LC_12_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_er_LC_12_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.T01_er_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29946),
            .lcout(shift_flag_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48754),
            .ce(N__39520),
            .sr(N__48147));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_12_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_12_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_12_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42568),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48748),
            .ce(N__39875),
            .sr(N__48153));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42535),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48748),
            .ce(N__39875),
            .sr(N__48153));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39849),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48748),
            .ce(N__39875),
            .sr(N__48153));
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_12_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_12_16_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_7_LC_12_16_5  (
            .in0(N__46154),
            .in1(N__46978),
            .in2(N__38998),
            .in3(N__43879),
            .lcout(measured_delay_tr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48742),
            .ce(),
            .sr(N__48160));
    defparam \phase_controller_inst1.state_1_LC_12_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_12_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_12_16_7 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_1_LC_12_16_7  (
            .in0(N__29977),
            .in1(N__39673),
            .in2(N__29947),
            .in3(N__29905),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48742),
            .ce(),
            .sr(N__48160));
    defparam \current_shift_inst.timer_s1.running_LC_12_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_12_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_12_17_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_12_17_2  (
            .in0(N__29881),
            .in1(N__33766),
            .in2(_gnd_net_),
            .in3(N__29832),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48735),
            .ce(),
            .sr(N__48170));
    defparam \phase_controller_inst1.S1_LC_12_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_12_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_12_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39597),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48735),
            .ce(),
            .sr(N__48170));
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_12_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_12_17_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_12_17_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_8_LC_12_17_5  (
            .in0(N__46155),
            .in1(N__46924),
            .in2(N__39038),
            .in3(N__43878),
            .lcout(measured_delay_tr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48735),
            .ce(),
            .sr(N__48170));
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_12_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_12_18_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_12_18_2 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_17_LC_12_18_2  (
            .in0(N__49124),
            .in1(N__47233),
            .in2(_gnd_net_),
            .in3(N__46238),
            .lcout(measured_delay_tr_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48730),
            .ce(N__46350),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_12_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_12_18_5 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_12_18_5 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_1_LC_12_18_5  (
            .in0(N__46531),
            .in1(N__48894),
            .in2(N__46167),
            .in3(N__46447),
            .lcout(measured_delay_tr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48730),
            .ce(N__46350),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_12_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_12_18_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_12_18_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_19_LC_12_18_7  (
            .in0(N__46239),
            .in1(N__49125),
            .in2(_gnd_net_),
            .in3(N__47122),
            .lcout(measured_delay_tr_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48730),
            .ce(N__46350),
            .sr(N__48182));
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_12_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_12_19_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_16_LC_12_19_3  (
            .in0(N__49115),
            .in1(N__47293),
            .in2(_gnd_net_),
            .in3(N__46250),
            .lcout(measured_delay_tr_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48722),
            .ce(N__46345),
            .sr(N__48190));
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_12_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_12_19_4 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_12_19_4 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_3_LC_12_19_4  (
            .in0(N__46087),
            .in1(N__46527),
            .in2(N__46166),
            .in3(N__46446),
            .lcout(measured_delay_tr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48722),
            .ce(N__46345),
            .sr(N__48190));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_20_0 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_20_0  (
            .in0(N__32897),
            .in1(N__32690),
            .in2(N__32570),
            .in3(N__30124),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48715),
            .ce(),
            .sr(N__48197));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_20_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_20_1  (
            .in0(N__32526),
            .in1(N__32898),
            .in2(N__32732),
            .in3(N__30112),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48715),
            .ce(),
            .sr(N__48197));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_12_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_12_20_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_12_20_4  (
            .in0(N__30019),
            .in1(N__46569),
            .in2(N__38798),
            .in3(N__30004),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_14_LC_12_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_14_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_14_LC_12_20_6 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_14_LC_12_20_6  (
            .in0(N__46284),
            .in1(N__47427),
            .in2(N__36821),
            .in3(N__43876),
            .lcout(measured_delay_tr_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48715),
            .ce(),
            .sr(N__48197));
    defparam \delay_measurement_inst.delay_tr_reg_15_LC_12_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_15_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_15_LC_12_20_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_15_LC_12_20_7  (
            .in0(N__43877),
            .in1(N__46285),
            .in2(N__38883),
            .in3(N__47365),
            .lcout(measured_delay_tr_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48715),
            .ce(),
            .sr(N__48197));
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_12_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_12_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_i_31_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34894),
            .lcout(\current_shift_inst.z_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_12_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_12_21_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_12_21_4  (
            .in0(N__39994),
            .in1(N__39931),
            .in2(N__33964),
            .in3(N__33914),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_12_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_12_22_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIC90O_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(N__31846),
            .in2(_gnd_net_),
            .in3(N__31760),
            .lcout(\current_shift_inst.timer_phase.N_188_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_12_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_12_23_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_12_23_4  (
            .in0(N__32349),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32402),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_12_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_12_23_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(N__32401),
            .in2(_gnd_net_),
            .in3(N__32348),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_12_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_12_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(N__30055),
            .in2(N__32317),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_24_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_12_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_12_24_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_12_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33055),
            .in3(N__30049),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_12_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_12_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_12_24_2  (
            .in0(_gnd_net_),
            .in1(N__30145),
            .in2(N__33031),
            .in3(N__30139),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_12_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_12_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_12_24_3  (
            .in0(_gnd_net_),
            .in1(N__33006),
            .in2(_gnd_net_),
            .in3(N__30136),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_12_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_12_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_12_24_4  (
            .in0(_gnd_net_),
            .in1(N__32985),
            .in2(_gnd_net_),
            .in3(N__30133),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_12_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_12_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_12_24_5  (
            .in0(_gnd_net_),
            .in1(N__32961),
            .in2(_gnd_net_),
            .in3(N__30130),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_12_24_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_12_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(N__32940),
            .in2(_gnd_net_),
            .in3(N__30127),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_12_24_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_12_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_12_24_7  (
            .in0(_gnd_net_),
            .in1(N__32044),
            .in2(_gnd_net_),
            .in3(N__30115),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_12_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_12_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_12_25_0  (
            .in0(_gnd_net_),
            .in1(N__32008),
            .in2(_gnd_net_),
            .in3(N__30103),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ),
            .ltout(),
            .carryin(bfn_12_25_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_12_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_12_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_12_25_1  (
            .in0(_gnd_net_),
            .in1(N__32421),
            .in2(_gnd_net_),
            .in3(N__30100),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_12_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_12_25_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_12_25_2  (
            .in0(_gnd_net_),
            .in1(N__32286),
            .in2(_gnd_net_),
            .in3(N__30097),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_12_25_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_12_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_12_25_3  (
            .in0(_gnd_net_),
            .in1(N__32265),
            .in2(_gnd_net_),
            .in3(N__30211),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_12_25_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_12_25_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_12_25_4  (
            .in0(_gnd_net_),
            .in1(N__32244),
            .in2(_gnd_net_),
            .in3(N__30208),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_12_25_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_12_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_12_25_5  (
            .in0(_gnd_net_),
            .in1(N__32223),
            .in2(_gnd_net_),
            .in3(N__30205),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_12_25_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_12_25_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_12_25_6  (
            .in0(_gnd_net_),
            .in1(N__32202),
            .in2(_gnd_net_),
            .in3(N__30202),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_12_25_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_12_25_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_12_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32145),
            .in3(N__30190),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_12_26_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_12_26_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_12_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_12_26_0  (
            .in0(_gnd_net_),
            .in1(N__32442),
            .in2(_gnd_net_),
            .in3(N__30187),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ),
            .ltout(),
            .carryin(bfn_12_26_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_12_26_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_12_26_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_12_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_12_26_1  (
            .in0(_gnd_net_),
            .in1(N__32181),
            .in2(_gnd_net_),
            .in3(N__30184),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_12_26_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_12_26_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_12_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_12_26_2  (
            .in0(_gnd_net_),
            .in1(N__33075),
            .in2(_gnd_net_),
            .in3(N__30181),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_5_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30178),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_13_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_13_6_3 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_14_LC_13_6_3  (
            .in0(N__30523),
            .in1(N__33628),
            .in2(N__33360),
            .in3(N__30484),
            .lcout(measured_delay_hc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48834),
            .ce(),
            .sr(N__48091));
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_13_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_13_6_7 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_13_6_7 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_3_LC_13_6_7  (
            .in0(N__36063),
            .in1(N__30485),
            .in2(N__33648),
            .in3(N__30357),
            .lcout(measured_delay_hc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48834),
            .ce(),
            .sr(N__48091));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_13_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_13_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_13_7_0  (
            .in0(N__31193),
            .in1(N__30335),
            .in2(_gnd_net_),
            .in3(N__30319),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__48824),
            .ce(N__31072),
            .sr(N__48096));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_13_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_13_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_13_7_1  (
            .in0(N__31205),
            .in1(N__30314),
            .in2(_gnd_net_),
            .in3(N__30298),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__48824),
            .ce(N__31072),
            .sr(N__48096));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_13_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_13_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_13_7_2  (
            .in0(N__31194),
            .in1(N__30293),
            .in2(_gnd_net_),
            .in3(N__30274),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__48824),
            .ce(N__31072),
            .sr(N__48096));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_13_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_13_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_13_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_13_7_3  (
            .in0(N__31206),
            .in1(N__30269),
            .in2(_gnd_net_),
            .in3(N__30250),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__48824),
            .ce(N__31072),
            .sr(N__48096));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_13_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_13_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_13_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_13_7_4  (
            .in0(N__31195),
            .in1(N__30247),
            .in2(_gnd_net_),
            .in3(N__30232),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__48824),
            .ce(N__31072),
            .sr(N__48096));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_13_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_13_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_13_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_13_7_5  (
            .in0(N__31207),
            .in1(N__30229),
            .in2(_gnd_net_),
            .in3(N__30214),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__48824),
            .ce(N__31072),
            .sr(N__48096));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_13_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_13_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_13_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_13_7_6  (
            .in0(N__31196),
            .in1(N__30725),
            .in2(_gnd_net_),
            .in3(N__30706),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__48824),
            .ce(N__31072),
            .sr(N__48096));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_13_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_13_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_13_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_13_7_7  (
            .in0(N__31208),
            .in1(N__30701),
            .in2(_gnd_net_),
            .in3(N__30682),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__48824),
            .ce(N__31072),
            .sr(N__48096));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_13_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_13_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_13_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_13_8_0  (
            .in0(N__31216),
            .in1(N__30677),
            .in2(_gnd_net_),
            .in3(N__30658),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__48814),
            .ce(N__31082),
            .sr(N__48104));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_13_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_13_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_13_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_13_8_1  (
            .in0(N__31200),
            .in1(N__30653),
            .in2(_gnd_net_),
            .in3(N__30634),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__48814),
            .ce(N__31082),
            .sr(N__48104));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_13_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_13_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_13_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_13_8_2  (
            .in0(N__31213),
            .in1(N__30629),
            .in2(_gnd_net_),
            .in3(N__30610),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__48814),
            .ce(N__31082),
            .sr(N__48104));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_13_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_13_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_13_8_3  (
            .in0(N__31197),
            .in1(N__30605),
            .in2(_gnd_net_),
            .in3(N__30586),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__48814),
            .ce(N__31082),
            .sr(N__48104));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_13_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_13_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_13_8_4  (
            .in0(N__31214),
            .in1(N__30583),
            .in2(_gnd_net_),
            .in3(N__30568),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__48814),
            .ce(N__31082),
            .sr(N__48104));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_13_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_13_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_13_8_5  (
            .in0(N__31198),
            .in1(N__30565),
            .in2(_gnd_net_),
            .in3(N__30550),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__48814),
            .ce(N__31082),
            .sr(N__48104));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_13_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_13_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_13_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_13_8_6  (
            .in0(N__31215),
            .in1(N__30545),
            .in2(_gnd_net_),
            .in3(N__30526),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__48814),
            .ce(N__31082),
            .sr(N__48104));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_13_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_13_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_13_8_7  (
            .in0(N__31199),
            .in1(N__30905),
            .in2(_gnd_net_),
            .in3(N__30886),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__48814),
            .ce(N__31082),
            .sr(N__48104));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_13_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_13_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_13_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_13_9_0  (
            .in0(N__31201),
            .in1(N__30881),
            .in2(_gnd_net_),
            .in3(N__30862),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__48807),
            .ce(N__31083),
            .sr(N__48110));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_13_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_13_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_13_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_13_9_1  (
            .in0(N__31217),
            .in1(N__30857),
            .in2(_gnd_net_),
            .in3(N__30838),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__48807),
            .ce(N__31083),
            .sr(N__48110));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_13_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_13_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_13_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_13_9_2  (
            .in0(N__31202),
            .in1(N__30833),
            .in2(_gnd_net_),
            .in3(N__30814),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__48807),
            .ce(N__31083),
            .sr(N__48110));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_13_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_13_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_13_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_13_9_3  (
            .in0(N__31218),
            .in1(N__30809),
            .in2(_gnd_net_),
            .in3(N__30790),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__48807),
            .ce(N__31083),
            .sr(N__48110));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_13_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_13_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_13_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_13_9_4  (
            .in0(N__31203),
            .in1(N__30787),
            .in2(_gnd_net_),
            .in3(N__30772),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__48807),
            .ce(N__31083),
            .sr(N__48110));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_13_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_13_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_13_9_5  (
            .in0(N__31219),
            .in1(N__30769),
            .in2(_gnd_net_),
            .in3(N__30754),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__48807),
            .ce(N__31083),
            .sr(N__48110));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_13_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_13_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_13_9_6  (
            .in0(N__31204),
            .in1(N__30749),
            .in2(_gnd_net_),
            .in3(N__30730),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__48807),
            .ce(N__31083),
            .sr(N__48110));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_13_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_13_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_13_9_7  (
            .in0(N__31220),
            .in1(N__31355),
            .in2(_gnd_net_),
            .in3(N__31336),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__48807),
            .ce(N__31083),
            .sr(N__48110));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_13_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_13_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_13_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_13_10_0  (
            .in0(N__31209),
            .in1(N__31331),
            .in2(_gnd_net_),
            .in3(N__31312),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__48796),
            .ce(N__31084),
            .sr(N__48119));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_13_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_13_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_13_10_1  (
            .in0(N__31221),
            .in1(N__31307),
            .in2(_gnd_net_),
            .in3(N__31288),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__48796),
            .ce(N__31084),
            .sr(N__48119));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_13_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_13_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_13_10_2  (
            .in0(N__31210),
            .in1(N__31283),
            .in2(_gnd_net_),
            .in3(N__31264),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__48796),
            .ce(N__31084),
            .sr(N__48119));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_13_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_13_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_13_10_3  (
            .in0(N__31222),
            .in1(N__31259),
            .in2(_gnd_net_),
            .in3(N__31240),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__48796),
            .ce(N__31084),
            .sr(N__48119));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_13_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_13_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_13_10_4  (
            .in0(N__31211),
            .in1(N__31237),
            .in2(_gnd_net_),
            .in3(N__31225),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__48796),
            .ce(N__31084),
            .sr(N__48119));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_13_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_13_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_13_10_5  (
            .in0(N__31096),
            .in1(N__31212),
            .in2(_gnd_net_),
            .in3(N__31099),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48796),
            .ce(N__31084),
            .sr(N__48119));
    defparam \phase_controller_slave.state_RNO_0_3_LC_13_12_6 .C_ON=1'b0;
    defparam \phase_controller_slave.state_RNO_0_3_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.state_RNO_0_3_LC_13_12_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_slave.state_RNO_0_3_LC_13_12_6  (
            .in0(N__30992),
            .in1(N__45713),
            .in2(_gnd_net_),
            .in3(N__45922),
            .lcout(\phase_controller_slave.N_213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39853),
            .lcout(\current_shift_inst.elapsed_time_ns_1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48772),
            .ce(N__39878),
            .sr(N__48135));
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_14_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_14_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_14_0  (
            .in0(N__42230),
            .in1(N__41978),
            .in2(N__42196),
            .in3(N__42600),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48762),
            .ce(N__31464),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_14_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_14_1 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_14_1  (
            .in0(N__42601),
            .in1(N__42191),
            .in2(N__42002),
            .in3(N__42231),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48762),
            .ce(N__31464),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_13_14_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_13_14_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_13_14_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_0_LC_13_14_2  (
            .in0(N__45433),
            .in1(N__45361),
            .in2(N__45655),
            .in3(N__45872),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48762),
            .ce(N__31464),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_13_14_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_13_14_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_13_14_3 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_1_LC_13_14_3  (
            .in0(N__45873),
            .in1(N__45643),
            .in2(N__45391),
            .in3(N__45434),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48762),
            .ce(N__31464),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_0_LC_13_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_0_LC_13_14_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_state_0_LC_13_14_5 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.tr_state_0_LC_13_14_5  (
            .in0(N__43987),
            .in1(N__44006),
            .in2(_gnd_net_),
            .in3(N__43951),
            .lcout(\delay_measurement_inst.tr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48762),
            .ce(N__31464),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31387),
            .lcout(\current_shift_inst.un4_control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_15_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(N__31381),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_13_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_13_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38743),
            .lcout(\current_shift_inst.un4_control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_13_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_13_16_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__40632),
            .in2(_gnd_net_),
            .in3(N__34468),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_13_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_13_16_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__40911),
            .in2(_gnd_net_),
            .in3(N__34708),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_13_16_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_13_16_2  (
            .in0(N__34339),
            .in1(N__40340),
            .in2(N__40423),
            .in3(N__34303),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_13_16_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__41662),
            .in2(_gnd_net_),
            .in3(N__34549),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_13_16_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_13_16_4  (
            .in0(N__40269),
            .in1(N__40341),
            .in2(N__34311),
            .in3(N__34258),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_13_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_13_16_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_13_16_5  (
            .in0(N__40193),
            .in1(N__34861),
            .in2(N__34233),
            .in3(N__41183),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_13_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_13_16_6  (
            .in0(N__40912),
            .in1(N__40838),
            .in2(N__34718),
            .in3(N__34669),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_13_16_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_13_16_7  (
            .in0(N__34819),
            .in1(N__41043),
            .in2(N__41116),
            .in3(N__34784),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_0_25_LC_13_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_13_17_0 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \current_shift_inst.control_input_RNO_0_25_LC_13_17_0  (
            .in0(N__41890),
            .in1(N__37408),
            .in2(N__41851),
            .in3(N__34913),
            .lcout(\current_shift_inst.un38_control_input_0_axb_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_13_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_13_17_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__41115),
            .in2(_gnd_net_),
            .in3(N__34833),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_13_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_13_17_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_13_17_2  (
            .in0(N__41469),
            .in1(N__41405),
            .in2(N__35056),
            .in3(N__35024),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_13_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_13_17_4 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIL91O_LC_13_17_4  (
            .in0(N__31791),
            .in1(N__31845),
            .in2(_gnd_net_),
            .in3(N__31761),
            .lcout(\current_shift_inst.timer_phase.N_192_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_13_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_13_17_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__41468),
            .in2(_gnd_net_),
            .in3(N__35050),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_13_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_13_17_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__41406),
            .in2(_gnd_net_),
            .in3(N__35023),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_13_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_13_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__41338),
            .in2(_gnd_net_),
            .in3(N__34985),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_RNIMR6L_0_LC_13_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_RNIMR6L_0_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.tr_state_RNIMR6L_0_LC_13_18_0 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \delay_measurement_inst.tr_state_RNIMR6L_0_LC_13_18_0  (
            .in0(N__43947),
            .in1(N__43981),
            .in2(_gnd_net_),
            .in3(N__44010),
            .lcout(\delay_measurement_inst.tr_state_RNIMR6LZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_13_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_13_18_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_13_18_1  (
            .in0(N__35117),
            .in1(N__41526),
            .in2(N__41590),
            .in3(N__35080),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_13_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_13_18_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_13_18_2  (
            .in0(N__41527),
            .in1(N__41470),
            .in2(N__35090),
            .in3(N__35054),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_13_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_13_18_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_13_18_4  (
            .in0(N__41407),
            .in1(N__41337),
            .in2(N__35029),
            .in3(N__34984),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_13_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_13_18_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_13_18_5  (
            .in0(N__34515),
            .in1(N__40628),
            .in2(N__40705),
            .in3(N__34479),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_13_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_13_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_13_19_0 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_13_19_0  (
            .in0(N__46382),
            .in1(N__39164),
            .in2(N__39122),
            .in3(N__39080),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48731),
            .ce(N__46641),
            .sr(N__48183));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_13_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_13_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_13_19_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_13_19_2  (
            .in0(N__39286),
            .in1(N__39165),
            .in2(N__39261),
            .in3(N__39079),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48731),
            .ce(N__46641),
            .sr(N__48183));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_13_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_13_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_13_19_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_13_19_3  (
            .in0(N__39081),
            .in1(N__39112),
            .in2(_gnd_net_),
            .in3(N__39166),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48731),
            .ce(N__46641),
            .sr(N__48183));
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_13_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_13_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIB31B_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31844),
            .lcout(\current_shift_inst.timer_phase.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_13_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_13_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_13_20_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_13_20_0  (
            .in0(N__45134),
            .in1(N__45053),
            .in2(N__38799),
            .in3(N__45006),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48724),
            .ce(N__46628),
            .sr(N__48191));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_13_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_13_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_13_20_1 .LUT_INIT=16'b0000111100000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_13_20_1  (
            .in0(N__45007),
            .in1(N__45135),
            .in2(N__45058),
            .in3(N__38962),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48724),
            .ce(N__46628),
            .sr(N__48191));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_13_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_13_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_13_20_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_13_20_2  (
            .in0(N__45136),
            .in1(N__39003),
            .in2(_gnd_net_),
            .in3(N__45004),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48724),
            .ce(N__46628),
            .sr(N__48191));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_13_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_13_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_13_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39832),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48724),
            .ce(N__46628),
            .sr(N__48191));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_13_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_13_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_13_20_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_13_20_4  (
            .in0(N__39037),
            .in1(N__45133),
            .in2(_gnd_net_),
            .in3(N__45005),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48724),
            .ce(N__46628),
            .sr(N__48191));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_13_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_13_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_13_20_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_13_20_5  (
            .in0(N__45132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38869),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48724),
            .ce(N__46628),
            .sr(N__48191));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_13_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_13_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_13_20_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_13_20_6  (
            .in0(N__38867),
            .in1(N__45131),
            .in2(_gnd_net_),
            .in3(N__36811),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48724),
            .ce(N__46628),
            .sr(N__48191));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_13_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_13_20_7 .LUT_INIT=16'b1111010011110101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_13_20_7  (
            .in0(N__36973),
            .in1(N__38868),
            .in2(N__39220),
            .in3(N__38833),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48724),
            .ce(N__46628),
            .sr(N__48191));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__31927),
            .in2(N__31942),
            .in3(N__32316),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__31909),
            .in2(N__31921),
            .in3(N__33054),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__31891),
            .in2(N__31903),
            .in3(N__33030),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(N__31885),
            .in2(N__46666),
            .in3(N__33007),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(N__31870),
            .in2(N__31879),
            .in3(N__32986),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__31852),
            .in2(N__31864),
            .in3(N__32965),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_21_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_21_6  (
            .in0(N__32941),
            .in1(N__32059),
            .in2(N__32068),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_21_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(N__32026),
            .in2(N__32053),
            .in3(N__32043),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__31990),
            .in2(N__32020),
            .in3(N__32007),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__31984),
            .in2(N__37057),
            .in3(N__32422),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__31978),
            .in2(N__37042),
            .in3(N__32287),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(N__31972),
            .in2(N__37027),
            .in3(N__32266),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(N__31966),
            .in2(N__36952),
            .in3(N__32245),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(N__31948),
            .in2(N__31960),
            .in3(N__32224),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_22_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(N__32152),
            .in2(N__32167),
            .in3(N__32203),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_22_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(N__32125),
            .in2(N__44035),
            .in3(N__32146),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_23_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__32119),
            .in2(N__32086),
            .in3(N__32443),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_23_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__32101),
            .in2(N__32113),
            .in3(N__32182),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_23_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__32095),
            .in2(N__32077),
            .in3(N__33076),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32089),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_13_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_13_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_13_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39786),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48708),
            .ce(N__46642),
            .sr(N__48211));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_13_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_13_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_13_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39740),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48708),
            .ce(N__46642),
            .sr(N__48211));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_13_24_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_13_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_13_24_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_13_24_0  (
            .in0(N__32899),
            .in1(N__32573),
            .in2(N__32777),
            .in3(N__32428),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48705),
            .ce(),
            .sr(N__48216));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_13_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_13_24_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_13_24_1  (
            .in0(N__32407),
            .in1(N__32315),
            .in2(_gnd_net_),
            .in3(N__32350),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_13_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_13_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_13_24_2 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_13_24_2  (
            .in0(N__32902),
            .in1(N__32576),
            .in2(N__32320),
            .in3(N__32757),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48705),
            .ce(),
            .sr(N__48216));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_13_24_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_13_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_13_24_3 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_13_24_3  (
            .in0(N__32293),
            .in1(N__32758),
            .in2(N__32594),
            .in3(N__32903),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48705),
            .ce(),
            .sr(N__48216));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_13_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_13_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_13_24_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_13_24_4  (
            .in0(N__32900),
            .in1(N__32574),
            .in2(N__32778),
            .in3(N__32272),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48705),
            .ce(),
            .sr(N__48216));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_13_24_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_13_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_13_24_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_13_24_5  (
            .in0(N__32571),
            .in1(N__32759),
            .in2(N__32925),
            .in3(N__32251),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48705),
            .ce(),
            .sr(N__48216));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_13_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_13_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_13_24_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_13_24_6  (
            .in0(N__32901),
            .in1(N__32575),
            .in2(N__32779),
            .in3(N__32230),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48705),
            .ce(),
            .sr(N__48216));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_13_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_13_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_13_24_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_13_24_7  (
            .in0(N__32572),
            .in1(N__32760),
            .in2(N__32926),
            .in3(N__32209),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48705),
            .ce(),
            .sr(N__48216));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_13_25_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_13_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_13_25_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_13_25_0  (
            .in0(N__32581),
            .in1(N__32907),
            .in2(N__32773),
            .in3(N__32188),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48222));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_13_25_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_13_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_13_25_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_13_25_1  (
            .in0(N__32904),
            .in1(N__32584),
            .in2(N__32770),
            .in3(N__33082),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48222));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_13_25_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_13_25_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_13_25_2 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_13_25_2  (
            .in0(N__33061),
            .in1(N__32737),
            .in2(N__32595),
            .in3(N__32913),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48222));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_13_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_13_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_13_25_3 .LUT_INIT=16'b1010101010000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_13_25_3  (
            .in0(N__33037),
            .in1(N__32744),
            .in2(N__32923),
            .in3(N__32590),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48222));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_13_25_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_13_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_13_25_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_13_25_4  (
            .in0(N__32582),
            .in1(N__32908),
            .in2(N__32774),
            .in3(N__33013),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48222));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_13_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_13_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_13_25_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_13_25_5  (
            .in0(N__32905),
            .in1(N__32585),
            .in2(N__32771),
            .in3(N__32992),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48222));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_13_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_13_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_13_25_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_13_25_6  (
            .in0(N__32583),
            .in1(N__32909),
            .in2(N__32775),
            .in3(N__32971),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48222));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_13_25_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_13_25_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_13_25_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_13_25_7  (
            .in0(N__32906),
            .in1(N__32586),
            .in2(N__32772),
            .in3(N__32947),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48703),
            .ce(),
            .sr(N__48222));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_13_26_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_13_26_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_13_26_5 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_13_26_5  (
            .in0(N__32924),
            .in1(N__32785),
            .in2(N__32776),
            .in3(N__32580),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48701),
            .ce(),
            .sr(N__48224));
    defparam \phase_controller_inst1.S2_LC_13_27_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_27_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39694),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48700),
            .ce(),
            .sr(N__48229));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_14_8_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_14_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_14_8_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_19_LC_14_8_5  (
            .in0(N__42270),
            .in1(N__42042),
            .in2(N__42195),
            .in3(N__44845),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48825),
            .ce(),
            .sr(N__48097));
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_14_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_14_8_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_31_LC_14_8_6  (
            .in0(N__33632),
            .in1(N__36339),
            .in2(_gnd_net_),
            .in3(N__33455),
            .lcout(measured_delay_hc_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48825),
            .ce(),
            .sr(N__48097));
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_9_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_9_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_12_LC_14_9_5  (
            .in0(N__36319),
            .in1(N__33412),
            .in2(_gnd_net_),
            .in3(N__36646),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48815),
            .ce(N__36226),
            .sr(N__48105));
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_14_10_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_14_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_14_10_0 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_14_LC_14_10_0  (
            .in0(N__36584),
            .in1(_gnd_net_),
            .in2(N__36367),
            .in3(N__33364),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48808),
            .ce(N__36231),
            .sr(N__48111));
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_14_10_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_14_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_14_10_1 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_16_LC_14_10_1  (
            .in0(N__33309),
            .in1(N__36344),
            .in2(_gnd_net_),
            .in3(N__36585),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48808),
            .ce(N__36231),
            .sr(N__48111));
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_14_10_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_14_10_2 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_17_LC_14_10_2  (
            .in0(N__36586),
            .in1(_gnd_net_),
            .in2(N__36368),
            .in3(N__33259),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48808),
            .ce(N__36231),
            .sr(N__48111));
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_14_10_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_14_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_14_10_3 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_18_LC_14_10_3  (
            .in0(N__33211),
            .in1(N__36348),
            .in2(_gnd_net_),
            .in3(N__36587),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48808),
            .ce(N__36231),
            .sr(N__48111));
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_14_10_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_14_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_14_10_4 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_19_LC_14_10_4  (
            .in0(N__36340),
            .in1(N__33163),
            .in2(_gnd_net_),
            .in3(N__33129),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48808),
            .ce(N__36231),
            .sr(N__48111));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_14_10_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_14_10_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(N__45456),
            .in2(_gnd_net_),
            .in3(N__45365),
            .lcout(\phase_controller_slave.stoper_tr.time_passed11 ),
            .ltout(\phase_controller_slave.stoper_tr.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_10_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_10_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33691),
            .in3(N__45870),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_11_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(N__33688),
            .in2(N__38407),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_11_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__38380),
            .in2(_gnd_net_),
            .in3(N__33682),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_11_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(N__33790),
            .in2(N__38362),
            .in3(N__33679),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_11_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(N__38329),
            .in2(_gnd_net_),
            .in3(N__33676),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_11_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__38311),
            .in2(_gnd_net_),
            .in3(N__33673),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_11_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__38281),
            .in2(_gnd_net_),
            .in3(N__33670),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_11_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(N__38251),
            .in2(_gnd_net_),
            .in3(N__33667),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_11_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__38218),
            .in2(_gnd_net_),
            .in3(N__33718),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_12_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__38611),
            .in2(_gnd_net_),
            .in3(N__33715),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_12_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_12_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38581),
            .in3(N__33712),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_12_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__45778),
            .in2(_gnd_net_),
            .in3(N__33709),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_12_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__38524),
            .in2(_gnd_net_),
            .in3(N__33706),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_12_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_12_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38506),
            .in3(N__33703),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_12_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__38458),
            .in2(_gnd_net_),
            .in3(N__33700),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_12_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__38425),
            .in2(_gnd_net_),
            .in3(N__33697),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_12_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(N__38734),
            .in2(_gnd_net_),
            .in3(N__33694),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_13_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__38713),
            .in2(_gnd_net_),
            .in3(N__33799),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_13_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_13_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38695),
            .in3(N__33796),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_13_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__38674),
            .in2(_gnd_net_),
            .in3(N__33793),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_14_13_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_14_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__45900),
            .in2(_gnd_net_),
            .in3(N__45861),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_14_13_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_14_13_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__42219),
            .in2(_gnd_net_),
            .in3(N__41967),
            .lcout(\phase_controller_slave.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33779),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_14_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_14_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__33742),
            .in2(N__34143),
            .in3(N__34136),
            .lcout(\current_shift_inst.un38_control_input_0 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_14_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_14_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__33736),
            .in2(_gnd_net_),
            .in3(N__33730),
            .lcout(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_14_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_14_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__33727),
            .in2(_gnd_net_),
            .in3(N__33721),
            .lcout(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_14_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_14_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__36784),
            .in2(_gnd_net_),
            .in3(N__33826),
            .lcout(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_14_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_14_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__36778),
            .in2(_gnd_net_),
            .in3(N__33823),
            .lcout(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_14_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_14_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__36874),
            .in2(_gnd_net_),
            .in3(N__33820),
            .lcout(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_14_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_14_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__36868),
            .in2(_gnd_net_),
            .in3(N__33817),
            .lcout(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_14_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_14_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__36862),
            .in2(_gnd_net_),
            .in3(N__33814),
            .lcout(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_14_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__36856),
            .in2(_gnd_net_),
            .in3(N__33811),
            .lcout(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_14_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__36850),
            .in2(_gnd_net_),
            .in3(N__33808),
            .lcout(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_14_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__36844),
            .in2(_gnd_net_),
            .in3(N__33805),
            .lcout(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_14_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__36934),
            .in2(_gnd_net_),
            .in3(N__33802),
            .lcout(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_14_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__37192),
            .in2(_gnd_net_),
            .in3(N__33853),
            .lcout(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_14_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__43525),
            .in2(_gnd_net_),
            .in3(N__33850),
            .lcout(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_14_15_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36916),
            .in3(N__33847),
            .lcout(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_14_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36907),
            .in3(N__33844),
            .lcout(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_14_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__36922),
            .in2(_gnd_net_),
            .in3(N__33841),
            .lcout(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_14_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__36898),
            .in2(_gnd_net_),
            .in3(N__33838),
            .lcout(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_14_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__36928),
            .in2(_gnd_net_),
            .in3(N__33835),
            .lcout(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_14_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__36880),
            .in2(_gnd_net_),
            .in3(N__33832),
            .lcout(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_14_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__37201),
            .in2(_gnd_net_),
            .in3(N__33829),
            .lcout(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_14_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_14_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__36838),
            .in2(_gnd_net_),
            .in3(N__33880),
            .lcout(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_14_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_14_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__36892),
            .in2(_gnd_net_),
            .in3(N__33877),
            .lcout(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_14_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_14_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__43510),
            .in2(_gnd_net_),
            .in3(N__33874),
            .lcout(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_14_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__37063),
            .in2(_gnd_net_),
            .in3(N__33871),
            .lcout(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_14_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__37081),
            .in2(_gnd_net_),
            .in3(N__33868),
            .lcout(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_14_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__36886),
            .in2(_gnd_net_),
            .in3(N__33865),
            .lcout(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_14_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_14_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__37069),
            .in2(_gnd_net_),
            .in3(N__33862),
            .lcout(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_14_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_14_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__37075),
            .in2(_gnd_net_),
            .in3(N__33859),
            .lcout(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_14_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_14_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__37087),
            .in2(_gnd_net_),
            .in3(N__33856),
            .lcout(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_29 ),
            .carryout(\current_shift_inst.un4_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_14_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_14_17_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__37409),
            .in2(_gnd_net_),
            .in3(N__34192),
            .lcout(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_14_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_14_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__41036),
            .in2(_gnd_net_),
            .in3(N__34783),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_14_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_14_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__34161),
            .in2(N__34117),
            .in3(N__34144),
            .lcout(G_407),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\current_shift_inst.z_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_14_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_14_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__34095),
            .in2(N__34078),
            .in3(N__37328),
            .lcout(G_406),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_0 ),
            .carryout(\current_shift_inst.z_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_14_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_14_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_2_c_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__37267),
            .in2(N__34058),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_1 ),
            .carryout(\current_shift_inst.z_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_14_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_14_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_3_c_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__37255),
            .in2(N__34032),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_2 ),
            .carryout(\current_shift_inst.z_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_14_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_14_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_4_c_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__33989),
            .in2(N__37243),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_3 ),
            .carryout(\current_shift_inst.z_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_14_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_14_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_5_c_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__37228),
            .in2(N__33943),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_4 ),
            .carryout(\current_shift_inst.z_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_14_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_14_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_6_c_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__33897),
            .in2(N__37216),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_5 ),
            .carryout(\current_shift_inst.z_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_14_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_14_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_7_c_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__34505),
            .in2(N__37582),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_6 ),
            .carryout(\current_shift_inst.z_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_14_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_14_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_8_c_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__37564),
            .in2(N__34478),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\current_shift_inst.z_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_14_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_14_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_9_c_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__34421),
            .in2(N__37549),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_8 ),
            .carryout(\current_shift_inst.z_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_14_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_14_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_10_c_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__37534),
            .in2(N__34393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_9 ),
            .carryout(\current_shift_inst.z_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_14_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_14_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_11_c_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__37522),
            .in2(N__34356),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_10 ),
            .carryout(\current_shift_inst.z_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_14_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_14_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_12_c_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__34307),
            .in2(N__37510),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_11 ),
            .carryout(\current_shift_inst.z_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_14_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_14_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_13_c_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__37495),
            .in2(N__34268),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_12 ),
            .carryout(\current_shift_inst.z_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_14_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_14_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_14_c_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__34219),
            .in2(N__37483),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_13 ),
            .carryout(\current_shift_inst.z_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_14_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_14_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_15_c_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__34865),
            .in2(N__37705),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_14 ),
            .carryout(\current_shift_inst.z_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_14_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_14_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_16_c_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__34829),
            .in2(N__37687),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\current_shift_inst.z_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_14_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_14_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_17_c_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__37669),
            .in2(N__34794),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_16 ),
            .carryout(\current_shift_inst.z_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_14_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_14_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_18_c_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__34748),
            .in2(N__37654),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_17 ),
            .carryout(\current_shift_inst.z_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_14_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_14_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_19_c_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__37636),
            .in2(N__34722),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_18 ),
            .carryout(\current_shift_inst.z_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_14_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_14_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_20_c_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__37624),
            .in2(N__34687),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_19 ),
            .carryout(\current_shift_inst.z_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_14_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_14_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_21_c_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__37609),
            .in2(N__34635),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_20 ),
            .carryout(\current_shift_inst.z_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_14_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_14_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_22_c_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__37597),
            .in2(N__34594),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_21 ),
            .carryout(\current_shift_inst.z_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_14_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_14_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_23_c_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__34550),
            .in2(N__37855),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_22 ),
            .carryout(\current_shift_inst.z_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_14_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_14_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_24_c_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__35118),
            .in2(N__37837),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\current_shift_inst.z_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_14_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_14_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_25_c_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__37819),
            .in2(N__35091),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_24 ),
            .carryout(\current_shift_inst.z_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_14_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_14_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_26_c_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__35055),
            .in2(N__37804),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_25 ),
            .carryout(\current_shift_inst.z_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_14_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_14_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_27_c_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__35028),
            .in2(N__37786),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_26 ),
            .carryout(\current_shift_inst.z_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_14_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_14_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_28_c_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__37768),
            .in2(N__35001),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_27 ),
            .carryout(\current_shift_inst.z_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_14_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_14_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_29_c_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__34958),
            .in2(N__37753),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_28 ),
            .carryout(\current_shift_inst.z_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_14_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_14_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_30_c_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__37735),
            .in2(N__34926),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_29 ),
            .carryout(\current_shift_inst.z_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_14_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_14_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.un10_control_input_z_s_31_LC_14_21_7  (
            .in0(N__37427),
            .in1(N__37717),
            .in2(N__41847),
            .in3(N__34897),
            .lcout(\current_shift_inst.z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.counter_0_LC_14_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_0_LC_14_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_0_LC_14_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_0_LC_14_22_0  (
            .in0(N__35584),
            .in1(N__40118),
            .in2(_gnd_net_),
            .in3(N__35158),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_0 ),
            .clk(N__48717),
            .ce(N__35480),
            .sr(N__48198));
    defparam \current_shift_inst.timer_phase.counter_1_LC_14_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_1_LC_14_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_1_LC_14_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_1_LC_14_22_1  (
            .in0(N__35579),
            .in1(N__40083),
            .in2(_gnd_net_),
            .in3(N__35155),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_1 ),
            .clk(N__48717),
            .ce(N__35480),
            .sr(N__48198));
    defparam \current_shift_inst.timer_phase.counter_2_LC_14_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_2_LC_14_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_2_LC_14_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_2_LC_14_22_2  (
            .in0(N__35585),
            .in1(N__40016),
            .in2(_gnd_net_),
            .in3(N__35152),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_2 ),
            .clk(N__48717),
            .ce(N__35480),
            .sr(N__48198));
    defparam \current_shift_inst.timer_phase.counter_3_LC_14_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_3_LC_14_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_3_LC_14_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_3_LC_14_22_3  (
            .in0(N__35580),
            .in1(N__39953),
            .in2(_gnd_net_),
            .in3(N__35149),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_3 ),
            .clk(N__48717),
            .ce(N__35480),
            .sr(N__48198));
    defparam \current_shift_inst.timer_phase.counter_4_LC_14_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_4_LC_14_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_4_LC_14_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_4_LC_14_22_4  (
            .in0(N__35586),
            .in1(N__40721),
            .in2(_gnd_net_),
            .in3(N__35146),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_4 ),
            .clk(N__48717),
            .ce(N__35480),
            .sr(N__48198));
    defparam \current_shift_inst.timer_phase.counter_5_LC_14_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_5_LC_14_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_5_LC_14_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_5_LC_14_22_5  (
            .in0(N__35581),
            .in1(N__40652),
            .in2(_gnd_net_),
            .in3(N__35143),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_5 ),
            .clk(N__48717),
            .ce(N__35480),
            .sr(N__48198));
    defparam \current_shift_inst.timer_phase.counter_6_LC_14_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_6_LC_14_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_6_LC_14_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_6_LC_14_22_6  (
            .in0(N__35583),
            .in1(N__40580),
            .in2(_gnd_net_),
            .in3(N__35140),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_6 ),
            .clk(N__48717),
            .ce(N__35480),
            .sr(N__48198));
    defparam \current_shift_inst.timer_phase.counter_7_LC_14_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_7_LC_14_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_7_LC_14_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_7_LC_14_22_7  (
            .in0(N__35582),
            .in1(N__40520),
            .in2(_gnd_net_),
            .in3(N__35137),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_7 ),
            .clk(N__48717),
            .ce(N__35480),
            .sr(N__48198));
    defparam \current_shift_inst.timer_phase.counter_8_LC_14_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_8_LC_14_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_8_LC_14_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_8_LC_14_23_0  (
            .in0(N__35590),
            .in1(N__40442),
            .in2(_gnd_net_),
            .in3(N__35134),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_8 ),
            .clk(N__48711),
            .ce(N__35476),
            .sr(N__48206));
    defparam \current_shift_inst.timer_phase.counter_9_LC_14_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_9_LC_14_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_9_LC_14_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_9_LC_14_23_1  (
            .in0(N__35594),
            .in1(N__40358),
            .in2(_gnd_net_),
            .in3(N__35185),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_9 ),
            .clk(N__48711),
            .ce(N__35476),
            .sr(N__48206));
    defparam \current_shift_inst.timer_phase.counter_10_LC_14_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_10_LC_14_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_10_LC_14_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_10_LC_14_23_2  (
            .in0(N__35587),
            .in1(N__40298),
            .in2(_gnd_net_),
            .in3(N__35182),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_10 ),
            .clk(N__48711),
            .ce(N__35476),
            .sr(N__48206));
    defparam \current_shift_inst.timer_phase.counter_11_LC_14_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_11_LC_14_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_11_LC_14_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_11_LC_14_23_3  (
            .in0(N__35591),
            .in1(N__40217),
            .in2(_gnd_net_),
            .in3(N__35179),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_11 ),
            .clk(N__48711),
            .ce(N__35476),
            .sr(N__48206));
    defparam \current_shift_inst.timer_phase.counter_12_LC_14_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_12_LC_14_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_12_LC_14_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_12_LC_14_23_4  (
            .in0(N__35588),
            .in1(N__41207),
            .in2(_gnd_net_),
            .in3(N__35176),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_12 ),
            .clk(N__48711),
            .ce(N__35476),
            .sr(N__48206));
    defparam \current_shift_inst.timer_phase.counter_13_LC_14_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_13_LC_14_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_13_LC_14_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_13_LC_14_23_5  (
            .in0(N__35592),
            .in1(N__41132),
            .in2(_gnd_net_),
            .in3(N__35173),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_13 ),
            .clk(N__48711),
            .ce(N__35476),
            .sr(N__48206));
    defparam \current_shift_inst.timer_phase.counter_14_LC_14_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_14_LC_14_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_14_LC_14_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_14_LC_14_23_6  (
            .in0(N__35589),
            .in1(N__41063),
            .in2(_gnd_net_),
            .in3(N__35170),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_14 ),
            .clk(N__48711),
            .ce(N__35476),
            .sr(N__48206));
    defparam \current_shift_inst.timer_phase.counter_15_LC_14_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_15_LC_14_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_15_LC_14_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_15_LC_14_23_7  (
            .in0(N__35593),
            .in1(N__41000),
            .in2(_gnd_net_),
            .in3(N__35167),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_15 ),
            .clk(N__48711),
            .ce(N__35476),
            .sr(N__48206));
    defparam \current_shift_inst.timer_phase.counter_16_LC_14_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_16_LC_14_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_16_LC_14_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_16_LC_14_24_0  (
            .in0(N__35595),
            .in1(N__40928),
            .in2(_gnd_net_),
            .in3(N__35164),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_16 ),
            .clk(N__48709),
            .ce(N__35481),
            .sr(N__48212));
    defparam \current_shift_inst.timer_phase.counter_17_LC_14_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_17_LC_14_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_17_LC_14_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_17_LC_14_24_1  (
            .in0(N__35601),
            .in1(N__40862),
            .in2(_gnd_net_),
            .in3(N__35161),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_17 ),
            .clk(N__48709),
            .ce(N__35481),
            .sr(N__48212));
    defparam \current_shift_inst.timer_phase.counter_18_LC_14_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_18_LC_14_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_18_LC_14_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_18_LC_14_24_2  (
            .in0(N__35596),
            .in1(N__40793),
            .in2(_gnd_net_),
            .in3(N__35212),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_18 ),
            .clk(N__48709),
            .ce(N__35481),
            .sr(N__48212));
    defparam \current_shift_inst.timer_phase.counter_19_LC_14_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_19_LC_14_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_19_LC_14_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_19_LC_14_24_3  (
            .in0(N__35602),
            .in1(N__41750),
            .in2(_gnd_net_),
            .in3(N__35209),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_19 ),
            .clk(N__48709),
            .ce(N__35481),
            .sr(N__48212));
    defparam \current_shift_inst.timer_phase.counter_20_LC_14_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_20_LC_14_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_20_LC_14_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_20_LC_14_24_4  (
            .in0(N__35597),
            .in1(N__41678),
            .in2(_gnd_net_),
            .in3(N__35206),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_20 ),
            .clk(N__48709),
            .ce(N__35481),
            .sr(N__48212));
    defparam \current_shift_inst.timer_phase.counter_21_LC_14_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_21_LC_14_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_21_LC_14_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_21_LC_14_24_5  (
            .in0(N__35603),
            .in1(N__41606),
            .in2(_gnd_net_),
            .in3(N__35203),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_21 ),
            .clk(N__48709),
            .ce(N__35481),
            .sr(N__48212));
    defparam \current_shift_inst.timer_phase.counter_22_LC_14_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_22_LC_14_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_22_LC_14_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_22_LC_14_24_6  (
            .in0(N__35598),
            .in1(N__41546),
            .in2(_gnd_net_),
            .in3(N__35200),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_22 ),
            .clk(N__48709),
            .ce(N__35481),
            .sr(N__48212));
    defparam \current_shift_inst.timer_phase.counter_23_LC_14_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_23_LC_14_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_23_LC_14_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_23_LC_14_24_7  (
            .in0(N__35604),
            .in1(N__41484),
            .in2(_gnd_net_),
            .in3(N__35197),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_23 ),
            .clk(N__48709),
            .ce(N__35481),
            .sr(N__48212));
    defparam \current_shift_inst.timer_phase.counter_24_LC_14_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_24_LC_14_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_24_LC_14_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_24_LC_14_25_0  (
            .in0(N__35605),
            .in1(N__41426),
            .in2(_gnd_net_),
            .in3(N__35194),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_24 ),
            .clk(N__48706),
            .ce(N__35482),
            .sr(N__48217));
    defparam \current_shift_inst.timer_phase.counter_25_LC_14_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_25_LC_14_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_25_LC_14_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_25_LC_14_25_1  (
            .in0(N__35599),
            .in1(N__41354),
            .in2(_gnd_net_),
            .in3(N__35191),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_25 ),
            .clk(N__48706),
            .ce(N__35482),
            .sr(N__48217));
    defparam \current_shift_inst.timer_phase.counter_26_LC_14_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_26_LC_14_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_26_LC_14_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_26_LC_14_25_2  (
            .in0(N__35606),
            .in1(N__41270),
            .in2(_gnd_net_),
            .in3(N__35188),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_26 ),
            .clk(N__48706),
            .ce(N__35482),
            .sr(N__48217));
    defparam \current_shift_inst.timer_phase.counter_27_LC_14_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_27_LC_14_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_27_LC_14_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_27_LC_14_25_3  (
            .in0(N__35600),
            .in1(N__41927),
            .in2(_gnd_net_),
            .in3(N__35614),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_27 ),
            .clk(N__48706),
            .ce(N__35482),
            .sr(N__48217));
    defparam \current_shift_inst.timer_phase.counter_28_LC_14_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_28_LC_14_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_28_LC_14_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_28_LC_14_25_4  (
            .in0(N__35607),
            .in1(N__41286),
            .in2(_gnd_net_),
            .in3(N__35611),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_28 ),
            .clk(N__48706),
            .ce(N__35482),
            .sr(N__48217));
    defparam \current_shift_inst.timer_phase.counter_29_LC_14_25_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.counter_29_LC_14_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_29_LC_14_25_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_phase.counter_29_LC_14_25_5  (
            .in0(N__41904),
            .in1(N__35608),
            .in2(_gnd_net_),
            .in3(N__35485),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48706),
            .ce(N__35482),
            .sr(N__48217));
    defparam SB_DFF_inst_DELAY_TR1_LC_15_5_5.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR1_LC_15_5_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR1_LC_15_5_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_DELAY_TR1_LC_15_5_5 (
            .in0(N__35443),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(delay_tr_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48854),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR2_LC_15_6_6.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR2_LC_15_6_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR2_LC_15_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR2_LC_15_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35434),
            .lcout(delay_tr_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48846),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_15_7_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_15_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_15_7_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_7_LC_15_7_7  (
            .in0(N__36667),
            .in1(N__36335),
            .in2(_gnd_net_),
            .in3(N__35428),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48840),
            .ce(N__36222),
            .sr(N__48089));
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_15_8_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_15_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_15_8_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_2_LC_15_8_1  (
            .in0(N__36663),
            .in1(N__36315),
            .in2(N__35801),
            .in3(N__35374),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48835),
            .ce(N__36232),
            .sr(N__48092));
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_15_8_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_15_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_15_8_2 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_15_8_2  (
            .in0(N__35319),
            .in1(N__35791),
            .in2(N__36357),
            .in3(N__36661),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48835),
            .ce(N__36232),
            .sr(N__48092));
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_15_8_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_15_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_15_8_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_4_LC_15_8_3  (
            .in0(N__36665),
            .in1(N__36317),
            .in2(N__35803),
            .in3(N__35265),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48835),
            .ce(N__36232),
            .sr(N__48092));
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_15_8_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_15_8_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_5_LC_15_8_4  (
            .in0(N__36318),
            .in1(N__36151),
            .in2(_gnd_net_),
            .in3(N__36666),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48835),
            .ce(N__36232),
            .sr(N__48092));
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_15_8_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_15_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_15_8_5 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_3_LC_15_8_5  (
            .in0(N__36664),
            .in1(N__36316),
            .in2(N__35802),
            .in3(N__36085),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48835),
            .ce(N__36232),
            .sr(N__48092));
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_15_8_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_13_LC_15_8_6  (
            .in0(N__36314),
            .in1(N__36031),
            .in2(_gnd_net_),
            .in3(N__36662),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48835),
            .ce(N__36232),
            .sr(N__48092));
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_15_9_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_15_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_15_9_1 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_9_LC_15_9_1  (
            .in0(N__36653),
            .in1(N__35983),
            .in2(N__36361),
            .in3(N__35780),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48826),
            .ce(N__36227),
            .sr(N__48098));
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_15_9_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_15_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_15_9_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_10_LC_15_9_2  (
            .in0(N__35932),
            .in1(N__36321),
            .in2(_gnd_net_),
            .in3(N__36648),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48826),
            .ce(N__36227),
            .sr(N__48098));
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_15_9_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_15_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_15_9_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_11_LC_15_9_3  (
            .in0(N__36649),
            .in1(_gnd_net_),
            .in2(N__36358),
            .in3(N__35890),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48826),
            .ce(N__36227),
            .sr(N__48098));
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_15_9_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_15_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_15_9_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_0_LC_15_9_4  (
            .in0(N__35778),
            .in1(N__36320),
            .in2(N__35848),
            .in3(N__36647),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48826),
            .ce(N__36227),
            .sr(N__48098));
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_15_9_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_15_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_15_9_5 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_1_LC_15_9_5  (
            .in0(N__36651),
            .in1(N__35779),
            .in2(N__36359),
            .in3(N__35708),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48826),
            .ce(N__36227),
            .sr(N__48098));
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_15_9_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_15_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_15_9_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_15_LC_15_9_6  (
            .in0(N__35668),
            .in1(N__36325),
            .in2(_gnd_net_),
            .in3(N__36650),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48826),
            .ce(N__36227),
            .sr(N__48098));
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_15_9_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_15_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_15_9_7 .LUT_INIT=16'b0000100000001000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_8_LC_15_9_7  (
            .in0(N__36652),
            .in1(N__36491),
            .in2(N__36360),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48826),
            .ce(N__36227),
            .sr(N__48098));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_15_10_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_15_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_15_10_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_7_LC_15_10_0  (
            .in0(N__42005),
            .in1(N__42152),
            .in2(N__42306),
            .in3(N__44227),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48816),
            .ce(),
            .sr(N__48106));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_15_10_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_15_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_15_10_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_9_LC_15_10_2  (
            .in0(N__42006),
            .in1(N__42153),
            .in2(N__42307),
            .in3(N__44710),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48816),
            .ce(),
            .sr(N__48106));
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_15_10_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_15_10_3 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_15_10_3  (
            .in0(N__42151),
            .in1(_gnd_net_),
            .in2(N__42271),
            .in3(N__42004),
            .lcout(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_10_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_10_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_10_4  (
            .in0(N__45896),
            .in1(N__38406),
            .in2(_gnd_net_),
            .in3(N__45871),
            .lcout(),
            .ltout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_10_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_10_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_10_5  (
            .in0(N__45626),
            .in1(N__45458),
            .in2(N__36235),
            .in3(N__45374),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48816),
            .ce(),
            .sr(N__48106));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_15_10_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_15_10_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_15_10_6  (
            .in0(N__42003),
            .in1(N__42150),
            .in2(_gnd_net_),
            .in3(N__42250),
            .lcout(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_15_10_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_15_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_15_10_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_10_LC_15_10_7  (
            .in0(N__45625),
            .in1(N__45457),
            .in2(N__45394),
            .in3(N__36178),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48816),
            .ce(),
            .sr(N__48106));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_15_11_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_15_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_15_11_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_2_LC_15_11_0  (
            .in0(N__45507),
            .in1(N__45390),
            .in2(N__45650),
            .in3(N__36169),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48809),
            .ce(),
            .sr(N__48112));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_15_11_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_15_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_15_11_1 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_3_LC_15_11_1  (
            .in0(N__45384),
            .in1(N__45512),
            .in2(N__36160),
            .in3(N__45619),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48809),
            .ce(),
            .sr(N__48112));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_15_11_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_15_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_15_11_2 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_4_LC_15_11_2  (
            .in0(N__45508),
            .in1(N__36736),
            .in2(N__45647),
            .in3(N__45387),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48809),
            .ce(),
            .sr(N__48112));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_15_11_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_15_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_15_11_3 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_5_LC_15_11_3  (
            .in0(N__45385),
            .in1(N__45513),
            .in2(N__36730),
            .in3(N__45620),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48809),
            .ce(),
            .sr(N__48112));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_15_11_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_15_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_15_11_4 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_6_LC_15_11_4  (
            .in0(N__45509),
            .in1(N__36721),
            .in2(N__45648),
            .in3(N__45388),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48809),
            .ce(),
            .sr(N__48112));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_15_11_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_15_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_15_11_5 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_7_LC_15_11_5  (
            .in0(N__45386),
            .in1(N__45514),
            .in2(N__36715),
            .in3(N__45621),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48809),
            .ce(),
            .sr(N__48112));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_15_11_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_15_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_15_11_6 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_8_LC_15_11_6  (
            .in0(N__45510),
            .in1(N__36706),
            .in2(N__45649),
            .in3(N__45389),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48809),
            .ce(),
            .sr(N__48112));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_11_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_11_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_11_7  (
            .in0(N__45383),
            .in1(N__45511),
            .in2(N__36700),
            .in3(N__45618),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48809),
            .ce(),
            .sr(N__48112));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_12_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_12_0 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_12_0  (
            .in0(N__45378),
            .in1(N__45630),
            .in2(N__36691),
            .in3(N__45506),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48797),
            .ce(),
            .sr(N__48120));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_12_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_12_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_12_1  (
            .in0(N__45499),
            .in1(N__45379),
            .in2(N__45651),
            .in3(N__36682),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48797),
            .ce(),
            .sr(N__48120));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_12_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_12_2 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_12_2  (
            .in0(N__45375),
            .in1(N__45627),
            .in2(N__36676),
            .in3(N__45503),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48797),
            .ce(),
            .sr(N__48120));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_12_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_12_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_12_3  (
            .in0(N__45500),
            .in1(N__45380),
            .in2(N__45652),
            .in3(N__36772),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48797),
            .ce(),
            .sr(N__48120));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_15_12_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_15_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_15_12_4 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_16_LC_15_12_4  (
            .in0(N__45376),
            .in1(N__45628),
            .in2(N__36766),
            .in3(N__45504),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48797),
            .ce(),
            .sr(N__48120));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_12_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_12_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_12_5  (
            .in0(N__45501),
            .in1(N__45381),
            .in2(N__45653),
            .in3(N__36757),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48797),
            .ce(),
            .sr(N__48120));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_15_12_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_15_12_6 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_18_LC_15_12_6  (
            .in0(N__45377),
            .in1(N__45629),
            .in2(N__36751),
            .in3(N__45505),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48797),
            .ce(),
            .sr(N__48120));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_12_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_12_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_12_7  (
            .in0(N__45502),
            .in1(N__45382),
            .in2(N__45654),
            .in3(N__36742),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48797),
            .ce(),
            .sr(N__48120));
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_15_13_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_15_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_15_13_0 .LUT_INIT=16'b0100010001000101;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_6_LC_15_13_0  (
            .in0(N__45034),
            .in1(N__38955),
            .in2(N__45165),
            .in3(N__44974),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48789),
            .ce(N__45212),
            .sr(N__48126));
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_15_13_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_15_13_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_4_LC_15_13_1  (
            .in0(N__44973),
            .in1(N__45157),
            .in2(N__46570),
            .in3(N__45033),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48789),
            .ce(N__45212),
            .sr(N__48126));
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_15_13_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_15_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_15_13_2 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_7_LC_15_13_2  (
            .in0(N__39004),
            .in1(_gnd_net_),
            .in2(N__45166),
            .in3(N__44972),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48789),
            .ce(N__45212),
            .sr(N__48126));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_15_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_15_13_3 .LUT_INIT=16'b0001010100010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_15_13_3  (
            .in0(N__38896),
            .in1(N__36828),
            .in2(N__39219),
            .in3(N__38825),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_15_13_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_15_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_15_13_4 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_8_LC_15_13_4  (
            .in0(N__45164),
            .in1(_gnd_net_),
            .in2(N__36832),
            .in3(N__39045),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48789),
            .ce(N__45212),
            .sr(N__48126));
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_15_13_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_15_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_15_13_6 .LUT_INIT=16'b1111111100110001;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_9_LC_15_13_6  (
            .in0(N__38826),
            .in1(N__37011),
            .in2(N__38912),
            .in3(N__39214),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48789),
            .ce(N__45212),
            .sr(N__48126));
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_15_13_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_15_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_15_13_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_14_LC_15_13_7  (
            .in0(N__38897),
            .in1(N__45156),
            .in2(_gnd_net_),
            .in3(N__36829),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48789),
            .ce(N__45212),
            .sr(N__48126));
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_15_14_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_15_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_15_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_10_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__37005),
            .in2(_gnd_net_),
            .in3(N__37108),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48781),
            .ce(N__45211),
            .sr(N__48130));
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_15_14_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_15_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_15_14_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_11_LC_15_14_1  (
            .in0(N__37129),
            .in1(_gnd_net_),
            .in2(N__37012),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48781),
            .ce(N__45211),
            .sr(N__48130));
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_15_14_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_15_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_15_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_12_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__37009),
            .in2(_gnd_net_),
            .in3(N__37180),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48781),
            .ce(N__45211),
            .sr(N__48130));
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_15_14_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_15_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_15_14_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_13_LC_15_14_3  (
            .in0(N__37010),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37152),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48781),
            .ce(N__45211),
            .sr(N__48130));
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_15_14_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_15_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_15_14_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_15_LC_15_14_4  (
            .in0(N__45155),
            .in1(_gnd_net_),
            .in2(N__38917),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48781),
            .ce(N__45211),
            .sr(N__48130));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39364),
            .lcout(\current_shift_inst.un4_control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39355),
            .lcout(\current_shift_inst.un4_control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39346),
            .lcout(\current_shift_inst.un4_control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_15_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_15_15_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__39123),
            .in2(_gnd_net_),
            .in3(N__46386),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_15_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_15_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_15_15_1  (
            .in0(N__37179),
            .in1(N__37128),
            .in2(N__37153),
            .in3(N__37107),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39337),
            .lcout(\current_shift_inst.un4_control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39328),
            .lcout(\current_shift_inst.un4_control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39319),
            .lcout(\current_shift_inst.un4_control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39310),
            .lcout(\current_shift_inst.un4_control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39301),
            .lcout(\current_shift_inst.un4_control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_15_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_15_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39493),
            .lcout(\current_shift_inst.un4_control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_15_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_15_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39292),
            .lcout(\current_shift_inst.un4_control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_15_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_15_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39382),
            .lcout(\current_shift_inst.un4_control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39400),
            .lcout(\current_shift_inst.un4_control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39418),
            .lcout(\current_shift_inst.un4_control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39409),
            .lcout(\current_shift_inst.un4_control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_15_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_15_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39391),
            .lcout(\current_shift_inst.un4_control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39484),
            .lcout(\current_shift_inst.un4_control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_15_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_15_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39454),
            .lcout(\current_shift_inst.un4_control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_15_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_15_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39373),
            .lcout(\current_shift_inst.un4_control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_15_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_15_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39889),
            .lcout(\current_shift_inst.un4_control_input_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39463),
            .lcout(\current_shift_inst.un4_control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_15_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_15_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39898),
            .lcout(\current_shift_inst.un4_control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_15_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_15_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39445),
            .lcout(\current_shift_inst.un4_control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_15_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_15_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39472),
            .lcout(\current_shift_inst.un4_control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__36989),
            .in2(_gnd_net_),
            .in3(N__37106),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48750),
            .ce(N__46643),
            .sr(N__48154));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_18_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_15_18_1  (
            .in0(N__36990),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37127),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48750),
            .ce(N__46643),
            .sr(N__48154));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__36991),
            .in2(_gnd_net_),
            .in3(N__37172),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48750),
            .ce(N__46643),
            .sr(N__48154));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_18_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_15_18_3  (
            .in0(N__36992),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37148),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48750),
            .ce(N__46643),
            .sr(N__48154));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_15_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_15_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39502),
            .lcout(\current_shift_inst.un4_control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_15_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_15_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39433),
            .lcout(\current_shift_inst.un4_control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_15_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_15_19_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_15_19_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_12_LC_15_19_0  (
            .in0(N__49102),
            .in1(N__44081),
            .in2(_gnd_net_),
            .in3(N__46696),
            .lcout(measured_delay_tr_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48744),
            .ce(N__46343),
            .sr(N__48161));
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_15_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_15_19_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_15_19_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_13_LC_15_19_1  (
            .in0(N__44082),
            .in1(N__49103),
            .in2(_gnd_net_),
            .in3(N__47482),
            .lcout(measured_delay_tr_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48744),
            .ce(N__46343),
            .sr(N__48161));
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_15_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_15_19_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_15_19_2 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_5_LC_15_19_2  (
            .in0(N__46417),
            .in1(N__46502),
            .in2(N__45973),
            .in3(N__46165),
            .lcout(measured_delay_tr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48744),
            .ce(N__46343),
            .sr(N__48161));
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_15_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_15_19_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_15_19_3 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_11_LC_15_19_3  (
            .in0(N__44080),
            .in1(N__49101),
            .in2(_gnd_net_),
            .in3(N__46744),
            .lcout(measured_delay_tr_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48744),
            .ce(N__46343),
            .sr(N__48161));
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_15_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_15_19_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_10_LC_15_19_4  (
            .in0(N__49100),
            .in1(N__44079),
            .in2(_gnd_net_),
            .in3(N__46789),
            .lcout(measured_delay_tr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48744),
            .ce(N__46343),
            .sr(N__48161));
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_15_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_15_19_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_15_19_5 .LUT_INIT=16'b0100010111001111;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_6_LC_15_19_5  (
            .in0(N__46503),
            .in1(N__47020),
            .in2(N__46168),
            .in3(N__46418),
            .lcout(measured_delay_tr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48744),
            .ce(N__46343),
            .sr(N__48161));
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_15_19_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_15_19_7 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_9_LC_15_19_7  (
            .in0(N__44083),
            .in1(N__49104),
            .in2(N__46864),
            .in3(N__46416),
            .lcout(measured_delay_tr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48744),
            .ce(N__46343),
            .sr(N__48161));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_15_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_15_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_15_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40084),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48737),
            .ce(N__41821),
            .sr(N__48171));
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_15_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_15_20_2 .LUT_INIT=16'b0101010101100101;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_15_20_2  (
            .in0(N__40101),
            .in1(N__37286),
            .in2(N__37443),
            .in3(N__37321),
            .lcout(\current_shift_inst.N_1742_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_15_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_15_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40129),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48737),
            .ce(N__41821),
            .sr(N__48171));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_15_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_15_20_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_15_20_5  (
            .in0(N__37322),
            .in1(N__40102),
            .in2(N__37293),
            .in3(N__37431),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_15_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_15_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__37317),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\current_shift_inst.z_5_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_15_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_15_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__37285),
            .in2(N__43357),
            .in3(N__37258),
            .lcout(\current_shift_inst.z_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_1 ),
            .carryout(\current_shift_inst.z_5_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_15_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_15_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__40095),
            .in2(N__43361),
            .in3(N__37246),
            .lcout(\current_shift_inst.z_5_3 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_2 ),
            .carryout(\current_shift_inst.z_5_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_15_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_15_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__40037),
            .in2(N__43358),
            .in3(N__37231),
            .lcout(\current_shift_inst.z_5_4 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_3 ),
            .carryout(\current_shift_inst.z_5_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_15_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_15_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__39971),
            .in2(N__43362),
            .in3(N__37219),
            .lcout(\current_shift_inst.z_5_5 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_4 ),
            .carryout(\current_shift_inst.z_5_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_15_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_15_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__39917),
            .in2(N__43359),
            .in3(N__37204),
            .lcout(\current_shift_inst.z_5_6 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_5 ),
            .carryout(\current_shift_inst.z_5_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_15_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_15_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__40679),
            .in2(N__43363),
            .in3(N__37567),
            .lcout(\current_shift_inst.z_5_7 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_6 ),
            .carryout(\current_shift_inst.z_5_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_15_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_15_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__40606),
            .in2(N__43360),
            .in3(N__37552),
            .lcout(\current_shift_inst.z_5_8 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_7 ),
            .carryout(\current_shift_inst.z_5_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_15_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_15_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__40541),
            .in2(N__43467),
            .in3(N__37537),
            .lcout(\current_shift_inst.z_5_9 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\current_shift_inst.z_5_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_15_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_15_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__40472),
            .in2(N__43450),
            .in3(N__37525),
            .lcout(\current_shift_inst.z_5_10 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_9 ),
            .carryout(\current_shift_inst.z_5_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_15_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_15_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__40393),
            .in2(N__43464),
            .in3(N__37513),
            .lcout(\current_shift_inst.z_5_11 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_10 ),
            .carryout(\current_shift_inst.z_5_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_15_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_15_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__40319),
            .in2(N__43451),
            .in3(N__37498),
            .lcout(\current_shift_inst.z_5_12 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_11 ),
            .carryout(\current_shift_inst.z_5_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_15_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_15_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__40243),
            .in2(N__43465),
            .in3(N__37486),
            .lcout(\current_shift_inst.z_5_13 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_12 ),
            .carryout(\current_shift_inst.z_5_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_15_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_15_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__40163),
            .in2(N__43452),
            .in3(N__37468),
            .lcout(\current_shift_inst.z_5_14 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_13 ),
            .carryout(\current_shift_inst.z_5_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_15_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_15_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__41159),
            .in2(N__43466),
            .in3(N__37690),
            .lcout(\current_shift_inst.z_5_15 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_14 ),
            .carryout(\current_shift_inst.z_5_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_15_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_15_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(N__41090),
            .in2(N__43453),
            .in3(N__37672),
            .lcout(\current_shift_inst.z_5_16 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_15 ),
            .carryout(\current_shift_inst.z_5_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_15_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_15_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__41021),
            .in2(N__43454),
            .in3(N__37657),
            .lcout(\current_shift_inst.z_5_17 ),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\current_shift_inst.z_5_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_15_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_15_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(N__40958),
            .in2(N__43468),
            .in3(N__37639),
            .lcout(\current_shift_inst.z_5_18 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_17 ),
            .carryout(\current_shift_inst.z_5_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_15_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_15_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__40887),
            .in2(N__43455),
            .in3(N__37627),
            .lcout(\current_shift_inst.z_5_19 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_18 ),
            .carryout(\current_shift_inst.z_5_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_15_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_15_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__40814),
            .in2(N__43469),
            .in3(N__37612),
            .lcout(\current_shift_inst.z_5_20 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_19 ),
            .carryout(\current_shift_inst.z_5_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_15_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_15_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(N__40748),
            .in2(N__43456),
            .in3(N__37600),
            .lcout(\current_shift_inst.z_5_21 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_20 ),
            .carryout(\current_shift_inst.z_5_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_15_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_15_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__41705),
            .in2(N__43470),
            .in3(N__37585),
            .lcout(\current_shift_inst.z_5_22 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_21 ),
            .carryout(\current_shift_inst.z_5_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_15_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_15_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__41638),
            .in2(N__43457),
            .in3(N__37840),
            .lcout(\current_shift_inst.z_5_23 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_22 ),
            .carryout(\current_shift_inst.z_5_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_15_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_15_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_15_23_7  (
            .in0(_gnd_net_),
            .in1(N__41570),
            .in2(N__43471),
            .in3(N__37822),
            .lcout(\current_shift_inst.z_5_24 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_23 ),
            .carryout(\current_shift_inst.z_5_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_15_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_15_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(N__41510),
            .in2(N__43458),
            .in3(N__37807),
            .lcout(\current_shift_inst.z_5_25 ),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\current_shift_inst.z_5_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_15_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_15_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__41450),
            .in2(N__43461),
            .in3(N__37789),
            .lcout(\current_shift_inst.z_5_26 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_25 ),
            .carryout(\current_shift_inst.z_5_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_15_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_15_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(N__41384),
            .in2(N__43459),
            .in3(N__37771),
            .lcout(\current_shift_inst.z_5_27 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_26 ),
            .carryout(\current_shift_inst.z_5_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_15_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_15_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__41311),
            .in2(N__43462),
            .in3(N__37756),
            .lcout(\current_shift_inst.z_5_28 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_27 ),
            .carryout(\current_shift_inst.z_5_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_15_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_15_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(N__41231),
            .in2(N__43460),
            .in3(N__37738),
            .lcout(\current_shift_inst.z_5_29 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_28 ),
            .carryout(\current_shift_inst.z_5_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_15_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_15_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(N__41873),
            .in2(N__43463),
            .in3(N__37723),
            .lcout(\current_shift_inst.z_5_30 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_29 ),
            .carryout(\current_shift_inst.z_5_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_15_24_6 .C_ON=1'b0;
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_15_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_15_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37720),
            .lcout(\current_shift_inst.z_5_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC1_LC_16_4_6.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC1_LC_16_4_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC1_LC_16_4_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_DELAY_HC1_LC_16_4_6 (
            .in0(N__37975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(delay_hc_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48862),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_16_8_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_16_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37957),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_16_8_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_16_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__37948),
            .in2(N__37942),
            .in3(N__44393),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_16_8_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_16_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__37924),
            .in2(N__37933),
            .in3(N__44376),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_16_8_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_16_8_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_16_8_3  (
            .in0(N__44340),
            .in1(N__37909),
            .in2(N__37918),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_16_8_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_16_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__37891),
            .in2(N__37903),
            .in3(N__44319),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_16_8_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_16_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(N__37876),
            .in2(N__37885),
            .in3(N__44292),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_16_8_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_16_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__37861),
            .in2(N__37870),
            .in3(N__44268),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_16_8_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_16_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_16_8_7  (
            .in0(N__44244),
            .in1(N__38098),
            .in2(N__38110),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_16_9_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_16_9_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_16_9_0  (
            .in0(N__44748),
            .in1(N__38083),
            .in2(N__38092),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_16_9_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_16_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__38068),
            .in2(N__38077),
            .in3(N__44721),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_16_9_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_16_9_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_16_9_2  (
            .in0(N__44694),
            .in1(N__38053),
            .in2(N__38062),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_16_9_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_16_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__38038),
            .in2(N__38047),
            .in3(N__44673),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_16_9_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_16_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__38020),
            .in2(N__38032),
            .in3(N__44652),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_16_9_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_16_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__38005),
            .in2(N__38014),
            .in3(N__44631),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_16_9_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_16_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__37981),
            .in2(N__37999),
            .in3(N__44610),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_16_9_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_16_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(N__38194),
            .in2(N__38206),
            .in3(N__44589),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_16_10_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_16_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__38176),
            .in2(N__38188),
            .in3(N__44943),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_16_10_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_16_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__38158),
            .in2(N__38170),
            .in3(N__44922),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_16_10_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_16_10_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_16_10_2  (
            .in0(N__44889),
            .in1(N__38140),
            .in2(N__38152),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_16_10_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_16_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__38119),
            .in2(N__38134),
            .in3(N__44865),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_10_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38113),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_16_10_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_16_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__42630),
            .in2(_gnd_net_),
            .in3(N__42590),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_16_10_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_16_10_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_16_10_7  (
            .in0(N__42591),
            .in1(_gnd_net_),
            .in2(N__42634),
            .in3(N__44397),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_11_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__38386),
            .in2(N__39244),
            .in3(N__38402),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_11_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_11_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_11_1  (
            .in0(N__38379),
            .in1(N__38368),
            .in2(N__39058),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_11_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_11_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_11_2  (
            .in0(N__38358),
            .in1(N__38347),
            .in2(N__39232),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_11_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__38317),
            .in2(N__38341),
            .in3(N__38328),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_11_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__38299),
            .in2(N__38758),
            .in3(N__38310),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_11_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__38269),
            .in2(N__38293),
            .in3(N__38280),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_11_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__38239),
            .in2(N__38263),
            .in3(N__38250),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_11_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__38626),
            .in2(N__38233),
            .in3(N__38217),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_12_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__38599),
            .in2(N__38620),
            .in3(N__38610),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_12_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__38560),
            .in2(N__38593),
            .in3(N__38577),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_12_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__38542),
            .in2(N__38554),
            .in3(N__45774),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_12_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__38512),
            .in2(N__38536),
            .in3(N__38523),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_12_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_12_4  (
            .in0(N__38502),
            .in1(N__38476),
            .in2(N__38491),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_12_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__38446),
            .in2(N__38470),
            .in3(N__38457),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_12_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(N__38413),
            .in2(N__38440),
            .in3(N__38424),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_12_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(N__45235),
            .in2(N__38722),
            .in3(N__38733),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_13_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(N__38701),
            .in2(N__38653),
            .in3(N__38712),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_13_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__38680),
            .in2(N__38644),
            .in3(N__38691),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_13_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__38662),
            .in2(N__38635),
            .in3(N__38673),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_13_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38656),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_16_13_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_16_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_16_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_17_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39787),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48798),
            .ce(N__45223),
            .sr(N__48121));
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_16_13_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_16_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_16_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_18_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39831),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48798),
            .ce(N__45223),
            .sr(N__48121));
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_16_13_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_16_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_16_13_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_19_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__39741),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48798),
            .ce(N__45223),
            .sr(N__48121));
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_16_14_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_16_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_16_14_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_1_LC_16_14_0  (
            .in0(N__39279),
            .in1(N__39146),
            .in2(N__39268),
            .in3(N__39089),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48790),
            .ce(N__45219),
            .sr(N__48127));
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_16_14_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_16_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_16_14_1 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_3_LC_16_14_1  (
            .in0(N__39091),
            .in1(_gnd_net_),
            .in2(N__39150),
            .in3(N__39129),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48790),
            .ce(N__45219),
            .sr(N__48127));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_16_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_16_14_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_16_14_3  (
            .in0(N__38824),
            .in1(N__39215),
            .in2(N__38926),
            .in3(N__39181),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_16_14_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_16_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_16_14_4 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_2_LC_16_14_4  (
            .in0(N__39130),
            .in1(N__46390),
            .in2(N__39094),
            .in3(N__39090),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48790),
            .ce(N__45219),
            .sr(N__48127));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_16_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_16_14_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_16_14_5  (
            .in0(N__39046),
            .in1(N__39002),
            .in2(_gnd_net_),
            .in3(N__38954),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_16_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_16_14_6 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__38913),
            .in2(N__38836),
            .in3(N__38823),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_16_14_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_16_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_16_14_7 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_5_LC_16_14_7  (
            .in0(N__38800),
            .in1(N__45141),
            .in2(N__38761),
            .in3(N__44975),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48790),
            .ce(N__45219),
            .sr(N__48127));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__42498),
            .in2(N__42567),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__48782),
            .ce(N__39880),
            .sr(N__48131));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__42474),
            .in2(N__42531),
            .in3(N__39358),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__48782),
            .ce(N__39880),
            .sr(N__48131));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__42499),
            .in2(N__42450),
            .in3(N__39349),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__48782),
            .ce(N__39880),
            .sr(N__48131));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__42475),
            .in2(N__42420),
            .in3(N__39340),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__48782),
            .ce(N__39880),
            .sr(N__48131));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__42390),
            .in2(N__42451),
            .in3(N__39331),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__48782),
            .ce(N__39880),
            .sr(N__48131));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__42366),
            .in2(N__42421),
            .in3(N__39322),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__48782),
            .ce(N__39880),
            .sr(N__48131));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__42391),
            .in2(N__42859),
            .in3(N__39313),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__48782),
            .ce(N__39880),
            .sr(N__48131));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__42367),
            .in2(N__42828),
            .in3(N__39304),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__48782),
            .ce(N__39880),
            .sr(N__48131));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__42858),
            .in2(N__42796),
            .in3(N__39295),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__48773),
            .ce(N__39879),
            .sr(N__48136));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__42765),
            .in2(N__42829),
            .in3(N__39436),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__48773),
            .ce(N__39879),
            .sr(N__48136));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__42795),
            .in2(N__42741),
            .in3(N__39424),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__48773),
            .ce(N__39879),
            .sr(N__48136));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__42766),
            .in2(N__42711),
            .in3(N__39421),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__48773),
            .ce(N__39879),
            .sr(N__48136));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(N__42681),
            .in2(N__42742),
            .in3(N__39412),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__48773),
            .ce(N__39879),
            .sr(N__48136));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(N__42657),
            .in2(N__42712),
            .in3(N__39403),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__48773),
            .ce(N__39879),
            .sr(N__48136));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(N__42682),
            .in2(N__43114),
            .in3(N__39394),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__48773),
            .ce(N__39879),
            .sr(N__48136));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_16_7  (
            .in0(_gnd_net_),
            .in1(N__42658),
            .in2(N__43084),
            .in3(N__39385),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__48773),
            .ce(N__39879),
            .sr(N__48136));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(N__43113),
            .in2(N__43053),
            .in3(N__39376),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__48763),
            .ce(N__39877),
            .sr(N__48142));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__43083),
            .in2(N__43024),
            .in3(N__39367),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__48763),
            .ce(N__39877),
            .sr(N__48142));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(N__42993),
            .in2(N__43054),
            .in3(N__39496),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__48763),
            .ce(N__39877),
            .sr(N__48142));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(N__43023),
            .in2(N__42969),
            .in3(N__39487),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__48763),
            .ce(N__39877),
            .sr(N__48142));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__42994),
            .in2(N__42940),
            .in3(N__39478),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__48763),
            .ce(N__39877),
            .sr(N__48142));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__42909),
            .in2(N__42970),
            .in3(N__39475),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__48763),
            .ce(N__39877),
            .sr(N__48142));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__42939),
            .in2(N__42886),
            .in3(N__39466),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__48763),
            .ce(N__39877),
            .sr(N__48142));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(N__42910),
            .in2(N__43837),
            .in3(N__39457),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__48763),
            .ce(N__39877),
            .sr(N__48142));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(N__42885),
            .in2(N__43806),
            .in3(N__39448),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__48756),
            .ce(N__39876),
            .sr(N__48148));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__43836),
            .in2(N__43777),
            .in3(N__39439),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__48756),
            .ce(N__39876),
            .sr(N__48148));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(N__43747),
            .in2(N__43807),
            .in3(N__39892),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__48756),
            .ce(N__39876),
            .sr(N__48148));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__43776),
            .in2(N__43597),
            .in3(N__39883),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__48756),
            .ce(N__39876),
            .sr(N__48148));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39856),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_16_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_16_19_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_16_19_0  (
            .in0(N__39824),
            .in1(N__39782),
            .in2(N__39745),
            .in3(N__45263),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5PP_2_LC_16_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5PP_2_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5PP_2_LC_16_19_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5PP_2_LC_16_19_1  (
            .in0(N__46474),
            .in1(N__47428),
            .in2(N__46086),
            .in3(N__46030),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_16_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_16_19_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_16_19_2  (
            .in0(N__46916),
            .in1(N__46970),
            .in2(_gnd_net_),
            .in3(N__47019),
            .lcout(\delay_measurement_inst.N_425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.T01_sbtinv_LC_16_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_sbtinv_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.T01_sbtinv_LC_16_19_3 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \phase_controller_inst1.T01_sbtinv_LC_16_19_3  (
            .in0(N__39690),
            .in1(N__39642),
            .in2(N__39604),
            .in3(N__39553),
            .lcout(\phase_controller_inst1.N_221_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9DQM6_10_LC_16_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9DQM6_10_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9DQM6_10_LC_16_19_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9DQM6_10_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__44097),
            .in2(_gnd_net_),
            .in3(N__46219),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_424_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_16_19_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_16_19_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_16_19_7  (
            .in0(N__40147),
            .in1(N__46501),
            .in2(N__39505),
            .in3(N__40138),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_16_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_16_20_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_16_20_1  (
            .in0(N__47354),
            .in1(N__44098),
            .in2(_gnd_net_),
            .in3(N__46220),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_4_LC_16_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_4_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_4_LC_16_20_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_4_LC_16_20_4  (
            .in0(N__47418),
            .in1(N__46029),
            .in2(N__47363),
            .in3(N__45968),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICTS5M_31_LC_16_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICTS5M_31_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICTS5M_31_LC_16_20_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICTS5M_31_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__48275),
            .in2(_gnd_net_),
            .in3(N__43851),
            .lcout(\delay_measurement_inst.N_280_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_16_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_16_21_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_16_21_5  (
            .in0(N__47172),
            .in1(N__47232),
            .in2(N__47117),
            .in3(N__47289),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_16_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_16_21_6 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_16_21_6  (
            .in0(N__46079),
            .in1(N__46463),
            .in2(N__40141),
            .in3(N__46852),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_16_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_16_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_16_22_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(N__40125),
            .in2(N__40018),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_3 ),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ),
            .clk(N__48732),
            .ce(N__41820),
            .sr(N__48184));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_16_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_16_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_16_22_1  (
            .in0(_gnd_net_),
            .in1(N__40082),
            .in2(N__39955),
            .in3(N__40021),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ),
            .clk(N__48732),
            .ce(N__41820),
            .sr(N__48184));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_16_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_16_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_16_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(N__40017),
            .in2(N__40728),
            .in3(N__39958),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ),
            .clk(N__48732),
            .ce(N__41820),
            .sr(N__48184));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_16_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_16_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(N__39954),
            .in2(N__40659),
            .in3(N__39901),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ),
            .clk(N__48732),
            .ce(N__41820),
            .sr(N__48184));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_16_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_16_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_16_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(N__40581),
            .in2(N__40729),
            .in3(N__40663),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ),
            .clk(N__48732),
            .ce(N__41820),
            .sr(N__48184));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_16_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_16_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_16_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_16_22_5  (
            .in0(_gnd_net_),
            .in1(N__40521),
            .in2(N__40660),
            .in3(N__40585),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ),
            .clk(N__48732),
            .ce(N__41820),
            .sr(N__48184));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_16_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_16_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_16_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_16_22_6  (
            .in0(_gnd_net_),
            .in1(N__40582),
            .in2(N__40453),
            .in3(N__40525),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ),
            .clk(N__48732),
            .ce(N__41820),
            .sr(N__48184));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_16_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_16_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_16_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_16_22_7  (
            .in0(_gnd_net_),
            .in1(N__40522),
            .in2(N__40369),
            .in3(N__40456),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ),
            .clk(N__48732),
            .ce(N__41820),
            .sr(N__48184));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_16_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_16_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_16_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(N__40446),
            .in2(N__40299),
            .in3(N__40372),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_11 ),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ),
            .clk(N__48725),
            .ce(N__41819),
            .sr(N__48192));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_16_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_16_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_16_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_16_23_1  (
            .in0(_gnd_net_),
            .in1(N__40368),
            .in2(N__40219),
            .in3(N__40303),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ),
            .clk(N__48725),
            .ce(N__41819),
            .sr(N__48192));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_16_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_16_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_16_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_16_23_2  (
            .in0(_gnd_net_),
            .in1(N__41208),
            .in2(N__40300),
            .in3(N__40222),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ),
            .clk(N__48725),
            .ce(N__41819),
            .sr(N__48192));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_16_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_16_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_16_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(N__40218),
            .in2(N__41139),
            .in3(N__41212),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ),
            .clk(N__48725),
            .ce(N__41819),
            .sr(N__48192));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_16_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_16_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_16_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(N__41209),
            .in2(N__41070),
            .in3(N__41143),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ),
            .clk(N__48725),
            .ce(N__41819),
            .sr(N__48192));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_16_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_16_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_16_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_16_23_5  (
            .in0(_gnd_net_),
            .in1(N__41001),
            .in2(N__41140),
            .in3(N__41074),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ),
            .clk(N__48725),
            .ce(N__41819),
            .sr(N__48192));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_16_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_16_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_16_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_16_23_6  (
            .in0(_gnd_net_),
            .in1(N__40939),
            .in2(N__41071),
            .in3(N__41005),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ),
            .clk(N__48725),
            .ce(N__41819),
            .sr(N__48192));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_16_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_16_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_16_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_16_23_7  (
            .in0(_gnd_net_),
            .in1(N__41002),
            .in2(N__40873),
            .in3(N__40942),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ),
            .clk(N__48725),
            .ce(N__41819),
            .sr(N__48192));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_16_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_16_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_16_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_16_24_0  (
            .in0(_gnd_net_),
            .in1(N__40938),
            .in2(N__40795),
            .in3(N__40876),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_19 ),
            .ltout(),
            .carryin(bfn_16_24_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ),
            .clk(N__48718),
            .ce(N__41818),
            .sr(N__48199));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_16_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_16_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_16_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_16_24_1  (
            .in0(_gnd_net_),
            .in1(N__40866),
            .in2(N__41752),
            .in3(N__40798),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ),
            .clk(N__48718),
            .ce(N__41818),
            .sr(N__48199));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_16_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_16_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_16_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_16_24_2  (
            .in0(_gnd_net_),
            .in1(N__40794),
            .in2(N__41685),
            .in3(N__40732),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ),
            .clk(N__48718),
            .ce(N__41818),
            .sr(N__48199));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_16_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_16_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_16_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(N__41751),
            .in2(N__41613),
            .in3(N__41689),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ),
            .clk(N__48718),
            .ce(N__41818),
            .sr(N__48199));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_16_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_16_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_16_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_16_24_4  (
            .in0(_gnd_net_),
            .in1(N__41547),
            .in2(N__41686),
            .in3(N__41617),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ),
            .clk(N__48718),
            .ce(N__41818),
            .sr(N__48199));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_16_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_16_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_16_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_16_24_5  (
            .in0(_gnd_net_),
            .in1(N__41490),
            .in2(N__41614),
            .in3(N__41554),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ),
            .clk(N__48718),
            .ce(N__41818),
            .sr(N__48199));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_16_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_16_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_16_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_16_24_6  (
            .in0(_gnd_net_),
            .in1(N__41431),
            .in2(N__41551),
            .in3(N__41494),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ),
            .clk(N__48718),
            .ce(N__41818),
            .sr(N__48199));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_16_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_16_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_16_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_16_24_7  (
            .in0(_gnd_net_),
            .in1(N__41491),
            .in2(N__41365),
            .in3(N__41434),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ),
            .clk(N__48718),
            .ce(N__41818),
            .sr(N__48199));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_16_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_16_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_16_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_16_25_0  (
            .in0(_gnd_net_),
            .in1(N__41430),
            .in2(N__41271),
            .in3(N__41368),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_27 ),
            .ltout(),
            .carryin(bfn_16_25_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ),
            .clk(N__48712),
            .ce(N__41817),
            .sr(N__48207));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_16_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_16_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_16_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_16_25_1  (
            .in0(_gnd_net_),
            .in1(N__41364),
            .in2(N__41932),
            .in3(N__41290),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ),
            .clk(N__48712),
            .ce(N__41817),
            .sr(N__48207));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_16_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_16_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_16_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_16_25_2  (
            .in0(_gnd_net_),
            .in1(N__41287),
            .in2(N__41272),
            .in3(N__41215),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ),
            .clk(N__48712),
            .ce(N__41817),
            .sr(N__48207));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_16_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_16_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_16_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_16_25_3  (
            .in0(_gnd_net_),
            .in1(N__41931),
            .in2(N__41908),
            .in3(N__41857),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ),
            .clk(N__48712),
            .ce(N__41817),
            .sr(N__48207));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_16_25_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_16_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_16_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_16_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41854),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48712),
            .ce(N__41817),
            .sr(N__48207));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_16_26_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_16_26_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_16_26_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_16_26_3  (
            .in0(N__47548),
            .in1(N__47581),
            .in2(N__47518),
            .in3(N__47617),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_16_26_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_16_26_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_16_26_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_16_26_4  (
            .in0(N__47056),
            .in1(N__41797),
            .in2(N__41800),
            .in3(N__41791),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_27_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_27_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_27_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_27_6  (
            .in0(N__47686),
            .in1(N__47716),
            .in2(N__47656),
            .in3(N__47752),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_16_28_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_16_28_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_16_28_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_16_28_6  (
            .in0(_gnd_net_),
            .in1(N__49144),
            .in2(_gnd_net_),
            .in3(N__49192),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_17_5_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_17_5_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_17_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_17_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41782),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48863),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_17_6_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_17_6_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_17_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_17_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41767),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48859),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_17_8_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_17_8_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_5_LC_17_8_0  (
            .in0(N__42310),
            .in1(N__42174),
            .in2(N__44281),
            .in3(N__42057),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48847),
            .ce(),
            .sr(N__48088));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_17_8_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_17_8_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_8_LC_17_8_1  (
            .in0(N__42054),
            .in1(N__42314),
            .in2(N__42190),
            .in3(N__44737),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48847),
            .ce(),
            .sr(N__48088));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_8_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_8_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_8_2  (
            .in0(N__42308),
            .in1(N__42172),
            .in2(N__44905),
            .in3(N__42055),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48847),
            .ce(),
            .sr(N__48088));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_17_8_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_17_8_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_2_LC_17_8_3  (
            .in0(N__42051),
            .in1(N__42311),
            .in2(N__42187),
            .in3(N__44365),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48847),
            .ce(),
            .sr(N__48088));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_17_8_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_17_8_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_6_LC_17_8_5  (
            .in0(N__42053),
            .in1(N__42313),
            .in2(N__42189),
            .in3(N__44257),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48847),
            .ce(),
            .sr(N__48088));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_17_8_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_17_8_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_4_LC_17_8_6  (
            .in0(N__42309),
            .in1(N__42173),
            .in2(N__44308),
            .in3(N__42056),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48847),
            .ce(),
            .sr(N__48088));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_17_8_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_17_8_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_3_LC_17_8_7  (
            .in0(N__42052),
            .in1(N__42312),
            .in2(N__42188),
            .in3(N__44329),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48847),
            .ce(),
            .sr(N__48088));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_17_9_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_17_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_17_9_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_10_LC_17_9_0  (
            .in0(N__42315),
            .in1(N__42047),
            .in2(N__42175),
            .in3(N__44683),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48841),
            .ce(),
            .sr(N__48090));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_9_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_9_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_9_1  (
            .in0(N__42045),
            .in1(N__42136),
            .in2(N__42333),
            .in3(N__44878),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48841),
            .ce(),
            .sr(N__48090));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_9_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_9_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_9_2  (
            .in0(N__42317),
            .in1(N__42049),
            .in2(N__42177),
            .in3(N__44641),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48841),
            .ce(),
            .sr(N__48090));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_17_9_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_17_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_17_9_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_13_LC_17_9_3  (
            .in0(N__42043),
            .in1(N__42134),
            .in2(N__42331),
            .in3(N__44620),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48841),
            .ce(),
            .sr(N__48090));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_9_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_9_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_9_4  (
            .in0(N__42318),
            .in1(N__42050),
            .in2(N__42178),
            .in3(N__44578),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48841),
            .ce(),
            .sr(N__48090));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_17_9_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_17_9_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_14_LC_17_9_5  (
            .in0(N__42044),
            .in1(N__42135),
            .in2(N__42332),
            .in3(N__44599),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48841),
            .ce(),
            .sr(N__48090));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_17_9_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_17_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_17_9_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_11_LC_17_9_6  (
            .in0(N__42316),
            .in1(N__42048),
            .in2(N__42176),
            .in3(N__44662),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48841),
            .ce(),
            .sr(N__48090));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_17_9_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_17_9_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_1_LC_17_9_7  (
            .in0(N__42046),
            .in1(N__42137),
            .in2(N__42334),
            .in3(N__42343),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48841),
            .ce(),
            .sr(N__48090));
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_17_10_0 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_17_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_0_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__44798),
            .in2(_gnd_net_),
            .in3(N__44821),
            .lcout(),
            .ltout(\phase_controller_slave.N_214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_LC_17_10_1 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_hc_LC_17_10_1 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \phase_controller_slave.start_timer_hc_LC_17_10_1  (
            .in0(N__42132),
            .in1(N__44833),
            .in2(N__42337),
            .in3(N__45937),
            .lcout(\phase_controller_slave.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48836),
            .ce(),
            .sr(N__48093));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_10_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_10_2 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_10_2  (
            .in0(N__42305),
            .in1(N__42133),
            .in2(N__42061),
            .in3(N__44932),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48836),
            .ce(),
            .sr(N__48093));
    defparam \phase_controller_slave.state_2_LC_17_10_3 .C_ON=1'b0;
    defparam \phase_controller_slave.state_2_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_2_LC_17_10_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_slave.state_2_LC_17_10_3  (
            .in0(N__44822),
            .in1(N__45822),
            .in2(N__44805),
            .in3(N__45760),
            .lcout(\phase_controller_slave.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48836),
            .ce(),
            .sr(N__48093));
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_17_10_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_17_10_5 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_LC_17_10_5  (
            .in0(N__44823),
            .in1(N__42629),
            .in2(N__41944),
            .in3(N__42589),
            .lcout(\phase_controller_slave.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48836),
            .ce(),
            .sr(N__48093));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_10_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__42628),
            .in2(_gnd_net_),
            .in3(N__42588),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_17_11_0  (
            .in0(N__43703),
            .in1(N__42554),
            .in2(_gnd_net_),
            .in3(N__42538),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__48827),
            .ce(N__43576),
            .sr(N__48099));
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_17_11_1  (
            .in0(N__43711),
            .in1(N__42518),
            .in2(_gnd_net_),
            .in3(N__42502),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__48827),
            .ce(N__43576),
            .sr(N__48099));
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_17_11_2  (
            .in0(N__43704),
            .in1(N__42497),
            .in2(_gnd_net_),
            .in3(N__42478),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__48827),
            .ce(N__43576),
            .sr(N__48099));
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_17_11_3  (
            .in0(N__43712),
            .in1(N__42468),
            .in2(_gnd_net_),
            .in3(N__42454),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__48827),
            .ce(N__43576),
            .sr(N__48099));
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_17_11_4  (
            .in0(N__43705),
            .in1(N__42438),
            .in2(_gnd_net_),
            .in3(N__42424),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__48827),
            .ce(N__43576),
            .sr(N__48099));
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_17_11_5  (
            .in0(N__43713),
            .in1(N__42408),
            .in2(_gnd_net_),
            .in3(N__42394),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__48827),
            .ce(N__43576),
            .sr(N__48099));
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_17_11_6  (
            .in0(N__43706),
            .in1(N__42384),
            .in2(_gnd_net_),
            .in3(N__42370),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__48827),
            .ce(N__43576),
            .sr(N__48099));
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_17_11_7  (
            .in0(N__43714),
            .in1(N__42360),
            .in2(_gnd_net_),
            .in3(N__42346),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__48827),
            .ce(N__43576),
            .sr(N__48099));
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_17_12_0  (
            .in0(N__43718),
            .in1(N__42848),
            .in2(_gnd_net_),
            .in3(N__42832),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__48817),
            .ce(N__43571),
            .sr(N__48107));
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_17_12_1  (
            .in0(N__43726),
            .in1(N__42815),
            .in2(_gnd_net_),
            .in3(N__42799),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__48817),
            .ce(N__43571),
            .sr(N__48107));
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_17_12_2  (
            .in0(N__43715),
            .in1(N__42791),
            .in2(_gnd_net_),
            .in3(N__42769),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__48817),
            .ce(N__43571),
            .sr(N__48107));
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_17_12_3  (
            .in0(N__43723),
            .in1(N__42764),
            .in2(_gnd_net_),
            .in3(N__42745),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__48817),
            .ce(N__43571),
            .sr(N__48107));
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_17_12_4  (
            .in0(N__43716),
            .in1(N__42729),
            .in2(_gnd_net_),
            .in3(N__42715),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__48817),
            .ce(N__43571),
            .sr(N__48107));
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_17_12_5  (
            .in0(N__43724),
            .in1(N__42699),
            .in2(_gnd_net_),
            .in3(N__42685),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__48817),
            .ce(N__43571),
            .sr(N__48107));
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_17_12_6  (
            .in0(N__43717),
            .in1(N__42675),
            .in2(_gnd_net_),
            .in3(N__42661),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__48817),
            .ce(N__43571),
            .sr(N__48107));
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_17_12_7  (
            .in0(N__43725),
            .in1(N__42651),
            .in2(_gnd_net_),
            .in3(N__42637),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__48817),
            .ce(N__43571),
            .sr(N__48107));
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_17_13_0  (
            .in0(N__43707),
            .in1(N__43103),
            .in2(_gnd_net_),
            .in3(N__43087),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__48810),
            .ce(N__43561),
            .sr(N__48113));
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_17_13_1  (
            .in0(N__43719),
            .in1(N__43073),
            .in2(_gnd_net_),
            .in3(N__43057),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__48810),
            .ce(N__43561),
            .sr(N__48113));
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_17_13_2  (
            .in0(N__43708),
            .in1(N__43046),
            .in2(_gnd_net_),
            .in3(N__43027),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__48810),
            .ce(N__43561),
            .sr(N__48113));
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_17_13_3  (
            .in0(N__43720),
            .in1(N__43019),
            .in2(_gnd_net_),
            .in3(N__42997),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__48810),
            .ce(N__43561),
            .sr(N__48113));
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_17_13_4  (
            .in0(N__43709),
            .in1(N__42987),
            .in2(_gnd_net_),
            .in3(N__42973),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__48810),
            .ce(N__43561),
            .sr(N__48113));
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_17_13_5  (
            .in0(N__43721),
            .in1(N__42957),
            .in2(_gnd_net_),
            .in3(N__42943),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__48810),
            .ce(N__43561),
            .sr(N__48113));
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_17_13_6  (
            .in0(N__43710),
            .in1(N__42929),
            .in2(_gnd_net_),
            .in3(N__42913),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__48810),
            .ce(N__43561),
            .sr(N__48113));
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_17_13_7  (
            .in0(N__43722),
            .in1(N__42903),
            .in2(_gnd_net_),
            .in3(N__42889),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__48810),
            .ce(N__43561),
            .sr(N__48113));
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_17_14_0  (
            .in0(N__43643),
            .in1(N__42875),
            .in2(_gnd_net_),
            .in3(N__43840),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__48799),
            .ce(N__43572),
            .sr(N__48122));
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_17_14_1  (
            .in0(N__43647),
            .in1(N__43826),
            .in2(_gnd_net_),
            .in3(N__43810),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__48799),
            .ce(N__43572),
            .sr(N__48122));
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_17_14_2  (
            .in0(N__43644),
            .in1(N__43799),
            .in2(_gnd_net_),
            .in3(N__43780),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__48799),
            .ce(N__43572),
            .sr(N__48122));
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_17_14_3  (
            .in0(N__43648),
            .in1(N__43772),
            .in2(_gnd_net_),
            .in3(N__43750),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__48799),
            .ce(N__43572),
            .sr(N__48122));
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_17_14_4  (
            .in0(N__43645),
            .in1(N__43743),
            .in2(_gnd_net_),
            .in3(N__43729),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__48799),
            .ce(N__43572),
            .sr(N__48122));
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_14_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_17_14_5  (
            .in0(N__43590),
            .in1(N__43646),
            .in2(_gnd_net_),
            .in3(N__43600),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48799),
            .ce(N__43572),
            .sr(N__48122));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43531),
            .lcout(\current_shift_inst.un4_control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43516),
            .lcout(\current_shift_inst.un4_control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_17_17_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_17_17_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_17_17_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_17_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_17_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_tr_LC_17_18_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_17_18_0  (
            .in0(N__43985),
            .in1(N__44014),
            .in2(_gnd_net_),
            .in3(N__43943),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48764),
            .ce(),
            .sr(N__48143));
    defparam \delay_measurement_inst.prev_tr_sig_LC_17_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_tr_sig_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_tr_sig_LC_17_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_tr_sig_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43986),
            .lcout(\delay_measurement_inst.prev_tr_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48764),
            .ce(),
            .sr(N__48143));
    defparam \delay_measurement_inst.stop_timer_tr_LC_17_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_tr_LC_17_18_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__43908),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48764),
            .ce(),
            .sr(N__48143));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_17_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_17_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_17_18_4 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_17_18_4  (
            .in0(N__44131),
            .in1(N__44116),
            .in2(_gnd_net_),
            .in3(N__44058),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48764),
            .ce(),
            .sr(N__48143));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9IAF_1_LC_17_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9IAF_1_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9IAF_1_LC_17_19_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9IAF_1_LC_17_19_1  (
            .in0(N__47018),
            .in1(N__45969),
            .in2(N__46860),
            .in3(N__48895),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI200N_7_LC_17_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI200N_7_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI200N_7_LC_17_19_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI200N_7_LC_17_19_2  (
            .in0(N__46917),
            .in1(_gnd_net_),
            .in2(N__43924),
            .in3(N__46971),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_2_LC_17_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_2_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_2_LC_17_19_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_2_LC_17_19_3  (
            .in0(N__43921),
            .in1(N__46268),
            .in2(N__43915),
            .in3(N__46415),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_390_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5KUTL_31_LC_17_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5KUTL_31_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5KUTL_31_LC_17_19_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5KUTL_31_LC_17_19_4  (
            .in0(N__49095),
            .in1(N__43912),
            .in2(N__43888),
            .in3(N__43885),
            .lcout(\delay_measurement_inst.N_280_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_17_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_17_19_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__44114),
            .in2(_gnd_net_),
            .in3(N__44056),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_338_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_19_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_19_7 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_19_7  (
            .in0(N__44057),
            .in1(N__44127),
            .in2(_gnd_net_),
            .in3(N__44115),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_339_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_17_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_17_20_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_17_20_1  (
            .in0(N__46692),
            .in1(N__46740),
            .in2(N__47481),
            .in3(N__46788),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_17_20_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_17_20_2 .LUT_INIT=16'b0001000100110001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_17_20_2  (
            .in0(N__47425),
            .in1(N__47361),
            .in2(N__44086),
            .in3(N__46856),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_17_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_17_20_4 .LUT_INIT=16'b0000000011001101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_17_20_4  (
            .in0(N__47426),
            .in1(N__46270),
            .in2(N__47364),
            .in3(N__46241),
            .lcout(\delay_measurement_inst.N_409_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_17_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_17_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44059),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_17_21_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_17_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_17_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46051),
            .lcout(\delay_measurement_inst.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48745),
            .ce(N__48338),
            .sr(N__48162));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_17_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_17_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_17_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45270),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48738),
            .ce(N__46648),
            .sr(N__48172));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_23_0  (
            .in0(N__44545),
            .in1(N__48911),
            .in2(_gnd_net_),
            .in3(N__44020),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__48733),
            .ce(N__44440),
            .sr(N__48185));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_23_1  (
            .in0(N__44540),
            .in1(N__46046),
            .in2(_gnd_net_),
            .in3(N__44017),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__48733),
            .ce(N__44440),
            .sr(N__48185));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_23_2  (
            .in0(N__44546),
            .in1(N__45992),
            .in2(_gnd_net_),
            .in3(N__44158),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__48733),
            .ce(N__44440),
            .sr(N__48185));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_23_3  (
            .in0(N__44541),
            .in1(N__47039),
            .in2(_gnd_net_),
            .in3(N__44155),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__48733),
            .ce(N__44440),
            .sr(N__48185));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_23_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_23_4  (
            .in0(N__44547),
            .in1(N__46993),
            .in2(_gnd_net_),
            .in3(N__44152),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__48733),
            .ce(N__44440),
            .sr(N__48185));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_23_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_23_5  (
            .in0(N__44542),
            .in1(N__46939),
            .in2(_gnd_net_),
            .in3(N__44149),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__48733),
            .ce(N__44440),
            .sr(N__48185));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_23_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_23_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_23_6  (
            .in0(N__44544),
            .in1(N__46883),
            .in2(_gnd_net_),
            .in3(N__44146),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__48733),
            .ce(N__44440),
            .sr(N__48185));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_23_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_23_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_23_7  (
            .in0(N__44543),
            .in1(N__46808),
            .in2(_gnd_net_),
            .in3(N__44143),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__48733),
            .ce(N__44440),
            .sr(N__48185));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_24_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_24_0  (
            .in0(N__44551),
            .in1(N__46761),
            .in2(_gnd_net_),
            .in3(N__44140),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_24_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__48726),
            .ce(N__44442),
            .sr(N__48193));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_24_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_24_1  (
            .in0(N__44569),
            .in1(N__46713),
            .in2(_gnd_net_),
            .in3(N__44137),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__48726),
            .ce(N__44442),
            .sr(N__48193));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_24_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_24_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_24_2  (
            .in0(N__44548),
            .in1(N__47501),
            .in2(_gnd_net_),
            .in3(N__44134),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__48726),
            .ce(N__44442),
            .sr(N__48193));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_24_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_24_3  (
            .in0(N__44566),
            .in1(N__47447),
            .in2(_gnd_net_),
            .in3(N__44185),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__48726),
            .ce(N__44442),
            .sr(N__48193));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_24_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_24_4  (
            .in0(N__44549),
            .in1(N__47380),
            .in2(_gnd_net_),
            .in3(N__44182),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__48726),
            .ce(N__44442),
            .sr(N__48193));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_24_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_24_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_24_5  (
            .in0(N__44567),
            .in1(N__47308),
            .in2(_gnd_net_),
            .in3(N__44179),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__48726),
            .ce(N__44442),
            .sr(N__48193));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_24_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_24_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_24_6  (
            .in0(N__44550),
            .in1(N__47252),
            .in2(_gnd_net_),
            .in3(N__44176),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__48726),
            .ce(N__44442),
            .sr(N__48193));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_24_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_24_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_24_7  (
            .in0(N__44568),
            .in1(N__47198),
            .in2(_gnd_net_),
            .in3(N__44173),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__48726),
            .ce(N__44442),
            .sr(N__48193));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_25_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_25_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_25_0  (
            .in0(N__44552),
            .in1(N__47139),
            .in2(_gnd_net_),
            .in3(N__44170),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_25_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__48719),
            .ce(N__44441),
            .sr(N__48200));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_25_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_25_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_25_1  (
            .in0(N__44556),
            .in1(N__47073),
            .in2(_gnd_net_),
            .in3(N__44167),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__48719),
            .ce(N__44441),
            .sr(N__48200));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_25_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_25_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_25_2  (
            .in0(N__44553),
            .in1(N__47771),
            .in2(_gnd_net_),
            .in3(N__44164),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__48719),
            .ce(N__44441),
            .sr(N__48200));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_25_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_25_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_25_3  (
            .in0(N__44557),
            .in1(N__47735),
            .in2(_gnd_net_),
            .in3(N__44161),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__48719),
            .ce(N__44441),
            .sr(N__48200));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_25_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_25_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_25_4  (
            .in0(N__44554),
            .in1(N__47701),
            .in2(_gnd_net_),
            .in3(N__44212),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__48719),
            .ce(N__44441),
            .sr(N__48200));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_25_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_25_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_25_5  (
            .in0(N__44558),
            .in1(N__47671),
            .in2(_gnd_net_),
            .in3(N__44209),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__48719),
            .ce(N__44441),
            .sr(N__48200));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_25_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_25_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_25_6  (
            .in0(N__44555),
            .in1(N__47636),
            .in2(_gnd_net_),
            .in3(N__44206),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__48719),
            .ce(N__44441),
            .sr(N__48200));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_25_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_25_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_25_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_25_7  (
            .in0(N__44559),
            .in1(N__47600),
            .in2(_gnd_net_),
            .in3(N__44203),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__48719),
            .ce(N__44441),
            .sr(N__48200));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_26_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_26_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_26_0  (
            .in0(N__44560),
            .in1(N__47565),
            .in2(_gnd_net_),
            .in3(N__44200),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_26_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__48713),
            .ce(N__44443),
            .sr(N__48208));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_26_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_26_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_26_1  (
            .in0(N__44564),
            .in1(N__47535),
            .in2(_gnd_net_),
            .in3(N__44197),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__48713),
            .ce(N__44443),
            .sr(N__48208));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_26_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_26_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_26_2  (
            .in0(N__44561),
            .in1(N__49211),
            .in2(_gnd_net_),
            .in3(N__44194),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__48713),
            .ce(N__44443),
            .sr(N__48208));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_26_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_26_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_26_3  (
            .in0(N__44565),
            .in1(N__49163),
            .in2(_gnd_net_),
            .in3(N__44191),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__48713),
            .ce(N__44443),
            .sr(N__48208));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_26_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_26_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_26_4  (
            .in0(N__44562),
            .in1(N__49225),
            .in2(_gnd_net_),
            .in3(N__44188),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__48713),
            .ce(N__44443),
            .sr(N__48208));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_26_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_26_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_26_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_26_5  (
            .in0(N__49177),
            .in1(N__44563),
            .in2(_gnd_net_),
            .in3(N__44446),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48713),
            .ce(N__44443),
            .sr(N__48208));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_8_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_8_0  (
            .in0(_gnd_net_),
            .in1(N__44407),
            .in2(N__44398),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_8_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_8_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_8_1  (
            .in0(_gnd_net_),
            .in1(N__44377),
            .in2(_gnd_net_),
            .in3(N__44359),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_8_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_8_2  (
            .in0(_gnd_net_),
            .in1(N__44356),
            .in2(N__44344),
            .in3(N__44323),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_8_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(N__44320),
            .in2(_gnd_net_),
            .in3(N__44296),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_8_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_8_4  (
            .in0(_gnd_net_),
            .in1(N__44293),
            .in2(_gnd_net_),
            .in3(N__44272),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_8_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_8_5  (
            .in0(_gnd_net_),
            .in1(N__44269),
            .in2(_gnd_net_),
            .in3(N__44251),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_8_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_8_6  (
            .in0(_gnd_net_),
            .in1(N__44248),
            .in2(_gnd_net_),
            .in3(N__44215),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_8_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_8_7  (
            .in0(_gnd_net_),
            .in1(N__44749),
            .in2(_gnd_net_),
            .in3(N__44731),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_9_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_9_0  (
            .in0(_gnd_net_),
            .in1(N__44728),
            .in2(_gnd_net_),
            .in3(N__44698),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ),
            .ltout(),
            .carryin(bfn_18_9_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_9_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_9_1  (
            .in0(_gnd_net_),
            .in1(N__44695),
            .in2(_gnd_net_),
            .in3(N__44677),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_9_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_9_2  (
            .in0(_gnd_net_),
            .in1(N__44674),
            .in2(_gnd_net_),
            .in3(N__44656),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_9_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_9_3  (
            .in0(_gnd_net_),
            .in1(N__44653),
            .in2(_gnd_net_),
            .in3(N__44635),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_9_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_9_4  (
            .in0(_gnd_net_),
            .in1(N__44632),
            .in2(_gnd_net_),
            .in3(N__44614),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_9_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_9_5  (
            .in0(_gnd_net_),
            .in1(N__44611),
            .in2(_gnd_net_),
            .in3(N__44593),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_9_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_9_6  (
            .in0(_gnd_net_),
            .in1(N__44590),
            .in2(_gnd_net_),
            .in3(N__44572),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_9_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_9_7  (
            .in0(_gnd_net_),
            .in1(N__44944),
            .in2(_gnd_net_),
            .in3(N__44926),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_10_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(N__44923),
            .in2(_gnd_net_),
            .in3(N__44893),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_10_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_10_1  (
            .in0(_gnd_net_),
            .in1(N__44890),
            .in2(_gnd_net_),
            .in3(N__44872),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_10_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_10_2  (
            .in0(_gnd_net_),
            .in1(N__44869),
            .in2(_gnd_net_),
            .in3(N__44848),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_18_10_4 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_18_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_1_LC_18_10_4  (
            .in0(_gnd_net_),
            .in1(N__45759),
            .in2(_gnd_net_),
            .in3(N__45818),
            .lcout(\phase_controller_slave.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_1_LC_18_11_0 .C_ON=1'b0;
    defparam \phase_controller_slave.state_1_LC_18_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_1_LC_18_11_0 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_slave.state_1_LC_18_11_0  (
            .in0(N__44824),
            .in1(N__49035),
            .in2(N__44806),
            .in3(N__49013),
            .lcout(\phase_controller_slave.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48837),
            .ce(),
            .sr(N__48094));
    defparam \phase_controller_slave.S2_LC_18_11_4 .C_ON=1'b0;
    defparam \phase_controller_slave.S2_LC_18_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S2_LC_18_11_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \phase_controller_slave.S2_LC_18_11_4  (
            .in0(N__45757),
            .in1(N__49034),
            .in2(N__44766),
            .in3(N__45727),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48837),
            .ce(),
            .sr(N__48094));
    defparam \phase_controller_slave.state_0_LC_18_11_7 .C_ON=1'b0;
    defparam \phase_controller_slave.state_0_LC_18_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_0_LC_18_11_7 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_slave.state_0_LC_18_11_7  (
            .in0(N__49014),
            .in1(N__48971),
            .in2(N__49039),
            .in3(N__48948),
            .lcout(\phase_controller_slave.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48837),
            .ce(),
            .sr(N__48094));
    defparam \phase_controller_slave.start_timer_tr_LC_18_12_1 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_LC_18_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_tr_LC_18_12_1 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_slave.start_timer_tr_LC_18_12_1  (
            .in0(N__48985),
            .in1(N__45930),
            .in2(N__45603),
            .in3(N__48934),
            .lcout(\phase_controller_slave.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48828),
            .ce(),
            .sr(N__48100));
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_18_12_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_18_12_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_18_12_2  (
            .in0(N__45555),
            .in1(N__45460),
            .in2(_gnd_net_),
            .in3(N__45392),
            .lcout(),
            .ltout(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_18_12_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_18_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_18_12_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_LC_18_12_3  (
            .in0(N__48972),
            .in1(N__45904),
            .in2(N__45877),
            .in3(N__45874),
            .lcout(\phase_controller_slave.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48828),
            .ce(),
            .sr(N__48100));
    defparam \phase_controller_slave.state_3_LC_18_12_6 .C_ON=1'b0;
    defparam \phase_controller_slave.state_3_LC_18_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_3_LC_18_12_6 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \phase_controller_slave.state_3_LC_18_12_6  (
            .in0(N__48933),
            .in1(N__45758),
            .in2(N__45823),
            .in3(N__45796),
            .lcout(\phase_controller_slave.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48828),
            .ce(),
            .sr(N__48100));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_18_12_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_18_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_18_12_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_11_LC_18_12_7  (
            .in0(N__45393),
            .in1(N__45556),
            .in2(N__45498),
            .in3(N__45787),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48828),
            .ce(),
            .sr(N__48100));
    defparam \phase_controller_slave.S1_LC_18_13_0 .C_ON=1'b0;
    defparam \phase_controller_slave.S1_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S1_LC_18_13_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_slave.S1_LC_18_13_0  (
            .in0(N__45666),
            .in1(N__45756),
            .in2(_gnd_net_),
            .in3(N__45726),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48818),
            .ce(),
            .sr(N__48108));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_18_14_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_18_14_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_18_14_6  (
            .in0(N__45560),
            .in1(N__45459),
            .in2(_gnd_net_),
            .in3(N__45326),
            .lcout(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_18_15_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_18_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_18_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_16_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45274),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48800),
            .ce(N__45196),
            .sr(N__48123));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_17_6 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_18_17_6  (
            .in0(N__45137),
            .in1(N__45052),
            .in2(N__46559),
            .in3(N__44993),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48783),
            .ce(N__46644),
            .sr(N__48132));
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_18_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_18_18_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_18_18_7 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_4_LC_18_18_7  (
            .in0(N__46028),
            .in1(N__46526),
            .in2(N__46153),
            .in3(N__46439),
            .lcout(measured_delay_tr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48774),
            .ce(N__46349),
            .sr(N__48137));
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_18_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_18_19_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_18_19_5 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_2_LC_18_19_5  (
            .in0(N__46516),
            .in1(N__46473),
            .in2(N__46135),
            .in3(N__46438),
            .lcout(measured_delay_tr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48765),
            .ce(N__46344),
            .sr(N__48144));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_18_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_18_20_0 .LUT_INIT=16'b0000111100000010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_18_20_0  (
            .in0(N__47362),
            .in1(N__46269),
            .in2(N__49114),
            .in3(N__46251),
            .lcout(\delay_measurement_inst.N_286_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_18_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_18_20_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_18_20_6  (
            .in0(N__47168),
            .in1(N__47228),
            .in2(N__47118),
            .in3(N__47282),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_18_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_18_20_7 .LUT_INIT=16'b1101110111011100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_18_20_7  (
            .in0(N__46252),
            .in1(N__49099),
            .in2(N__46177),
            .in3(N__46174),
            .lcout(\delay_measurement_inst.N_373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_23_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_23_0  (
            .in0(_gnd_net_),
            .in1(N__48912),
            .in2(N__45993),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_18_23_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__48739),
            .ce(N__48346),
            .sr(N__48173));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_23_1  (
            .in0(_gnd_net_),
            .in1(N__46047),
            .in2(N__47040),
            .in3(N__45997),
            .lcout(\delay_measurement_inst.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__48739),
            .ce(N__48346),
            .sr(N__48173));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_23_2  (
            .in0(_gnd_net_),
            .in1(N__46991),
            .in2(N__45994),
            .in3(N__45940),
            .lcout(\delay_measurement_inst.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__48739),
            .ce(N__48346),
            .sr(N__48173));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_23_3  (
            .in0(_gnd_net_),
            .in1(N__46937),
            .in2(N__47041),
            .in3(N__46996),
            .lcout(\delay_measurement_inst.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__48739),
            .ce(N__48346),
            .sr(N__48173));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_23_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(N__46992),
            .in2(N__46884),
            .in3(N__46942),
            .lcout(\delay_measurement_inst.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__48739),
            .ce(N__48346),
            .sr(N__48173));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_23_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_23_5  (
            .in0(_gnd_net_),
            .in1(N__46938),
            .in2(N__46809),
            .in3(N__46888),
            .lcout(\delay_measurement_inst.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__48739),
            .ce(N__48346),
            .sr(N__48173));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_23_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_23_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_23_6  (
            .in0(_gnd_net_),
            .in1(N__46760),
            .in2(N__46885),
            .in3(N__46813),
            .lcout(\delay_measurement_inst.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__48739),
            .ce(N__48346),
            .sr(N__48173));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_23_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_23_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_23_7  (
            .in0(_gnd_net_),
            .in1(N__46712),
            .in2(N__46810),
            .in3(N__46765),
            .lcout(\delay_measurement_inst.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__48739),
            .ce(N__48346),
            .sr(N__48173));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_24_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_24_0  (
            .in0(_gnd_net_),
            .in1(N__46762),
            .in2(N__47502),
            .in3(N__46717),
            .lcout(\delay_measurement_inst.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_18_24_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__48734),
            .ce(N__48343),
            .sr(N__48186));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_24_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_24_1  (
            .in0(_gnd_net_),
            .in1(N__46714),
            .in2(N__47448),
            .in3(N__46669),
            .lcout(\delay_measurement_inst.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__48734),
            .ce(N__48343),
            .sr(N__48186));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_24_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_24_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_24_2  (
            .in0(_gnd_net_),
            .in1(N__47378),
            .in2(N__47503),
            .in3(N__47452),
            .lcout(\delay_measurement_inst.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__48734),
            .ce(N__48343),
            .sr(N__48186));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_24_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_24_3  (
            .in0(_gnd_net_),
            .in1(N__47306),
            .in2(N__47449),
            .in3(N__47383),
            .lcout(\delay_measurement_inst.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__48734),
            .ce(N__48343),
            .sr(N__48186));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_24_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_24_4  (
            .in0(_gnd_net_),
            .in1(N__47379),
            .in2(N__47253),
            .in3(N__47311),
            .lcout(\delay_measurement_inst.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__48734),
            .ce(N__48343),
            .sr(N__48186));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_24_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_24_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_24_5  (
            .in0(_gnd_net_),
            .in1(N__47307),
            .in2(N__47199),
            .in3(N__47257),
            .lcout(\delay_measurement_inst.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__48734),
            .ce(N__48343),
            .sr(N__48186));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_24_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_24_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_24_6  (
            .in0(_gnd_net_),
            .in1(N__47138),
            .in2(N__47254),
            .in3(N__47203),
            .lcout(\delay_measurement_inst.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__48734),
            .ce(N__48343),
            .sr(N__48186));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_24_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_24_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_24_7  (
            .in0(_gnd_net_),
            .in1(N__47072),
            .in2(N__47200),
            .in3(N__47143),
            .lcout(\delay_measurement_inst.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__48734),
            .ce(N__48343),
            .sr(N__48186));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_25_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_25_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_25_0  (
            .in0(_gnd_net_),
            .in1(N__47140),
            .in2(N__47772),
            .in3(N__47077),
            .lcout(\delay_measurement_inst.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_18_25_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__48727),
            .ce(N__48345),
            .sr(N__48194));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_25_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_25_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_25_1  (
            .in0(_gnd_net_),
            .in1(N__47074),
            .in2(N__47736),
            .in3(N__47044),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__48727),
            .ce(N__48345),
            .sr(N__48194));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_25_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_25_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_25_2  (
            .in0(_gnd_net_),
            .in1(N__47699),
            .in2(N__47773),
            .in3(N__47740),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__48727),
            .ce(N__48345),
            .sr(N__48194));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_25_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_25_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_25_3  (
            .in0(_gnd_net_),
            .in1(N__47669),
            .in2(N__47737),
            .in3(N__47704),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__48727),
            .ce(N__48345),
            .sr(N__48194));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_25_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_25_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_25_4  (
            .in0(_gnd_net_),
            .in1(N__47700),
            .in2(N__47637),
            .in3(N__47674),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__48727),
            .ce(N__48345),
            .sr(N__48194));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_25_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_25_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_25_5  (
            .in0(_gnd_net_),
            .in1(N__47670),
            .in2(N__47601),
            .in3(N__47641),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__48727),
            .ce(N__48345),
            .sr(N__48194));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_25_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_25_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_25_6  (
            .in0(_gnd_net_),
            .in1(N__47564),
            .in2(N__47638),
            .in3(N__47605),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__48727),
            .ce(N__48345),
            .sr(N__48194));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_25_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_25_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_25_7  (
            .in0(_gnd_net_),
            .in1(N__47534),
            .in2(N__47602),
            .in3(N__47569),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__48727),
            .ce(N__48345),
            .sr(N__48194));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_26_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_26_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_26_0  (
            .in0(_gnd_net_),
            .in1(N__47566),
            .in2(N__49212),
            .in3(N__47539),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_18_26_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__48720),
            .ce(N__48344),
            .sr(N__48201));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_26_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_26_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_26_1  (
            .in0(_gnd_net_),
            .in1(N__47536),
            .in2(N__49164),
            .in3(N__47506),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__48720),
            .ce(N__48344),
            .sr(N__48201));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_26_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_26_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_26_2  (
            .in0(_gnd_net_),
            .in1(N__49224),
            .in2(N__49213),
            .in3(N__49180),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__48720),
            .ce(N__48344),
            .sr(N__48201));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_26_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_26_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_26_3  (
            .in0(_gnd_net_),
            .in1(N__49176),
            .in2(N__49165),
            .in3(N__49132),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__48720),
            .ce(N__48344),
            .sr(N__48201));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_26_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_26_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49129),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48720),
            .ce(N__48344),
            .sr(N__48201));
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_20_11_6 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_20_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_tr_RNO_0_LC_20_11_6  (
            .in0(_gnd_net_),
            .in1(N__49033),
            .in2(_gnd_net_),
            .in3(N__49015),
            .lcout(\phase_controller_slave.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_20_12_5 .C_ON=1'b0;
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.state_RNIVDE2_0_LC_20_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.state_RNIVDE2_0_LC_20_12_5  (
            .in0(_gnd_net_),
            .in1(N__48973),
            .in2(_gnd_net_),
            .in3(N__48952),
            .lcout(\phase_controller_slave.N_211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48922),
            .lcout(\delay_measurement_inst.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48791),
            .ce(N__48339),
            .sr(N__48138));
endmodule // MAIN
