-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jul 15 2025 13:11:57

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__47202\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47108\ : std_logic;
signal \N__47101\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47035\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46718\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46496\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46493\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46223\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46130\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46103\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45143\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45068\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44951\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44511\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44380\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43989\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43706\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43443\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42673\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42541\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42332\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41681\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41051\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38746\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal pwm_duty_input_4 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal un7_start_stop_0_a3 : std_logic;
signal \N_34_i_i\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_94\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_94_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_120\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118_cascade_\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_53\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_3_10_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_3_11_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_enablelt3_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal un5_counter_cry_1 : std_logic;
signal un5_counter_cry_2 : std_logic;
signal un5_counter_cry_3 : std_logic;
signal un5_counter_cry_4 : std_logic;
signal un5_counter_cry_5 : std_logic;
signal un5_counter_cry_6 : std_logic;
signal un5_counter_cry_7 : std_logic;
signal un5_counter_cry_8 : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal un5_counter_cry_9 : std_logic;
signal un5_counter_cry_10 : std_logic;
signal un5_counter_cry_11 : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_4_6_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_4_7_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \current_shift_inst.PI_CTRL.N_170_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_168\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \counterZ0Z_11\ : std_logic;
signal \counterZ0Z_6\ : std_logic;
signal \counterZ0Z_12\ : std_logic;
signal \counterZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un2_counterZ0Z_1_cascade_\ : std_logic;
signal \counterZ0Z_8\ : std_logic;
signal \counterZ0Z_7\ : std_logic;
signal \counterZ0Z_9\ : std_logic;
signal \counterZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un2_counterZ0Z_8\ : std_logic;
signal \counterZ0Z_2\ : std_logic;
signal \counterZ0Z_3\ : std_logic;
signal \counterZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un2_counterZ0Z_7\ : std_logic;
signal \counterZ0Z_1\ : std_logic;
signal \counterZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un2_counterZ0\ : std_logic;
signal clk_10khz_i : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_167\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_171_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_170\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_171\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_0\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_1_cry_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_8\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_13\ : std_logic;
signal \current_shift_inst.control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_14\ : std_logic;
signal \current_shift_inst.control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_15\ : std_logic;
signal \current_shift_inst.control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_16\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_17\ : std_logic;
signal \current_shift_inst.control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_18\ : std_logic;
signal \current_shift_inst.control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_19\ : std_logic;
signal \current_shift_inst.control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_20\ : std_logic;
signal \current_shift_inst.control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_21\ : std_logic;
signal \current_shift_inst.control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_22\ : std_logic;
signal \current_shift_inst.control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_23\ : std_logic;
signal \current_shift_inst.control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_24\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_25\ : std_logic;
signal \N_748_g\ : std_logic;
signal \current_shift_inst.control_input_1_axb_23\ : std_logic;
signal il_max_comp1_c : std_logic;
signal il_min_comp2_c : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \current_shift_inst.control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.control_input_1_axb_3\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_0_sqmuxa\ : std_logic;
signal \current_shift_inst.control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.control_input_1_axb_0\ : std_logic;
signal \current_shift_inst.control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.control_input_1_axb_7\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_8\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_16\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_1_axb_25\ : std_logic;
signal s4_phy_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_8\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_16\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal s3_phy_c : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_10_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_10_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.N_1819_i\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input_0_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_463_i\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_257\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_257_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_240\ : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal state_ns_i_a3_1 : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.N_185_i\ : std_logic;
signal \delay_measurement_inst.prev_tr_sigZ0\ : std_logic;
signal \delay_measurement_inst.tr_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_RNO_0_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal measured_delay_tr_15 : std_logic;
signal measured_delay_tr_14 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.N_185_i_g\ : std_logic;
signal s1_phy_c : std_logic;
signal delay_tr_input_c : std_logic;
signal delay_tr_d1 : std_logic;
signal delay_tr_d2 : std_logic;
signal il_min_comp1_c : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\ : std_logic;
signal \delay_measurement_inst.N_360_cascade_\ : std_logic;
signal measured_delay_tr_9 : std_logic;
signal \delay_measurement_inst.N_354_cascade_\ : std_logic;
signal measured_delay_tr_10 : std_logic;
signal measured_delay_tr_11 : std_logic;
signal measured_delay_tr_12 : std_logic;
signal \delay_measurement_inst.N_354\ : std_logic;
signal measured_delay_tr_13 : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_186_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_14_27_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_14_28_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31_cascade_\ : std_logic;
signal measured_delay_tr_6 : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0\ : std_logic;
signal \delay_measurement_inst.N_381_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_376\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_\ : std_logic;
signal \delay_measurement_inst.N_498_cascade_\ : std_logic;
signal \delay_measurement_inst.N_381\ : std_logic;
signal \delay_measurement_inst.N_384\ : std_logic;
signal \delay_measurement_inst.N_384_cascade_\ : std_logic;
signal measured_delay_tr_4 : std_logic;
signal measured_delay_tr_5 : std_logic;
signal measured_delay_tr_7 : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31\ : std_logic;
signal measured_delay_tr_8 : std_logic;
signal measured_delay_tr_3 : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_RNOZ0Z_0_cascade_\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal state_3 : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal s2_phy_c : std_logic;
signal measured_delay_tr_1 : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg_5_tz_1\ : std_logic;
signal measured_delay_tr_2 : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_461_i_g\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_462_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \phase_controller_inst1.state_RNI7NN7Z0Z_0\ : std_logic;
signal \phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal measured_delay_tr_16 : std_logic;
signal measured_delay_tr_19 : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_6\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_373_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_3\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_11\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_19\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_16_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_316_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlt31_5_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_406\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_406_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_7_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2Z0Z_18\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_11\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_10\ : std_logic;
signal measured_delay_hc_24 : std_logic;
signal measured_delay_hc_23 : std_logic;
signal measured_delay_hc_22 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7Z0Z_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_299_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_2_6\ : std_logic;
signal \delay_measurement_inst.N_332_cascade_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_318_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_440\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_0_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_328_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_318_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_331\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_328\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_319\ : std_logic;
signal \delay_measurement_inst.N_318_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_6_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_7_6\ : std_logic;
signal measured_delay_hc_21 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0Z0Z_19\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_408\ : std_logic;
signal measured_delay_hc_26 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_17\ : std_logic;
signal measured_delay_hc_20 : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_461_i\ : std_logic;
signal delay_hc_input_c : std_logic;
signal delay_hc_d1 : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_464_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \delay_measurement_inst.hc_stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal delay_hc_d2 : std_logic;
signal \delay_measurement_inst.prev_hc_sigZ0\ : std_logic;
signal measured_delay_hc_8 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_1\ : std_logic;
signal measured_delay_hc_7 : std_logic;
signal measured_delay_hc_5 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_388\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_405_cascade_\ : std_logic;
signal measured_delay_hc_4 : std_logic;
signal measured_delay_hc_10 : std_logic;
signal measured_delay_hc_11 : std_logic;
signal measured_delay_hc_12 : std_logic;
signal measured_delay_hc_13 : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_459\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3\ : std_logic;
signal measured_delay_hc_3 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3_cascade_\ : std_logic;
signal measured_delay_hc_14 : std_logic;
signal \phase_controller_inst1.stoper_hc.N_405\ : std_logic;
signal measured_delay_hc_9 : std_logic;
signal measured_delay_hc_30 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6Z0Z_19\ : std_logic;
signal measured_delay_hc_6 : std_logic;
signal measured_delay_hc_29 : std_logic;
signal measured_delay_hc_27 : std_logic;
signal measured_delay_hc_28 : std_logic;
signal measured_delay_hc_0 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_19\ : std_logic;
signal measured_delay_hc_19 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_16\ : std_logic;
signal measured_delay_hc_1 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_18\ : std_logic;
signal measured_delay_hc_18 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_3\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto6\ : std_logic;
signal \delay_measurement_inst.N_332\ : std_logic;
signal \delay_measurement_inst.N_318\ : std_logic;
signal \delay_measurement_inst.N_295\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto15\ : std_logic;
signal measured_delay_hc_15 : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_463_i_g\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_17\ : std_logic;
signal measured_delay_tr_17 : std_logic;
signal \delay_measurement_inst.N_498\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_18\ : std_logic;
signal measured_delay_tr_18 : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal red_c_i : std_logic;
signal \phase_controller_inst2.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_453\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal measured_delay_hc_16 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_449\ : std_logic;
signal measured_delay_hc_31 : std_logic;
signal measured_delay_hc_17 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal measured_delay_hc_25 : std_logic;
signal \delay_measurement_inst.N_312\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.N_298\ : std_logic;
signal measured_delay_hc_2 : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__20197\&\N__20238\&\N__20195\&\N__20237\&\N__20196\&\N__20236\&\N__20198\&\N__20233\&\N__20191\&\N__20232\&\N__20192\&\N__20234\&\N__20193\&\N__20235\&\N__20194\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34373\&\N__34370\&'0'&'0'&'0'&\N__34368\&\N__34372\&\N__34369\&\N__34371\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__20261\&\N__20278\&\N__20262\&\N__20279\&\N__20263\&\N__18851\&\N__17877\&\N__17934\&\N__17952\&\N__17916\&\N__17898\&\N__17853\&\N__33170\&\N__33227\&\N__33200\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34564\&\N__34561\&'0'&'0'&'0'&\N__34559\&\N__34563\&\N__34560\&\N__34562\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__18576\,
            RESETB => \N__42506\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__34374\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__34367\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__34565\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__34558\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__47200\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47202\,
            DIN => \N__47201\,
            DOUT => \N__47200\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47202\,
            PADOUT => \N__47201\,
            PADIN => \N__47200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47191\,
            DIN => \N__47190\,
            DOUT => \N__47189\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47191\,
            PADOUT => \N__47190\,
            PADIN => \N__47189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47182\,
            DIN => \N__47181\,
            DOUT => \N__47180\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47182\,
            PADOUT => \N__47181\,
            PADIN => \N__47180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47173\,
            DIN => \N__47172\,
            DOUT => \N__47171\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47173\,
            PADOUT => \N__47172\,
            PADIN => \N__47171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21351\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47164\,
            DIN => \N__47163\,
            DOUT => \N__47162\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47164\,
            PADOUT => \N__47163\,
            PADIN => \N__47162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47155\,
            DIN => \N__47154\,
            DOUT => \N__47153\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47155\,
            PADOUT => \N__47154\,
            PADIN => \N__47153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36021\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47146\,
            DIN => \N__47145\,
            DOUT => \N__47144\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47146\,
            PADOUT => \N__47145\,
            PADIN => \N__47144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47137\,
            DIN => \N__47136\,
            DOUT => \N__47135\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47137\,
            PADOUT => \N__47136\,
            PADIN => \N__47135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47128\,
            DIN => \N__47127\,
            DOUT => \N__47126\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47128\,
            PADOUT => \N__47127\,
            PADIN => \N__47126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47119\,
            DIN => \N__47118\,
            DOUT => \N__47117\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47119\,
            PADOUT => \N__47118\,
            PADIN => \N__47117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33021\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47110\,
            DIN => \N__47109\,
            DOUT => \N__47108\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47110\,
            PADOUT => \N__47109\,
            PADIN => \N__47108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25611\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47101\,
            DIN => \N__47100\,
            DOUT => \N__47099\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47101\,
            PADOUT => \N__47100\,
            PADIN => \N__47099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47092\,
            DIN => \N__47091\,
            DOUT => \N__47090\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47092\,
            PADOUT => \N__47091\,
            PADIN => \N__47090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26148\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11252\ : InMux
    port map (
            O => \N__47073\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__11251\ : InMux
    port map (
            O => \N__47070\,
            I => \N__47066\
        );

    \I__11250\ : InMux
    port map (
            O => \N__47069\,
            I => \N__47063\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__47066\,
            I => \N__47056\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__47063\,
            I => \N__47053\
        );

    \I__11247\ : InMux
    port map (
            O => \N__47062\,
            I => \N__47044\
        );

    \I__11246\ : InMux
    port map (
            O => \N__47061\,
            I => \N__47044\
        );

    \I__11245\ : InMux
    port map (
            O => \N__47060\,
            I => \N__47044\
        );

    \I__11244\ : InMux
    port map (
            O => \N__47059\,
            I => \N__47044\
        );

    \I__11243\ : Span4Mux_v
    port map (
            O => \N__47056\,
            I => \N__47041\
        );

    \I__11242\ : Span12Mux_v
    port map (
            O => \N__47053\,
            I => \N__47038\
        );

    \I__11241\ : LocalMux
    port map (
            O => \N__47044\,
            I => \N__47035\
        );

    \I__11240\ : Odrv4
    port map (
            O => \N__47041\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__11239\ : Odrv12
    port map (
            O => \N__47038\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__11238\ : Odrv12
    port map (
            O => \N__47035\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__11237\ : InMux
    port map (
            O => \N__47028\,
            I => \N__47025\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__47025\,
            I => \N__47022\
        );

    \I__11235\ : Span4Mux_h
    port map (
            O => \N__47022\,
            I => \N__47017\
        );

    \I__11234\ : InMux
    port map (
            O => \N__47021\,
            I => \N__47014\
        );

    \I__11233\ : InMux
    port map (
            O => \N__47020\,
            I => \N__47011\
        );

    \I__11232\ : Odrv4
    port map (
            O => \N__47017\,
            I => \phase_controller_inst1.stoper_hc.N_453\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__47014\,
            I => \phase_controller_inst1.stoper_hc.N_453\
        );

    \I__11230\ : LocalMux
    port map (
            O => \N__47011\,
            I => \phase_controller_inst1.stoper_hc.N_453\
        );

    \I__11229\ : CascadeMux
    port map (
            O => \N__47004\,
            I => \N__47001\
        );

    \I__11228\ : InMux
    port map (
            O => \N__47001\,
            I => \N__46998\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__46998\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__11226\ : InMux
    port map (
            O => \N__46995\,
            I => \N__46991\
        );

    \I__11225\ : CascadeMux
    port map (
            O => \N__46994\,
            I => \N__46988\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__46991\,
            I => \N__46985\
        );

    \I__11223\ : InMux
    port map (
            O => \N__46988\,
            I => \N__46979\
        );

    \I__11222\ : Span4Mux_h
    port map (
            O => \N__46985\,
            I => \N__46976\
        );

    \I__11221\ : InMux
    port map (
            O => \N__46984\,
            I => \N__46973\
        );

    \I__11220\ : InMux
    port map (
            O => \N__46983\,
            I => \N__46970\
        );

    \I__11219\ : InMux
    port map (
            O => \N__46982\,
            I => \N__46967\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__46979\,
            I => measured_delay_hc_16
        );

    \I__11217\ : Odrv4
    port map (
            O => \N__46976\,
            I => measured_delay_hc_16
        );

    \I__11216\ : LocalMux
    port map (
            O => \N__46973\,
            I => measured_delay_hc_16
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__46970\,
            I => measured_delay_hc_16
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__46967\,
            I => measured_delay_hc_16
        );

    \I__11213\ : CascadeMux
    port map (
            O => \N__46956\,
            I => \N__46953\
        );

    \I__11212\ : InMux
    port map (
            O => \N__46953\,
            I => \N__46950\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__46950\,
            I => \N__46947\
        );

    \I__11210\ : Odrv4
    port map (
            O => \N__46947\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__11209\ : CascadeMux
    port map (
            O => \N__46944\,
            I => \N__46931\
        );

    \I__11208\ : CascadeMux
    port map (
            O => \N__46943\,
            I => \N__46928\
        );

    \I__11207\ : CascadeMux
    port map (
            O => \N__46942\,
            I => \N__46925\
        );

    \I__11206\ : CascadeMux
    port map (
            O => \N__46941\,
            I => \N__46922\
        );

    \I__11205\ : InMux
    port map (
            O => \N__46940\,
            I => \N__46896\
        );

    \I__11204\ : InMux
    port map (
            O => \N__46939\,
            I => \N__46896\
        );

    \I__11203\ : InMux
    port map (
            O => \N__46938\,
            I => \N__46896\
        );

    \I__11202\ : InMux
    port map (
            O => \N__46937\,
            I => \N__46896\
        );

    \I__11201\ : InMux
    port map (
            O => \N__46936\,
            I => \N__46896\
        );

    \I__11200\ : InMux
    port map (
            O => \N__46935\,
            I => \N__46896\
        );

    \I__11199\ : InMux
    port map (
            O => \N__46934\,
            I => \N__46893\
        );

    \I__11198\ : InMux
    port map (
            O => \N__46931\,
            I => \N__46873\
        );

    \I__11197\ : InMux
    port map (
            O => \N__46928\,
            I => \N__46873\
        );

    \I__11196\ : InMux
    port map (
            O => \N__46925\,
            I => \N__46873\
        );

    \I__11195\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46873\
        );

    \I__11194\ : InMux
    port map (
            O => \N__46921\,
            I => \N__46873\
        );

    \I__11193\ : InMux
    port map (
            O => \N__46920\,
            I => \N__46873\
        );

    \I__11192\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46873\
        );

    \I__11191\ : InMux
    port map (
            O => \N__46918\,
            I => \N__46873\
        );

    \I__11190\ : InMux
    port map (
            O => \N__46917\,
            I => \N__46868\
        );

    \I__11189\ : InMux
    port map (
            O => \N__46916\,
            I => \N__46868\
        );

    \I__11188\ : InMux
    port map (
            O => \N__46915\,
            I => \N__46853\
        );

    \I__11187\ : InMux
    port map (
            O => \N__46914\,
            I => \N__46853\
        );

    \I__11186\ : InMux
    port map (
            O => \N__46913\,
            I => \N__46853\
        );

    \I__11185\ : InMux
    port map (
            O => \N__46912\,
            I => \N__46853\
        );

    \I__11184\ : InMux
    port map (
            O => \N__46911\,
            I => \N__46853\
        );

    \I__11183\ : InMux
    port map (
            O => \N__46910\,
            I => \N__46853\
        );

    \I__11182\ : InMux
    port map (
            O => \N__46909\,
            I => \N__46853\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__46896\,
            I => \N__46850\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__46893\,
            I => \N__46847\
        );

    \I__11179\ : InMux
    port map (
            O => \N__46892\,
            I => \N__46837\
        );

    \I__11178\ : InMux
    port map (
            O => \N__46891\,
            I => \N__46837\
        );

    \I__11177\ : InMux
    port map (
            O => \N__46890\,
            I => \N__46837\
        );

    \I__11176\ : LocalMux
    port map (
            O => \N__46873\,
            I => \N__46825\
        );

    \I__11175\ : LocalMux
    port map (
            O => \N__46868\,
            I => \N__46822\
        );

    \I__11174\ : LocalMux
    port map (
            O => \N__46853\,
            I => \N__46815\
        );

    \I__11173\ : Span4Mux_h
    port map (
            O => \N__46850\,
            I => \N__46815\
        );

    \I__11172\ : Span4Mux_h
    port map (
            O => \N__46847\,
            I => \N__46815\
        );

    \I__11171\ : InMux
    port map (
            O => \N__46846\,
            I => \N__46808\
        );

    \I__11170\ : InMux
    port map (
            O => \N__46845\,
            I => \N__46808\
        );

    \I__11169\ : InMux
    port map (
            O => \N__46844\,
            I => \N__46808\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__46837\,
            I => \N__46805\
        );

    \I__11167\ : InMux
    port map (
            O => \N__46836\,
            I => \N__46792\
        );

    \I__11166\ : InMux
    port map (
            O => \N__46835\,
            I => \N__46792\
        );

    \I__11165\ : InMux
    port map (
            O => \N__46834\,
            I => \N__46792\
        );

    \I__11164\ : InMux
    port map (
            O => \N__46833\,
            I => \N__46792\
        );

    \I__11163\ : InMux
    port map (
            O => \N__46832\,
            I => \N__46792\
        );

    \I__11162\ : InMux
    port map (
            O => \N__46831\,
            I => \N__46792\
        );

    \I__11161\ : InMux
    port map (
            O => \N__46830\,
            I => \N__46784\
        );

    \I__11160\ : InMux
    port map (
            O => \N__46829\,
            I => \N__46784\
        );

    \I__11159\ : InMux
    port map (
            O => \N__46828\,
            I => \N__46784\
        );

    \I__11158\ : Span4Mux_v
    port map (
            O => \N__46825\,
            I => \N__46781\
        );

    \I__11157\ : Span4Mux_h
    port map (
            O => \N__46822\,
            I => \N__46776\
        );

    \I__11156\ : Span4Mux_v
    port map (
            O => \N__46815\,
            I => \N__46776\
        );

    \I__11155\ : LocalMux
    port map (
            O => \N__46808\,
            I => \N__46769\
        );

    \I__11154\ : Span4Mux_h
    port map (
            O => \N__46805\,
            I => \N__46769\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__46792\,
            I => \N__46769\
        );

    \I__11152\ : InMux
    port map (
            O => \N__46791\,
            I => \N__46766\
        );

    \I__11151\ : LocalMux
    port map (
            O => \N__46784\,
            I => \phase_controller_inst1.stoper_hc.N_449\
        );

    \I__11150\ : Odrv4
    port map (
            O => \N__46781\,
            I => \phase_controller_inst1.stoper_hc.N_449\
        );

    \I__11149\ : Odrv4
    port map (
            O => \N__46776\,
            I => \phase_controller_inst1.stoper_hc.N_449\
        );

    \I__11148\ : Odrv4
    port map (
            O => \N__46769\,
            I => \phase_controller_inst1.stoper_hc.N_449\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__46766\,
            I => \phase_controller_inst1.stoper_hc.N_449\
        );

    \I__11146\ : CascadeMux
    port map (
            O => \N__46755\,
            I => \N__46751\
        );

    \I__11145\ : InMux
    port map (
            O => \N__46754\,
            I => \N__46748\
        );

    \I__11144\ : InMux
    port map (
            O => \N__46751\,
            I => \N__46743\
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__46748\,
            I => \N__46740\
        );

    \I__11142\ : InMux
    port map (
            O => \N__46747\,
            I => \N__46735\
        );

    \I__11141\ : InMux
    port map (
            O => \N__46746\,
            I => \N__46735\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__46743\,
            I => \N__46726\
        );

    \I__11139\ : Span4Mux_v
    port map (
            O => \N__46740\,
            I => \N__46721\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__46735\,
            I => \N__46721\
        );

    \I__11137\ : CascadeMux
    port map (
            O => \N__46734\,
            I => \N__46718\
        );

    \I__11136\ : InMux
    port map (
            O => \N__46733\,
            I => \N__46703\
        );

    \I__11135\ : InMux
    port map (
            O => \N__46732\,
            I => \N__46703\
        );

    \I__11134\ : InMux
    port map (
            O => \N__46731\,
            I => \N__46703\
        );

    \I__11133\ : InMux
    port map (
            O => \N__46730\,
            I => \N__46703\
        );

    \I__11132\ : InMux
    port map (
            O => \N__46729\,
            I => \N__46698\
        );

    \I__11131\ : Span4Mux_v
    port map (
            O => \N__46726\,
            I => \N__46693\
        );

    \I__11130\ : Span4Mux_h
    port map (
            O => \N__46721\,
            I => \N__46693\
        );

    \I__11129\ : InMux
    port map (
            O => \N__46718\,
            I => \N__46686\
        );

    \I__11128\ : InMux
    port map (
            O => \N__46717\,
            I => \N__46686\
        );

    \I__11127\ : InMux
    port map (
            O => \N__46716\,
            I => \N__46686\
        );

    \I__11126\ : InMux
    port map (
            O => \N__46715\,
            I => \N__46681\
        );

    \I__11125\ : InMux
    port map (
            O => \N__46714\,
            I => \N__46681\
        );

    \I__11124\ : InMux
    port map (
            O => \N__46713\,
            I => \N__46678\
        );

    \I__11123\ : InMux
    port map (
            O => \N__46712\,
            I => \N__46675\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__46703\,
            I => \N__46672\
        );

    \I__11121\ : InMux
    port map (
            O => \N__46702\,
            I => \N__46667\
        );

    \I__11120\ : InMux
    port map (
            O => \N__46701\,
            I => \N__46667\
        );

    \I__11119\ : LocalMux
    port map (
            O => \N__46698\,
            I => \N__46664\
        );

    \I__11118\ : Odrv4
    port map (
            O => \N__46693\,
            I => measured_delay_hc_31
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__46686\,
            I => measured_delay_hc_31
        );

    \I__11116\ : LocalMux
    port map (
            O => \N__46681\,
            I => measured_delay_hc_31
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__46678\,
            I => measured_delay_hc_31
        );

    \I__11114\ : LocalMux
    port map (
            O => \N__46675\,
            I => measured_delay_hc_31
        );

    \I__11113\ : Odrv4
    port map (
            O => \N__46672\,
            I => measured_delay_hc_31
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__46667\,
            I => measured_delay_hc_31
        );

    \I__11111\ : Odrv4
    port map (
            O => \N__46664\,
            I => measured_delay_hc_31
        );

    \I__11110\ : InMux
    port map (
            O => \N__46647\,
            I => \N__46644\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__46644\,
            I => \N__46638\
        );

    \I__11108\ : InMux
    port map (
            O => \N__46643\,
            I => \N__46634\
        );

    \I__11107\ : InMux
    port map (
            O => \N__46642\,
            I => \N__46631\
        );

    \I__11106\ : CascadeMux
    port map (
            O => \N__46641\,
            I => \N__46628\
        );

    \I__11105\ : Span4Mux_h
    port map (
            O => \N__46638\,
            I => \N__46625\
        );

    \I__11104\ : InMux
    port map (
            O => \N__46637\,
            I => \N__46622\
        );

    \I__11103\ : LocalMux
    port map (
            O => \N__46634\,
            I => \N__46619\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__46631\,
            I => \N__46616\
        );

    \I__11101\ : InMux
    port map (
            O => \N__46628\,
            I => \N__46613\
        );

    \I__11100\ : Span4Mux_v
    port map (
            O => \N__46625\,
            I => \N__46610\
        );

    \I__11099\ : LocalMux
    port map (
            O => \N__46622\,
            I => \N__46607\
        );

    \I__11098\ : Span4Mux_v
    port map (
            O => \N__46619\,
            I => \N__46602\
        );

    \I__11097\ : Span4Mux_h
    port map (
            O => \N__46616\,
            I => \N__46602\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__46613\,
            I => measured_delay_hc_17
        );

    \I__11095\ : Odrv4
    port map (
            O => \N__46610\,
            I => measured_delay_hc_17
        );

    \I__11094\ : Odrv12
    port map (
            O => \N__46607\,
            I => measured_delay_hc_17
        );

    \I__11093\ : Odrv4
    port map (
            O => \N__46602\,
            I => measured_delay_hc_17
        );

    \I__11092\ : CascadeMux
    port map (
            O => \N__46593\,
            I => \N__46590\
        );

    \I__11091\ : InMux
    port map (
            O => \N__46590\,
            I => \N__46587\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__46587\,
            I => \N__46584\
        );

    \I__11089\ : Odrv4
    port map (
            O => \N__46584\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__11088\ : CEMux
    port map (
            O => \N__46581\,
            I => \N__46574\
        );

    \I__11087\ : CEMux
    port map (
            O => \N__46580\,
            I => \N__46571\
        );

    \I__11086\ : CEMux
    port map (
            O => \N__46579\,
            I => \N__46568\
        );

    \I__11085\ : CEMux
    port map (
            O => \N__46578\,
            I => \N__46565\
        );

    \I__11084\ : CEMux
    port map (
            O => \N__46577\,
            I => \N__46562\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__46574\,
            I => \N__46558\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__46571\,
            I => \N__46555\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__46568\,
            I => \N__46552\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__46565\,
            I => \N__46549\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__46562\,
            I => \N__46546\
        );

    \I__11078\ : CEMux
    port map (
            O => \N__46561\,
            I => \N__46543\
        );

    \I__11077\ : Span4Mux_v
    port map (
            O => \N__46558\,
            I => \N__46540\
        );

    \I__11076\ : Span4Mux_v
    port map (
            O => \N__46555\,
            I => \N__46535\
        );

    \I__11075\ : Span4Mux_h
    port map (
            O => \N__46552\,
            I => \N__46535\
        );

    \I__11074\ : Span4Mux_v
    port map (
            O => \N__46549\,
            I => \N__46528\
        );

    \I__11073\ : Span4Mux_h
    port map (
            O => \N__46546\,
            I => \N__46528\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__46543\,
            I => \N__46528\
        );

    \I__11071\ : Span4Mux_h
    port map (
            O => \N__46540\,
            I => \N__46523\
        );

    \I__11070\ : Span4Mux_h
    port map (
            O => \N__46535\,
            I => \N__46523\
        );

    \I__11069\ : Span4Mux_v
    port map (
            O => \N__46528\,
            I => \N__46520\
        );

    \I__11068\ : Odrv4
    port map (
            O => \N__46523\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__11067\ : Odrv4
    port map (
            O => \N__46520\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__11066\ : InMux
    port map (
            O => \N__46515\,
            I => \N__46511\
        );

    \I__11065\ : InMux
    port map (
            O => \N__46514\,
            I => \N__46508\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__46511\,
            I => \N__46505\
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__46508\,
            I => measured_delay_hc_25
        );

    \I__11062\ : Odrv4
    port map (
            O => \N__46505\,
            I => measured_delay_hc_25
        );

    \I__11061\ : CascadeMux
    port map (
            O => \N__46500\,
            I => \N__46488\
        );

    \I__11060\ : CascadeMux
    port map (
            O => \N__46499\,
            I => \N__46485\
        );

    \I__11059\ : CascadeMux
    port map (
            O => \N__46498\,
            I => \N__46478\
        );

    \I__11058\ : CascadeMux
    port map (
            O => \N__46497\,
            I => \N__46475\
        );

    \I__11057\ : CascadeMux
    port map (
            O => \N__46496\,
            I => \N__46470\
        );

    \I__11056\ : CascadeMux
    port map (
            O => \N__46495\,
            I => \N__46466\
        );

    \I__11055\ : CascadeMux
    port map (
            O => \N__46494\,
            I => \N__46462\
        );

    \I__11054\ : CascadeMux
    port map (
            O => \N__46493\,
            I => \N__46456\
        );

    \I__11053\ : CascadeMux
    port map (
            O => \N__46492\,
            I => \N__46453\
        );

    \I__11052\ : InMux
    port map (
            O => \N__46491\,
            I => \N__46440\
        );

    \I__11051\ : InMux
    port map (
            O => \N__46488\,
            I => \N__46440\
        );

    \I__11050\ : InMux
    port map (
            O => \N__46485\,
            I => \N__46440\
        );

    \I__11049\ : InMux
    port map (
            O => \N__46484\,
            I => \N__46440\
        );

    \I__11048\ : InMux
    port map (
            O => \N__46483\,
            I => \N__46434\
        );

    \I__11047\ : InMux
    port map (
            O => \N__46482\,
            I => \N__46434\
        );

    \I__11046\ : InMux
    port map (
            O => \N__46481\,
            I => \N__46423\
        );

    \I__11045\ : InMux
    port map (
            O => \N__46478\,
            I => \N__46423\
        );

    \I__11044\ : InMux
    port map (
            O => \N__46475\,
            I => \N__46423\
        );

    \I__11043\ : InMux
    port map (
            O => \N__46474\,
            I => \N__46423\
        );

    \I__11042\ : InMux
    port map (
            O => \N__46473\,
            I => \N__46423\
        );

    \I__11041\ : InMux
    port map (
            O => \N__46470\,
            I => \N__46414\
        );

    \I__11040\ : InMux
    port map (
            O => \N__46469\,
            I => \N__46414\
        );

    \I__11039\ : InMux
    port map (
            O => \N__46466\,
            I => \N__46414\
        );

    \I__11038\ : InMux
    port map (
            O => \N__46465\,
            I => \N__46414\
        );

    \I__11037\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46409\
        );

    \I__11036\ : InMux
    port map (
            O => \N__46461\,
            I => \N__46409\
        );

    \I__11035\ : InMux
    port map (
            O => \N__46460\,
            I => \N__46406\
        );

    \I__11034\ : InMux
    port map (
            O => \N__46459\,
            I => \N__46395\
        );

    \I__11033\ : InMux
    port map (
            O => \N__46456\,
            I => \N__46395\
        );

    \I__11032\ : InMux
    port map (
            O => \N__46453\,
            I => \N__46395\
        );

    \I__11031\ : InMux
    port map (
            O => \N__46452\,
            I => \N__46395\
        );

    \I__11030\ : InMux
    port map (
            O => \N__46451\,
            I => \N__46395\
        );

    \I__11029\ : CascadeMux
    port map (
            O => \N__46450\,
            I => \N__46392\
        );

    \I__11028\ : CascadeMux
    port map (
            O => \N__46449\,
            I => \N__46389\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__46440\,
            I => \N__46384\
        );

    \I__11026\ : InMux
    port map (
            O => \N__46439\,
            I => \N__46381\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__46434\,
            I => \N__46375\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__46423\,
            I => \N__46370\
        );

    \I__11023\ : LocalMux
    port map (
            O => \N__46414\,
            I => \N__46370\
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__46409\,
            I => \N__46367\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__46406\,
            I => \N__46362\
        );

    \I__11020\ : LocalMux
    port map (
            O => \N__46395\,
            I => \N__46362\
        );

    \I__11019\ : InMux
    port map (
            O => \N__46392\,
            I => \N__46353\
        );

    \I__11018\ : InMux
    port map (
            O => \N__46389\,
            I => \N__46353\
        );

    \I__11017\ : InMux
    port map (
            O => \N__46388\,
            I => \N__46353\
        );

    \I__11016\ : InMux
    port map (
            O => \N__46387\,
            I => \N__46353\
        );

    \I__11015\ : Span4Mux_v
    port map (
            O => \N__46384\,
            I => \N__46347\
        );

    \I__11014\ : LocalMux
    port map (
            O => \N__46381\,
            I => \N__46347\
        );

    \I__11013\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46340\
        );

    \I__11012\ : InMux
    port map (
            O => \N__46379\,
            I => \N__46340\
        );

    \I__11011\ : InMux
    port map (
            O => \N__46378\,
            I => \N__46340\
        );

    \I__11010\ : Span4Mux_h
    port map (
            O => \N__46375\,
            I => \N__46335\
        );

    \I__11009\ : Span4Mux_h
    port map (
            O => \N__46370\,
            I => \N__46335\
        );

    \I__11008\ : Span4Mux_v
    port map (
            O => \N__46367\,
            I => \N__46328\
        );

    \I__11007\ : Span4Mux_h
    port map (
            O => \N__46362\,
            I => \N__46328\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__46353\,
            I => \N__46328\
        );

    \I__11005\ : InMux
    port map (
            O => \N__46352\,
            I => \N__46325\
        );

    \I__11004\ : Span4Mux_v
    port map (
            O => \N__46347\,
            I => \N__46320\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__46340\,
            I => \N__46320\
        );

    \I__11002\ : Odrv4
    port map (
            O => \N__46335\,
            I => \delay_measurement_inst.N_312\
        );

    \I__11001\ : Odrv4
    port map (
            O => \N__46328\,
            I => \delay_measurement_inst.N_312\
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__46325\,
            I => \delay_measurement_inst.N_312\
        );

    \I__10999\ : Odrv4
    port map (
            O => \N__46320\,
            I => \delay_measurement_inst.N_312\
        );

    \I__10998\ : CascadeMux
    port map (
            O => \N__46311\,
            I => \N__46308\
        );

    \I__10997\ : InMux
    port map (
            O => \N__46308\,
            I => \N__46305\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__46305\,
            I => \N__46301\
        );

    \I__10995\ : InMux
    port map (
            O => \N__46304\,
            I => \N__46298\
        );

    \I__10994\ : Span4Mux_v
    port map (
            O => \N__46301\,
            I => \N__46293\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__46298\,
            I => \N__46293\
        );

    \I__10992\ : Span4Mux_h
    port map (
            O => \N__46293\,
            I => \N__46289\
        );

    \I__10991\ : InMux
    port map (
            O => \N__46292\,
            I => \N__46286\
        );

    \I__10990\ : Odrv4
    port map (
            O => \N__46289\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__46286\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__10988\ : InMux
    port map (
            O => \N__46281\,
            I => \N__46256\
        );

    \I__10987\ : InMux
    port map (
            O => \N__46280\,
            I => \N__46256\
        );

    \I__10986\ : InMux
    port map (
            O => \N__46279\,
            I => \N__46256\
        );

    \I__10985\ : InMux
    port map (
            O => \N__46278\,
            I => \N__46256\
        );

    \I__10984\ : InMux
    port map (
            O => \N__46277\,
            I => \N__46243\
        );

    \I__10983\ : InMux
    port map (
            O => \N__46276\,
            I => \N__46243\
        );

    \I__10982\ : InMux
    port map (
            O => \N__46275\,
            I => \N__46232\
        );

    \I__10981\ : InMux
    port map (
            O => \N__46274\,
            I => \N__46232\
        );

    \I__10980\ : InMux
    port map (
            O => \N__46273\,
            I => \N__46232\
        );

    \I__10979\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46232\
        );

    \I__10978\ : InMux
    port map (
            O => \N__46271\,
            I => \N__46232\
        );

    \I__10977\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46223\
        );

    \I__10976\ : InMux
    port map (
            O => \N__46269\,
            I => \N__46223\
        );

    \I__10975\ : InMux
    port map (
            O => \N__46268\,
            I => \N__46223\
        );

    \I__10974\ : InMux
    port map (
            O => \N__46267\,
            I => \N__46223\
        );

    \I__10973\ : InMux
    port map (
            O => \N__46266\,
            I => \N__46215\
        );

    \I__10972\ : InMux
    port map (
            O => \N__46265\,
            I => \N__46215\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__46256\,
            I => \N__46212\
        );

    \I__10970\ : InMux
    port map (
            O => \N__46255\,
            I => \N__46209\
        );

    \I__10969\ : InMux
    port map (
            O => \N__46254\,
            I => \N__46206\
        );

    \I__10968\ : InMux
    port map (
            O => \N__46253\,
            I => \N__46193\
        );

    \I__10967\ : InMux
    port map (
            O => \N__46252\,
            I => \N__46193\
        );

    \I__10966\ : InMux
    port map (
            O => \N__46251\,
            I => \N__46193\
        );

    \I__10965\ : InMux
    port map (
            O => \N__46250\,
            I => \N__46193\
        );

    \I__10964\ : InMux
    port map (
            O => \N__46249\,
            I => \N__46193\
        );

    \I__10963\ : InMux
    port map (
            O => \N__46248\,
            I => \N__46193\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__46243\,
            I => \N__46190\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__46232\,
            I => \N__46185\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__46223\,
            I => \N__46185\
        );

    \I__10959\ : InMux
    port map (
            O => \N__46222\,
            I => \N__46178\
        );

    \I__10958\ : InMux
    port map (
            O => \N__46221\,
            I => \N__46178\
        );

    \I__10957\ : InMux
    port map (
            O => \N__46220\,
            I => \N__46178\
        );

    \I__10956\ : LocalMux
    port map (
            O => \N__46215\,
            I => \N__46171\
        );

    \I__10955\ : Span4Mux_v
    port map (
            O => \N__46212\,
            I => \N__46166\
        );

    \I__10954\ : LocalMux
    port map (
            O => \N__46209\,
            I => \N__46166\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__46206\,
            I => \N__46163\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__46193\,
            I => \N__46160\
        );

    \I__10951\ : Span4Mux_h
    port map (
            O => \N__46190\,
            I => \N__46153\
        );

    \I__10950\ : Span4Mux_h
    port map (
            O => \N__46185\,
            I => \N__46153\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__46178\,
            I => \N__46153\
        );

    \I__10948\ : InMux
    port map (
            O => \N__46177\,
            I => \N__46144\
        );

    \I__10947\ : InMux
    port map (
            O => \N__46176\,
            I => \N__46144\
        );

    \I__10946\ : InMux
    port map (
            O => \N__46175\,
            I => \N__46144\
        );

    \I__10945\ : InMux
    port map (
            O => \N__46174\,
            I => \N__46144\
        );

    \I__10944\ : Odrv12
    port map (
            O => \N__46171\,
            I => \delay_measurement_inst.N_298\
        );

    \I__10943\ : Odrv4
    port map (
            O => \N__46166\,
            I => \delay_measurement_inst.N_298\
        );

    \I__10942\ : Odrv4
    port map (
            O => \N__46163\,
            I => \delay_measurement_inst.N_298\
        );

    \I__10941\ : Odrv4
    port map (
            O => \N__46160\,
            I => \delay_measurement_inst.N_298\
        );

    \I__10940\ : Odrv4
    port map (
            O => \N__46153\,
            I => \delay_measurement_inst.N_298\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__46144\,
            I => \delay_measurement_inst.N_298\
        );

    \I__10938\ : InMux
    port map (
            O => \N__46131\,
            I => \N__46125\
        );

    \I__10937\ : InMux
    port map (
            O => \N__46130\,
            I => \N__46122\
        );

    \I__10936\ : InMux
    port map (
            O => \N__46129\,
            I => \N__46119\
        );

    \I__10935\ : InMux
    port map (
            O => \N__46128\,
            I => \N__46116\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__46125\,
            I => \N__46113\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__46122\,
            I => \N__46109\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__46119\,
            I => \N__46106\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__46116\,
            I => \N__46103\
        );

    \I__10930\ : Span4Mux_h
    port map (
            O => \N__46113\,
            I => \N__46100\
        );

    \I__10929\ : InMux
    port map (
            O => \N__46112\,
            I => \N__46097\
        );

    \I__10928\ : Span4Mux_v
    port map (
            O => \N__46109\,
            I => \N__46094\
        );

    \I__10927\ : Span4Mux_h
    port map (
            O => \N__46106\,
            I => \N__46091\
        );

    \I__10926\ : Span4Mux_v
    port map (
            O => \N__46103\,
            I => \N__46086\
        );

    \I__10925\ : Span4Mux_v
    port map (
            O => \N__46100\,
            I => \N__46086\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__46097\,
            I => measured_delay_hc_2
        );

    \I__10923\ : Odrv4
    port map (
            O => \N__46094\,
            I => measured_delay_hc_2
        );

    \I__10922\ : Odrv4
    port map (
            O => \N__46091\,
            I => measured_delay_hc_2
        );

    \I__10921\ : Odrv4
    port map (
            O => \N__46086\,
            I => measured_delay_hc_2
        );

    \I__10920\ : ClkMux
    port map (
            O => \N__46077\,
            I => \N__45627\
        );

    \I__10919\ : ClkMux
    port map (
            O => \N__46076\,
            I => \N__45627\
        );

    \I__10918\ : ClkMux
    port map (
            O => \N__46075\,
            I => \N__45627\
        );

    \I__10917\ : ClkMux
    port map (
            O => \N__46074\,
            I => \N__45627\
        );

    \I__10916\ : ClkMux
    port map (
            O => \N__46073\,
            I => \N__45627\
        );

    \I__10915\ : ClkMux
    port map (
            O => \N__46072\,
            I => \N__45627\
        );

    \I__10914\ : ClkMux
    port map (
            O => \N__46071\,
            I => \N__45627\
        );

    \I__10913\ : ClkMux
    port map (
            O => \N__46070\,
            I => \N__45627\
        );

    \I__10912\ : ClkMux
    port map (
            O => \N__46069\,
            I => \N__45627\
        );

    \I__10911\ : ClkMux
    port map (
            O => \N__46068\,
            I => \N__45627\
        );

    \I__10910\ : ClkMux
    port map (
            O => \N__46067\,
            I => \N__45627\
        );

    \I__10909\ : ClkMux
    port map (
            O => \N__46066\,
            I => \N__45627\
        );

    \I__10908\ : ClkMux
    port map (
            O => \N__46065\,
            I => \N__45627\
        );

    \I__10907\ : ClkMux
    port map (
            O => \N__46064\,
            I => \N__45627\
        );

    \I__10906\ : ClkMux
    port map (
            O => \N__46063\,
            I => \N__45627\
        );

    \I__10905\ : ClkMux
    port map (
            O => \N__46062\,
            I => \N__45627\
        );

    \I__10904\ : ClkMux
    port map (
            O => \N__46061\,
            I => \N__45627\
        );

    \I__10903\ : ClkMux
    port map (
            O => \N__46060\,
            I => \N__45627\
        );

    \I__10902\ : ClkMux
    port map (
            O => \N__46059\,
            I => \N__45627\
        );

    \I__10901\ : ClkMux
    port map (
            O => \N__46058\,
            I => \N__45627\
        );

    \I__10900\ : ClkMux
    port map (
            O => \N__46057\,
            I => \N__45627\
        );

    \I__10899\ : ClkMux
    port map (
            O => \N__46056\,
            I => \N__45627\
        );

    \I__10898\ : ClkMux
    port map (
            O => \N__46055\,
            I => \N__45627\
        );

    \I__10897\ : ClkMux
    port map (
            O => \N__46054\,
            I => \N__45627\
        );

    \I__10896\ : ClkMux
    port map (
            O => \N__46053\,
            I => \N__45627\
        );

    \I__10895\ : ClkMux
    port map (
            O => \N__46052\,
            I => \N__45627\
        );

    \I__10894\ : ClkMux
    port map (
            O => \N__46051\,
            I => \N__45627\
        );

    \I__10893\ : ClkMux
    port map (
            O => \N__46050\,
            I => \N__45627\
        );

    \I__10892\ : ClkMux
    port map (
            O => \N__46049\,
            I => \N__45627\
        );

    \I__10891\ : ClkMux
    port map (
            O => \N__46048\,
            I => \N__45627\
        );

    \I__10890\ : ClkMux
    port map (
            O => \N__46047\,
            I => \N__45627\
        );

    \I__10889\ : ClkMux
    port map (
            O => \N__46046\,
            I => \N__45627\
        );

    \I__10888\ : ClkMux
    port map (
            O => \N__46045\,
            I => \N__45627\
        );

    \I__10887\ : ClkMux
    port map (
            O => \N__46044\,
            I => \N__45627\
        );

    \I__10886\ : ClkMux
    port map (
            O => \N__46043\,
            I => \N__45627\
        );

    \I__10885\ : ClkMux
    port map (
            O => \N__46042\,
            I => \N__45627\
        );

    \I__10884\ : ClkMux
    port map (
            O => \N__46041\,
            I => \N__45627\
        );

    \I__10883\ : ClkMux
    port map (
            O => \N__46040\,
            I => \N__45627\
        );

    \I__10882\ : ClkMux
    port map (
            O => \N__46039\,
            I => \N__45627\
        );

    \I__10881\ : ClkMux
    port map (
            O => \N__46038\,
            I => \N__45627\
        );

    \I__10880\ : ClkMux
    port map (
            O => \N__46037\,
            I => \N__45627\
        );

    \I__10879\ : ClkMux
    port map (
            O => \N__46036\,
            I => \N__45627\
        );

    \I__10878\ : ClkMux
    port map (
            O => \N__46035\,
            I => \N__45627\
        );

    \I__10877\ : ClkMux
    port map (
            O => \N__46034\,
            I => \N__45627\
        );

    \I__10876\ : ClkMux
    port map (
            O => \N__46033\,
            I => \N__45627\
        );

    \I__10875\ : ClkMux
    port map (
            O => \N__46032\,
            I => \N__45627\
        );

    \I__10874\ : ClkMux
    port map (
            O => \N__46031\,
            I => \N__45627\
        );

    \I__10873\ : ClkMux
    port map (
            O => \N__46030\,
            I => \N__45627\
        );

    \I__10872\ : ClkMux
    port map (
            O => \N__46029\,
            I => \N__45627\
        );

    \I__10871\ : ClkMux
    port map (
            O => \N__46028\,
            I => \N__45627\
        );

    \I__10870\ : ClkMux
    port map (
            O => \N__46027\,
            I => \N__45627\
        );

    \I__10869\ : ClkMux
    port map (
            O => \N__46026\,
            I => \N__45627\
        );

    \I__10868\ : ClkMux
    port map (
            O => \N__46025\,
            I => \N__45627\
        );

    \I__10867\ : ClkMux
    port map (
            O => \N__46024\,
            I => \N__45627\
        );

    \I__10866\ : ClkMux
    port map (
            O => \N__46023\,
            I => \N__45627\
        );

    \I__10865\ : ClkMux
    port map (
            O => \N__46022\,
            I => \N__45627\
        );

    \I__10864\ : ClkMux
    port map (
            O => \N__46021\,
            I => \N__45627\
        );

    \I__10863\ : ClkMux
    port map (
            O => \N__46020\,
            I => \N__45627\
        );

    \I__10862\ : ClkMux
    port map (
            O => \N__46019\,
            I => \N__45627\
        );

    \I__10861\ : ClkMux
    port map (
            O => \N__46018\,
            I => \N__45627\
        );

    \I__10860\ : ClkMux
    port map (
            O => \N__46017\,
            I => \N__45627\
        );

    \I__10859\ : ClkMux
    port map (
            O => \N__46016\,
            I => \N__45627\
        );

    \I__10858\ : ClkMux
    port map (
            O => \N__46015\,
            I => \N__45627\
        );

    \I__10857\ : ClkMux
    port map (
            O => \N__46014\,
            I => \N__45627\
        );

    \I__10856\ : ClkMux
    port map (
            O => \N__46013\,
            I => \N__45627\
        );

    \I__10855\ : ClkMux
    port map (
            O => \N__46012\,
            I => \N__45627\
        );

    \I__10854\ : ClkMux
    port map (
            O => \N__46011\,
            I => \N__45627\
        );

    \I__10853\ : ClkMux
    port map (
            O => \N__46010\,
            I => \N__45627\
        );

    \I__10852\ : ClkMux
    port map (
            O => \N__46009\,
            I => \N__45627\
        );

    \I__10851\ : ClkMux
    port map (
            O => \N__46008\,
            I => \N__45627\
        );

    \I__10850\ : ClkMux
    port map (
            O => \N__46007\,
            I => \N__45627\
        );

    \I__10849\ : ClkMux
    port map (
            O => \N__46006\,
            I => \N__45627\
        );

    \I__10848\ : ClkMux
    port map (
            O => \N__46005\,
            I => \N__45627\
        );

    \I__10847\ : ClkMux
    port map (
            O => \N__46004\,
            I => \N__45627\
        );

    \I__10846\ : ClkMux
    port map (
            O => \N__46003\,
            I => \N__45627\
        );

    \I__10845\ : ClkMux
    port map (
            O => \N__46002\,
            I => \N__45627\
        );

    \I__10844\ : ClkMux
    port map (
            O => \N__46001\,
            I => \N__45627\
        );

    \I__10843\ : ClkMux
    port map (
            O => \N__46000\,
            I => \N__45627\
        );

    \I__10842\ : ClkMux
    port map (
            O => \N__45999\,
            I => \N__45627\
        );

    \I__10841\ : ClkMux
    port map (
            O => \N__45998\,
            I => \N__45627\
        );

    \I__10840\ : ClkMux
    port map (
            O => \N__45997\,
            I => \N__45627\
        );

    \I__10839\ : ClkMux
    port map (
            O => \N__45996\,
            I => \N__45627\
        );

    \I__10838\ : ClkMux
    port map (
            O => \N__45995\,
            I => \N__45627\
        );

    \I__10837\ : ClkMux
    port map (
            O => \N__45994\,
            I => \N__45627\
        );

    \I__10836\ : ClkMux
    port map (
            O => \N__45993\,
            I => \N__45627\
        );

    \I__10835\ : ClkMux
    port map (
            O => \N__45992\,
            I => \N__45627\
        );

    \I__10834\ : ClkMux
    port map (
            O => \N__45991\,
            I => \N__45627\
        );

    \I__10833\ : ClkMux
    port map (
            O => \N__45990\,
            I => \N__45627\
        );

    \I__10832\ : ClkMux
    port map (
            O => \N__45989\,
            I => \N__45627\
        );

    \I__10831\ : ClkMux
    port map (
            O => \N__45988\,
            I => \N__45627\
        );

    \I__10830\ : ClkMux
    port map (
            O => \N__45987\,
            I => \N__45627\
        );

    \I__10829\ : ClkMux
    port map (
            O => \N__45986\,
            I => \N__45627\
        );

    \I__10828\ : ClkMux
    port map (
            O => \N__45985\,
            I => \N__45627\
        );

    \I__10827\ : ClkMux
    port map (
            O => \N__45984\,
            I => \N__45627\
        );

    \I__10826\ : ClkMux
    port map (
            O => \N__45983\,
            I => \N__45627\
        );

    \I__10825\ : ClkMux
    port map (
            O => \N__45982\,
            I => \N__45627\
        );

    \I__10824\ : ClkMux
    port map (
            O => \N__45981\,
            I => \N__45627\
        );

    \I__10823\ : ClkMux
    port map (
            O => \N__45980\,
            I => \N__45627\
        );

    \I__10822\ : ClkMux
    port map (
            O => \N__45979\,
            I => \N__45627\
        );

    \I__10821\ : ClkMux
    port map (
            O => \N__45978\,
            I => \N__45627\
        );

    \I__10820\ : ClkMux
    port map (
            O => \N__45977\,
            I => \N__45627\
        );

    \I__10819\ : ClkMux
    port map (
            O => \N__45976\,
            I => \N__45627\
        );

    \I__10818\ : ClkMux
    port map (
            O => \N__45975\,
            I => \N__45627\
        );

    \I__10817\ : ClkMux
    port map (
            O => \N__45974\,
            I => \N__45627\
        );

    \I__10816\ : ClkMux
    port map (
            O => \N__45973\,
            I => \N__45627\
        );

    \I__10815\ : ClkMux
    port map (
            O => \N__45972\,
            I => \N__45627\
        );

    \I__10814\ : ClkMux
    port map (
            O => \N__45971\,
            I => \N__45627\
        );

    \I__10813\ : ClkMux
    port map (
            O => \N__45970\,
            I => \N__45627\
        );

    \I__10812\ : ClkMux
    port map (
            O => \N__45969\,
            I => \N__45627\
        );

    \I__10811\ : ClkMux
    port map (
            O => \N__45968\,
            I => \N__45627\
        );

    \I__10810\ : ClkMux
    port map (
            O => \N__45967\,
            I => \N__45627\
        );

    \I__10809\ : ClkMux
    port map (
            O => \N__45966\,
            I => \N__45627\
        );

    \I__10808\ : ClkMux
    port map (
            O => \N__45965\,
            I => \N__45627\
        );

    \I__10807\ : ClkMux
    port map (
            O => \N__45964\,
            I => \N__45627\
        );

    \I__10806\ : ClkMux
    port map (
            O => \N__45963\,
            I => \N__45627\
        );

    \I__10805\ : ClkMux
    port map (
            O => \N__45962\,
            I => \N__45627\
        );

    \I__10804\ : ClkMux
    port map (
            O => \N__45961\,
            I => \N__45627\
        );

    \I__10803\ : ClkMux
    port map (
            O => \N__45960\,
            I => \N__45627\
        );

    \I__10802\ : ClkMux
    port map (
            O => \N__45959\,
            I => \N__45627\
        );

    \I__10801\ : ClkMux
    port map (
            O => \N__45958\,
            I => \N__45627\
        );

    \I__10800\ : ClkMux
    port map (
            O => \N__45957\,
            I => \N__45627\
        );

    \I__10799\ : ClkMux
    port map (
            O => \N__45956\,
            I => \N__45627\
        );

    \I__10798\ : ClkMux
    port map (
            O => \N__45955\,
            I => \N__45627\
        );

    \I__10797\ : ClkMux
    port map (
            O => \N__45954\,
            I => \N__45627\
        );

    \I__10796\ : ClkMux
    port map (
            O => \N__45953\,
            I => \N__45627\
        );

    \I__10795\ : ClkMux
    port map (
            O => \N__45952\,
            I => \N__45627\
        );

    \I__10794\ : ClkMux
    port map (
            O => \N__45951\,
            I => \N__45627\
        );

    \I__10793\ : ClkMux
    port map (
            O => \N__45950\,
            I => \N__45627\
        );

    \I__10792\ : ClkMux
    port map (
            O => \N__45949\,
            I => \N__45627\
        );

    \I__10791\ : ClkMux
    port map (
            O => \N__45948\,
            I => \N__45627\
        );

    \I__10790\ : ClkMux
    port map (
            O => \N__45947\,
            I => \N__45627\
        );

    \I__10789\ : ClkMux
    port map (
            O => \N__45946\,
            I => \N__45627\
        );

    \I__10788\ : ClkMux
    port map (
            O => \N__45945\,
            I => \N__45627\
        );

    \I__10787\ : ClkMux
    port map (
            O => \N__45944\,
            I => \N__45627\
        );

    \I__10786\ : ClkMux
    port map (
            O => \N__45943\,
            I => \N__45627\
        );

    \I__10785\ : ClkMux
    port map (
            O => \N__45942\,
            I => \N__45627\
        );

    \I__10784\ : ClkMux
    port map (
            O => \N__45941\,
            I => \N__45627\
        );

    \I__10783\ : ClkMux
    port map (
            O => \N__45940\,
            I => \N__45627\
        );

    \I__10782\ : ClkMux
    port map (
            O => \N__45939\,
            I => \N__45627\
        );

    \I__10781\ : ClkMux
    port map (
            O => \N__45938\,
            I => \N__45627\
        );

    \I__10780\ : ClkMux
    port map (
            O => \N__45937\,
            I => \N__45627\
        );

    \I__10779\ : ClkMux
    port map (
            O => \N__45936\,
            I => \N__45627\
        );

    \I__10778\ : ClkMux
    port map (
            O => \N__45935\,
            I => \N__45627\
        );

    \I__10777\ : ClkMux
    port map (
            O => \N__45934\,
            I => \N__45627\
        );

    \I__10776\ : ClkMux
    port map (
            O => \N__45933\,
            I => \N__45627\
        );

    \I__10775\ : ClkMux
    port map (
            O => \N__45932\,
            I => \N__45627\
        );

    \I__10774\ : ClkMux
    port map (
            O => \N__45931\,
            I => \N__45627\
        );

    \I__10773\ : ClkMux
    port map (
            O => \N__45930\,
            I => \N__45627\
        );

    \I__10772\ : ClkMux
    port map (
            O => \N__45929\,
            I => \N__45627\
        );

    \I__10771\ : ClkMux
    port map (
            O => \N__45928\,
            I => \N__45627\
        );

    \I__10770\ : GlobalMux
    port map (
            O => \N__45627\,
            I => clk_100mhz_0
        );

    \I__10769\ : CascadeMux
    port map (
            O => \N__45624\,
            I => \N__45615\
        );

    \I__10768\ : CascadeMux
    port map (
            O => \N__45623\,
            I => \N__45612\
        );

    \I__10767\ : InMux
    port map (
            O => \N__45622\,
            I => \N__45609\
        );

    \I__10766\ : InMux
    port map (
            O => \N__45621\,
            I => \N__45606\
        );

    \I__10765\ : InMux
    port map (
            O => \N__45620\,
            I => \N__45603\
        );

    \I__10764\ : InMux
    port map (
            O => \N__45619\,
            I => \N__45600\
        );

    \I__10763\ : InMux
    port map (
            O => \N__45618\,
            I => \N__45597\
        );

    \I__10762\ : InMux
    port map (
            O => \N__45615\,
            I => \N__45594\
        );

    \I__10761\ : InMux
    port map (
            O => \N__45612\,
            I => \N__45591\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__45609\,
            I => \N__45588\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__45606\,
            I => \N__45585\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__45603\,
            I => \N__45582\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__45600\,
            I => \N__45536\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__45597\,
            I => \N__45470\
        );

    \I__10755\ : LocalMux
    port map (
            O => \N__45594\,
            I => \N__45462\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__45591\,
            I => \N__45449\
        );

    \I__10753\ : Glb2LocalMux
    port map (
            O => \N__45588\,
            I => \N__45165\
        );

    \I__10752\ : Glb2LocalMux
    port map (
            O => \N__45585\,
            I => \N__45165\
        );

    \I__10751\ : Glb2LocalMux
    port map (
            O => \N__45582\,
            I => \N__45165\
        );

    \I__10750\ : SRMux
    port map (
            O => \N__45581\,
            I => \N__45165\
        );

    \I__10749\ : SRMux
    port map (
            O => \N__45580\,
            I => \N__45165\
        );

    \I__10748\ : SRMux
    port map (
            O => \N__45579\,
            I => \N__45165\
        );

    \I__10747\ : SRMux
    port map (
            O => \N__45578\,
            I => \N__45165\
        );

    \I__10746\ : SRMux
    port map (
            O => \N__45577\,
            I => \N__45165\
        );

    \I__10745\ : SRMux
    port map (
            O => \N__45576\,
            I => \N__45165\
        );

    \I__10744\ : SRMux
    port map (
            O => \N__45575\,
            I => \N__45165\
        );

    \I__10743\ : SRMux
    port map (
            O => \N__45574\,
            I => \N__45165\
        );

    \I__10742\ : SRMux
    port map (
            O => \N__45573\,
            I => \N__45165\
        );

    \I__10741\ : SRMux
    port map (
            O => \N__45572\,
            I => \N__45165\
        );

    \I__10740\ : SRMux
    port map (
            O => \N__45571\,
            I => \N__45165\
        );

    \I__10739\ : SRMux
    port map (
            O => \N__45570\,
            I => \N__45165\
        );

    \I__10738\ : SRMux
    port map (
            O => \N__45569\,
            I => \N__45165\
        );

    \I__10737\ : SRMux
    port map (
            O => \N__45568\,
            I => \N__45165\
        );

    \I__10736\ : SRMux
    port map (
            O => \N__45567\,
            I => \N__45165\
        );

    \I__10735\ : SRMux
    port map (
            O => \N__45566\,
            I => \N__45165\
        );

    \I__10734\ : SRMux
    port map (
            O => \N__45565\,
            I => \N__45165\
        );

    \I__10733\ : SRMux
    port map (
            O => \N__45564\,
            I => \N__45165\
        );

    \I__10732\ : SRMux
    port map (
            O => \N__45563\,
            I => \N__45165\
        );

    \I__10731\ : SRMux
    port map (
            O => \N__45562\,
            I => \N__45165\
        );

    \I__10730\ : SRMux
    port map (
            O => \N__45561\,
            I => \N__45165\
        );

    \I__10729\ : SRMux
    port map (
            O => \N__45560\,
            I => \N__45165\
        );

    \I__10728\ : SRMux
    port map (
            O => \N__45559\,
            I => \N__45165\
        );

    \I__10727\ : SRMux
    port map (
            O => \N__45558\,
            I => \N__45165\
        );

    \I__10726\ : SRMux
    port map (
            O => \N__45557\,
            I => \N__45165\
        );

    \I__10725\ : SRMux
    port map (
            O => \N__45556\,
            I => \N__45165\
        );

    \I__10724\ : SRMux
    port map (
            O => \N__45555\,
            I => \N__45165\
        );

    \I__10723\ : SRMux
    port map (
            O => \N__45554\,
            I => \N__45165\
        );

    \I__10722\ : SRMux
    port map (
            O => \N__45553\,
            I => \N__45165\
        );

    \I__10721\ : SRMux
    port map (
            O => \N__45552\,
            I => \N__45165\
        );

    \I__10720\ : SRMux
    port map (
            O => \N__45551\,
            I => \N__45165\
        );

    \I__10719\ : SRMux
    port map (
            O => \N__45550\,
            I => \N__45165\
        );

    \I__10718\ : SRMux
    port map (
            O => \N__45549\,
            I => \N__45165\
        );

    \I__10717\ : SRMux
    port map (
            O => \N__45548\,
            I => \N__45165\
        );

    \I__10716\ : SRMux
    port map (
            O => \N__45547\,
            I => \N__45165\
        );

    \I__10715\ : SRMux
    port map (
            O => \N__45546\,
            I => \N__45165\
        );

    \I__10714\ : SRMux
    port map (
            O => \N__45545\,
            I => \N__45165\
        );

    \I__10713\ : SRMux
    port map (
            O => \N__45544\,
            I => \N__45165\
        );

    \I__10712\ : SRMux
    port map (
            O => \N__45543\,
            I => \N__45165\
        );

    \I__10711\ : SRMux
    port map (
            O => \N__45542\,
            I => \N__45165\
        );

    \I__10710\ : SRMux
    port map (
            O => \N__45541\,
            I => \N__45165\
        );

    \I__10709\ : SRMux
    port map (
            O => \N__45540\,
            I => \N__45165\
        );

    \I__10708\ : SRMux
    port map (
            O => \N__45539\,
            I => \N__45165\
        );

    \I__10707\ : Glb2LocalMux
    port map (
            O => \N__45536\,
            I => \N__45165\
        );

    \I__10706\ : SRMux
    port map (
            O => \N__45535\,
            I => \N__45165\
        );

    \I__10705\ : SRMux
    port map (
            O => \N__45534\,
            I => \N__45165\
        );

    \I__10704\ : SRMux
    port map (
            O => \N__45533\,
            I => \N__45165\
        );

    \I__10703\ : SRMux
    port map (
            O => \N__45532\,
            I => \N__45165\
        );

    \I__10702\ : SRMux
    port map (
            O => \N__45531\,
            I => \N__45165\
        );

    \I__10701\ : SRMux
    port map (
            O => \N__45530\,
            I => \N__45165\
        );

    \I__10700\ : SRMux
    port map (
            O => \N__45529\,
            I => \N__45165\
        );

    \I__10699\ : SRMux
    port map (
            O => \N__45528\,
            I => \N__45165\
        );

    \I__10698\ : SRMux
    port map (
            O => \N__45527\,
            I => \N__45165\
        );

    \I__10697\ : SRMux
    port map (
            O => \N__45526\,
            I => \N__45165\
        );

    \I__10696\ : SRMux
    port map (
            O => \N__45525\,
            I => \N__45165\
        );

    \I__10695\ : SRMux
    port map (
            O => \N__45524\,
            I => \N__45165\
        );

    \I__10694\ : SRMux
    port map (
            O => \N__45523\,
            I => \N__45165\
        );

    \I__10693\ : SRMux
    port map (
            O => \N__45522\,
            I => \N__45165\
        );

    \I__10692\ : SRMux
    port map (
            O => \N__45521\,
            I => \N__45165\
        );

    \I__10691\ : SRMux
    port map (
            O => \N__45520\,
            I => \N__45165\
        );

    \I__10690\ : SRMux
    port map (
            O => \N__45519\,
            I => \N__45165\
        );

    \I__10689\ : SRMux
    port map (
            O => \N__45518\,
            I => \N__45165\
        );

    \I__10688\ : SRMux
    port map (
            O => \N__45517\,
            I => \N__45165\
        );

    \I__10687\ : SRMux
    port map (
            O => \N__45516\,
            I => \N__45165\
        );

    \I__10686\ : SRMux
    port map (
            O => \N__45515\,
            I => \N__45165\
        );

    \I__10685\ : SRMux
    port map (
            O => \N__45514\,
            I => \N__45165\
        );

    \I__10684\ : SRMux
    port map (
            O => \N__45513\,
            I => \N__45165\
        );

    \I__10683\ : SRMux
    port map (
            O => \N__45512\,
            I => \N__45165\
        );

    \I__10682\ : SRMux
    port map (
            O => \N__45511\,
            I => \N__45165\
        );

    \I__10681\ : SRMux
    port map (
            O => \N__45510\,
            I => \N__45165\
        );

    \I__10680\ : SRMux
    port map (
            O => \N__45509\,
            I => \N__45165\
        );

    \I__10679\ : SRMux
    port map (
            O => \N__45508\,
            I => \N__45165\
        );

    \I__10678\ : SRMux
    port map (
            O => \N__45507\,
            I => \N__45165\
        );

    \I__10677\ : SRMux
    port map (
            O => \N__45506\,
            I => \N__45165\
        );

    \I__10676\ : SRMux
    port map (
            O => \N__45505\,
            I => \N__45165\
        );

    \I__10675\ : SRMux
    port map (
            O => \N__45504\,
            I => \N__45165\
        );

    \I__10674\ : SRMux
    port map (
            O => \N__45503\,
            I => \N__45165\
        );

    \I__10673\ : SRMux
    port map (
            O => \N__45502\,
            I => \N__45165\
        );

    \I__10672\ : SRMux
    port map (
            O => \N__45501\,
            I => \N__45165\
        );

    \I__10671\ : SRMux
    port map (
            O => \N__45500\,
            I => \N__45165\
        );

    \I__10670\ : SRMux
    port map (
            O => \N__45499\,
            I => \N__45165\
        );

    \I__10669\ : SRMux
    port map (
            O => \N__45498\,
            I => \N__45165\
        );

    \I__10668\ : SRMux
    port map (
            O => \N__45497\,
            I => \N__45165\
        );

    \I__10667\ : SRMux
    port map (
            O => \N__45496\,
            I => \N__45165\
        );

    \I__10666\ : SRMux
    port map (
            O => \N__45495\,
            I => \N__45165\
        );

    \I__10665\ : SRMux
    port map (
            O => \N__45494\,
            I => \N__45165\
        );

    \I__10664\ : SRMux
    port map (
            O => \N__45493\,
            I => \N__45165\
        );

    \I__10663\ : SRMux
    port map (
            O => \N__45492\,
            I => \N__45165\
        );

    \I__10662\ : SRMux
    port map (
            O => \N__45491\,
            I => \N__45165\
        );

    \I__10661\ : SRMux
    port map (
            O => \N__45490\,
            I => \N__45165\
        );

    \I__10660\ : SRMux
    port map (
            O => \N__45489\,
            I => \N__45165\
        );

    \I__10659\ : SRMux
    port map (
            O => \N__45488\,
            I => \N__45165\
        );

    \I__10658\ : SRMux
    port map (
            O => \N__45487\,
            I => \N__45165\
        );

    \I__10657\ : SRMux
    port map (
            O => \N__45486\,
            I => \N__45165\
        );

    \I__10656\ : SRMux
    port map (
            O => \N__45485\,
            I => \N__45165\
        );

    \I__10655\ : SRMux
    port map (
            O => \N__45484\,
            I => \N__45165\
        );

    \I__10654\ : SRMux
    port map (
            O => \N__45483\,
            I => \N__45165\
        );

    \I__10653\ : SRMux
    port map (
            O => \N__45482\,
            I => \N__45165\
        );

    \I__10652\ : SRMux
    port map (
            O => \N__45481\,
            I => \N__45165\
        );

    \I__10651\ : SRMux
    port map (
            O => \N__45480\,
            I => \N__45165\
        );

    \I__10650\ : SRMux
    port map (
            O => \N__45479\,
            I => \N__45165\
        );

    \I__10649\ : SRMux
    port map (
            O => \N__45478\,
            I => \N__45165\
        );

    \I__10648\ : SRMux
    port map (
            O => \N__45477\,
            I => \N__45165\
        );

    \I__10647\ : SRMux
    port map (
            O => \N__45476\,
            I => \N__45165\
        );

    \I__10646\ : SRMux
    port map (
            O => \N__45475\,
            I => \N__45165\
        );

    \I__10645\ : SRMux
    port map (
            O => \N__45474\,
            I => \N__45165\
        );

    \I__10644\ : SRMux
    port map (
            O => \N__45473\,
            I => \N__45165\
        );

    \I__10643\ : Glb2LocalMux
    port map (
            O => \N__45470\,
            I => \N__45165\
        );

    \I__10642\ : SRMux
    port map (
            O => \N__45469\,
            I => \N__45165\
        );

    \I__10641\ : SRMux
    port map (
            O => \N__45468\,
            I => \N__45165\
        );

    \I__10640\ : SRMux
    port map (
            O => \N__45467\,
            I => \N__45165\
        );

    \I__10639\ : SRMux
    port map (
            O => \N__45466\,
            I => \N__45165\
        );

    \I__10638\ : SRMux
    port map (
            O => \N__45465\,
            I => \N__45165\
        );

    \I__10637\ : Glb2LocalMux
    port map (
            O => \N__45462\,
            I => \N__45165\
        );

    \I__10636\ : SRMux
    port map (
            O => \N__45461\,
            I => \N__45165\
        );

    \I__10635\ : SRMux
    port map (
            O => \N__45460\,
            I => \N__45165\
        );

    \I__10634\ : SRMux
    port map (
            O => \N__45459\,
            I => \N__45165\
        );

    \I__10633\ : SRMux
    port map (
            O => \N__45458\,
            I => \N__45165\
        );

    \I__10632\ : SRMux
    port map (
            O => \N__45457\,
            I => \N__45165\
        );

    \I__10631\ : SRMux
    port map (
            O => \N__45456\,
            I => \N__45165\
        );

    \I__10630\ : SRMux
    port map (
            O => \N__45455\,
            I => \N__45165\
        );

    \I__10629\ : SRMux
    port map (
            O => \N__45454\,
            I => \N__45165\
        );

    \I__10628\ : SRMux
    port map (
            O => \N__45453\,
            I => \N__45165\
        );

    \I__10627\ : SRMux
    port map (
            O => \N__45452\,
            I => \N__45165\
        );

    \I__10626\ : Glb2LocalMux
    port map (
            O => \N__45449\,
            I => \N__45165\
        );

    \I__10625\ : SRMux
    port map (
            O => \N__45448\,
            I => \N__45165\
        );

    \I__10624\ : SRMux
    port map (
            O => \N__45447\,
            I => \N__45165\
        );

    \I__10623\ : SRMux
    port map (
            O => \N__45446\,
            I => \N__45165\
        );

    \I__10622\ : SRMux
    port map (
            O => \N__45445\,
            I => \N__45165\
        );

    \I__10621\ : SRMux
    port map (
            O => \N__45444\,
            I => \N__45165\
        );

    \I__10620\ : SRMux
    port map (
            O => \N__45443\,
            I => \N__45165\
        );

    \I__10619\ : SRMux
    port map (
            O => \N__45442\,
            I => \N__45165\
        );

    \I__10618\ : SRMux
    port map (
            O => \N__45441\,
            I => \N__45165\
        );

    \I__10617\ : SRMux
    port map (
            O => \N__45440\,
            I => \N__45165\
        );

    \I__10616\ : GlobalMux
    port map (
            O => \N__45165\,
            I => \N__45162\
        );

    \I__10615\ : gio2CtrlBuf
    port map (
            O => \N__45162\,
            I => red_c_g
        );

    \I__10614\ : CascadeMux
    port map (
            O => \N__45159\,
            I => \N__45156\
        );

    \I__10613\ : InMux
    port map (
            O => \N__45156\,
            I => \N__45153\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__45153\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__10611\ : InMux
    port map (
            O => \N__45150\,
            I => \N__45146\
        );

    \I__10610\ : InMux
    port map (
            O => \N__45149\,
            I => \N__45143\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__45146\,
            I => \N__45140\
        );

    \I__10608\ : LocalMux
    port map (
            O => \N__45143\,
            I => \N__45137\
        );

    \I__10607\ : Odrv4
    port map (
            O => \N__45140\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__10606\ : Odrv4
    port map (
            O => \N__45137\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__10605\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45129\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__45129\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__10603\ : InMux
    port map (
            O => \N__45126\,
            I => \N__45123\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__45123\,
            I => \N__45119\
        );

    \I__10601\ : InMux
    port map (
            O => \N__45122\,
            I => \N__45116\
        );

    \I__10600\ : Span4Mux_v
    port map (
            O => \N__45119\,
            I => \N__45111\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__45116\,
            I => \N__45111\
        );

    \I__10598\ : Odrv4
    port map (
            O => \N__45111\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__10597\ : CascadeMux
    port map (
            O => \N__45108\,
            I => \N__45105\
        );

    \I__10596\ : InMux
    port map (
            O => \N__45105\,
            I => \N__45102\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__45102\,
            I => \N__45099\
        );

    \I__10594\ : Odrv4
    port map (
            O => \N__45099\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__10593\ : InMux
    port map (
            O => \N__45096\,
            I => \N__45093\
        );

    \I__10592\ : LocalMux
    port map (
            O => \N__45093\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__10591\ : InMux
    port map (
            O => \N__45090\,
            I => \N__45087\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__45087\,
            I => \N__45084\
        );

    \I__10589\ : Span4Mux_h
    port map (
            O => \N__45084\,
            I => \N__45081\
        );

    \I__10588\ : Odrv4
    port map (
            O => \N__45081\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__10587\ : InMux
    port map (
            O => \N__45078\,
            I => \N__45074\
        );

    \I__10586\ : InMux
    port map (
            O => \N__45077\,
            I => \N__45071\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__45074\,
            I => \N__45068\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__45071\,
            I => \N__45065\
        );

    \I__10583\ : Span4Mux_v
    port map (
            O => \N__45068\,
            I => \N__45062\
        );

    \I__10582\ : Odrv4
    port map (
            O => \N__45065\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__10581\ : Odrv4
    port map (
            O => \N__45062\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__10580\ : CascadeMux
    port map (
            O => \N__45057\,
            I => \N__45054\
        );

    \I__10579\ : InMux
    port map (
            O => \N__45054\,
            I => \N__45051\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__45051\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__10577\ : CascadeMux
    port map (
            O => \N__45048\,
            I => \N__45045\
        );

    \I__10576\ : InMux
    port map (
            O => \N__45045\,
            I => \N__45042\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__45042\,
            I => \N__45039\
        );

    \I__10574\ : Odrv4
    port map (
            O => \N__45039\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__10573\ : InMux
    port map (
            O => \N__45036\,
            I => \N__45033\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__45033\,
            I => \N__45029\
        );

    \I__10571\ : InMux
    port map (
            O => \N__45032\,
            I => \N__45026\
        );

    \I__10570\ : Span4Mux_h
    port map (
            O => \N__45029\,
            I => \N__45023\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__45026\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__10568\ : Odrv4
    port map (
            O => \N__45023\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__10567\ : InMux
    port map (
            O => \N__45018\,
            I => \N__45015\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__45015\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__10565\ : InMux
    port map (
            O => \N__45012\,
            I => \N__45009\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__45009\,
            I => \N__45005\
        );

    \I__10563\ : InMux
    port map (
            O => \N__45008\,
            I => \N__45002\
        );

    \I__10562\ : Span4Mux_v
    port map (
            O => \N__45005\,
            I => \N__44999\
        );

    \I__10561\ : LocalMux
    port map (
            O => \N__45002\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10560\ : Odrv4
    port map (
            O => \N__44999\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10559\ : InMux
    port map (
            O => \N__44994\,
            I => \N__44991\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__44991\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\
        );

    \I__10557\ : InMux
    port map (
            O => \N__44988\,
            I => \N__44984\
        );

    \I__10556\ : InMux
    port map (
            O => \N__44987\,
            I => \N__44981\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__44984\,
            I => \N__44978\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__44981\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10553\ : Odrv4
    port map (
            O => \N__44978\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10552\ : InMux
    port map (
            O => \N__44973\,
            I => \N__44970\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__44970\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\
        );

    \I__10550\ : CascadeMux
    port map (
            O => \N__44967\,
            I => \N__44964\
        );

    \I__10549\ : InMux
    port map (
            O => \N__44964\,
            I => \N__44961\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__44961\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__10547\ : InMux
    port map (
            O => \N__44958\,
            I => \N__44954\
        );

    \I__10546\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44951\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__44954\,
            I => \N__44948\
        );

    \I__10544\ : LocalMux
    port map (
            O => \N__44951\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10543\ : Odrv4
    port map (
            O => \N__44948\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10542\ : InMux
    port map (
            O => \N__44943\,
            I => \N__44940\
        );

    \I__10541\ : LocalMux
    port map (
            O => \N__44940\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\
        );

    \I__10540\ : InMux
    port map (
            O => \N__44937\,
            I => \N__44933\
        );

    \I__10539\ : InMux
    port map (
            O => \N__44936\,
            I => \N__44930\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__44933\,
            I => \N__44927\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__44930\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10536\ : Odrv4
    port map (
            O => \N__44927\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10535\ : InMux
    port map (
            O => \N__44922\,
            I => \N__44919\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__44919\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\
        );

    \I__10533\ : CascadeMux
    port map (
            O => \N__44916\,
            I => \N__44913\
        );

    \I__10532\ : InMux
    port map (
            O => \N__44913\,
            I => \N__44910\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__44910\,
            I => \N__44907\
        );

    \I__10530\ : Odrv4
    port map (
            O => \N__44907\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__10529\ : InMux
    port map (
            O => \N__44904\,
            I => \N__44901\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__44901\,
            I => \N__44897\
        );

    \I__10527\ : InMux
    port map (
            O => \N__44900\,
            I => \N__44894\
        );

    \I__10526\ : Odrv4
    port map (
            O => \N__44897\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__10525\ : LocalMux
    port map (
            O => \N__44894\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__10524\ : InMux
    port map (
            O => \N__44889\,
            I => \N__44886\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__44886\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__10522\ : InMux
    port map (
            O => \N__44883\,
            I => \N__44880\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__44880\,
            I => \N__44876\
        );

    \I__10520\ : InMux
    port map (
            O => \N__44879\,
            I => \N__44873\
        );

    \I__10519\ : Odrv4
    port map (
            O => \N__44876\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__44873\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__10517\ : CascadeMux
    port map (
            O => \N__44868\,
            I => \N__44865\
        );

    \I__10516\ : InMux
    port map (
            O => \N__44865\,
            I => \N__44862\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__44862\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__10514\ : InMux
    port map (
            O => \N__44859\,
            I => \N__44856\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__44856\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__10512\ : InMux
    port map (
            O => \N__44853\,
            I => \N__44850\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__44850\,
            I => \N__44846\
        );

    \I__10510\ : InMux
    port map (
            O => \N__44849\,
            I => \N__44843\
        );

    \I__10509\ : Odrv4
    port map (
            O => \N__44846\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__44843\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__10507\ : CascadeMux
    port map (
            O => \N__44838\,
            I => \N__44835\
        );

    \I__10506\ : InMux
    port map (
            O => \N__44835\,
            I => \N__44832\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__44832\,
            I => \N__44829\
        );

    \I__10504\ : Odrv4
    port map (
            O => \N__44829\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__10503\ : InMux
    port map (
            O => \N__44826\,
            I => \N__44823\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__44823\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__10501\ : InMux
    port map (
            O => \N__44820\,
            I => \N__44817\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__44817\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__10499\ : InMux
    port map (
            O => \N__44814\,
            I => \N__44810\
        );

    \I__10498\ : InMux
    port map (
            O => \N__44813\,
            I => \N__44807\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__44810\,
            I => \N__44804\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__44807\,
            I => \N__44801\
        );

    \I__10495\ : Odrv12
    port map (
            O => \N__44804\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__10494\ : Odrv4
    port map (
            O => \N__44801\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__10493\ : CascadeMux
    port map (
            O => \N__44796\,
            I => \N__44793\
        );

    \I__10492\ : InMux
    port map (
            O => \N__44793\,
            I => \N__44790\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__44790\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__10490\ : CascadeMux
    port map (
            O => \N__44787\,
            I => \N__44784\
        );

    \I__10489\ : InMux
    port map (
            O => \N__44784\,
            I => \N__44781\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__44781\,
            I => \N__44778\
        );

    \I__10487\ : Odrv4
    port map (
            O => \N__44778\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__10486\ : InMux
    port map (
            O => \N__44775\,
            I => \N__44771\
        );

    \I__10485\ : InMux
    port map (
            O => \N__44774\,
            I => \N__44768\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__44771\,
            I => \N__44765\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__44768\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__10482\ : Odrv4
    port map (
            O => \N__44765\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__10481\ : InMux
    port map (
            O => \N__44760\,
            I => \N__44757\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__44757\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__10479\ : CascadeMux
    port map (
            O => \N__44754\,
            I => \N__44751\
        );

    \I__10478\ : InMux
    port map (
            O => \N__44751\,
            I => \N__44748\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__44748\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__10476\ : InMux
    port map (
            O => \N__44745\,
            I => \N__44741\
        );

    \I__10475\ : InMux
    port map (
            O => \N__44744\,
            I => \N__44738\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__44741\,
            I => \N__44735\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__44738\,
            I => \N__44730\
        );

    \I__10472\ : Span12Mux_v
    port map (
            O => \N__44735\,
            I => \N__44730\
        );

    \I__10471\ : Odrv12
    port map (
            O => \N__44730\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__10470\ : InMux
    port map (
            O => \N__44727\,
            I => \N__44724\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__44724\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__10468\ : CascadeMux
    port map (
            O => \N__44721\,
            I => \N__44718\
        );

    \I__10467\ : InMux
    port map (
            O => \N__44718\,
            I => \N__44715\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__44715\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__10465\ : InMux
    port map (
            O => \N__44712\,
            I => \N__44709\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__44709\,
            I => \N__44705\
        );

    \I__10463\ : InMux
    port map (
            O => \N__44708\,
            I => \N__44702\
        );

    \I__10462\ : Span4Mux_v
    port map (
            O => \N__44705\,
            I => \N__44699\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__44702\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__10460\ : Odrv4
    port map (
            O => \N__44699\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__10459\ : InMux
    port map (
            O => \N__44694\,
            I => \N__44691\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__44691\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__10457\ : CascadeMux
    port map (
            O => \N__44688\,
            I => \N__44685\
        );

    \I__10456\ : InMux
    port map (
            O => \N__44685\,
            I => \N__44682\
        );

    \I__10455\ : LocalMux
    port map (
            O => \N__44682\,
            I => \N__44679\
        );

    \I__10454\ : Odrv12
    port map (
            O => \N__44679\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14\
        );

    \I__10453\ : InMux
    port map (
            O => \N__44676\,
            I => \N__44673\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__44673\,
            I => \N__44670\
        );

    \I__10451\ : Odrv4
    port map (
            O => \N__44670\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8\
        );

    \I__10450\ : InMux
    port map (
            O => \N__44667\,
            I => \N__44657\
        );

    \I__10449\ : InMux
    port map (
            O => \N__44666\,
            I => \N__44657\
        );

    \I__10448\ : CascadeMux
    port map (
            O => \N__44665\,
            I => \N__44654\
        );

    \I__10447\ : CascadeMux
    port map (
            O => \N__44664\,
            I => \N__44650\
        );

    \I__10446\ : CascadeMux
    port map (
            O => \N__44663\,
            I => \N__44636\
        );

    \I__10445\ : CascadeMux
    port map (
            O => \N__44662\,
            I => \N__44633\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__44657\,
            I => \N__44628\
        );

    \I__10443\ : InMux
    port map (
            O => \N__44654\,
            I => \N__44623\
        );

    \I__10442\ : InMux
    port map (
            O => \N__44653\,
            I => \N__44623\
        );

    \I__10441\ : InMux
    port map (
            O => \N__44650\,
            I => \N__44606\
        );

    \I__10440\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44606\
        );

    \I__10439\ : InMux
    port map (
            O => \N__44648\,
            I => \N__44606\
        );

    \I__10438\ : InMux
    port map (
            O => \N__44647\,
            I => \N__44606\
        );

    \I__10437\ : InMux
    port map (
            O => \N__44646\,
            I => \N__44606\
        );

    \I__10436\ : InMux
    port map (
            O => \N__44645\,
            I => \N__44606\
        );

    \I__10435\ : InMux
    port map (
            O => \N__44644\,
            I => \N__44606\
        );

    \I__10434\ : InMux
    port map (
            O => \N__44643\,
            I => \N__44606\
        );

    \I__10433\ : CascadeMux
    port map (
            O => \N__44642\,
            I => \N__44603\
        );

    \I__10432\ : CascadeMux
    port map (
            O => \N__44641\,
            I => \N__44600\
        );

    \I__10431\ : CascadeMux
    port map (
            O => \N__44640\,
            I => \N__44597\
        );

    \I__10430\ : InMux
    port map (
            O => \N__44639\,
            I => \N__44586\
        );

    \I__10429\ : InMux
    port map (
            O => \N__44636\,
            I => \N__44586\
        );

    \I__10428\ : InMux
    port map (
            O => \N__44633\,
            I => \N__44586\
        );

    \I__10427\ : InMux
    port map (
            O => \N__44632\,
            I => \N__44586\
        );

    \I__10426\ : InMux
    port map (
            O => \N__44631\,
            I => \N__44586\
        );

    \I__10425\ : Span4Mux_h
    port map (
            O => \N__44628\,
            I => \N__44579\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__44623\,
            I => \N__44579\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__44606\,
            I => \N__44576\
        );

    \I__10422\ : InMux
    port map (
            O => \N__44603\,
            I => \N__44569\
        );

    \I__10421\ : InMux
    port map (
            O => \N__44600\,
            I => \N__44569\
        );

    \I__10420\ : InMux
    port map (
            O => \N__44597\,
            I => \N__44569\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__44586\,
            I => \N__44566\
        );

    \I__10418\ : InMux
    port map (
            O => \N__44585\,
            I => \N__44561\
        );

    \I__10417\ : InMux
    port map (
            O => \N__44584\,
            I => \N__44561\
        );

    \I__10416\ : Span4Mux_v
    port map (
            O => \N__44579\,
            I => \N__44554\
        );

    \I__10415\ : Span4Mux_v
    port map (
            O => \N__44576\,
            I => \N__44554\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__44569\,
            I => \N__44547\
        );

    \I__10413\ : Span4Mux_v
    port map (
            O => \N__44566\,
            I => \N__44547\
        );

    \I__10412\ : LocalMux
    port map (
            O => \N__44561\,
            I => \N__44547\
        );

    \I__10411\ : InMux
    port map (
            O => \N__44560\,
            I => \N__44544\
        );

    \I__10410\ : CascadeMux
    port map (
            O => \N__44559\,
            I => \N__44541\
        );

    \I__10409\ : Span4Mux_h
    port map (
            O => \N__44554\,
            I => \N__44538\
        );

    \I__10408\ : Span4Mux_v
    port map (
            O => \N__44547\,
            I => \N__44535\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__44544\,
            I => \N__44532\
        );

    \I__10406\ : InMux
    port map (
            O => \N__44541\,
            I => \N__44529\
        );

    \I__10405\ : Span4Mux_v
    port map (
            O => \N__44538\,
            I => \N__44526\
        );

    \I__10404\ : Span4Mux_v
    port map (
            O => \N__44535\,
            I => \N__44523\
        );

    \I__10403\ : Span12Mux_h
    port map (
            O => \N__44532\,
            I => \N__44520\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__44529\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__10401\ : Odrv4
    port map (
            O => \N__44526\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__10400\ : Odrv4
    port map (
            O => \N__44523\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__10399\ : Odrv12
    port map (
            O => \N__44520\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__10398\ : CascadeMux
    port map (
            O => \N__44511\,
            I => \N__44502\
        );

    \I__10397\ : CascadeMux
    port map (
            O => \N__44510\,
            I => \N__44499\
        );

    \I__10396\ : CascadeMux
    port map (
            O => \N__44509\,
            I => \N__44496\
        );

    \I__10395\ : CascadeMux
    port map (
            O => \N__44508\,
            I => \N__44493\
        );

    \I__10394\ : CascadeMux
    port map (
            O => \N__44507\,
            I => \N__44486\
        );

    \I__10393\ : CascadeMux
    port map (
            O => \N__44506\,
            I => \N__44483\
        );

    \I__10392\ : CascadeMux
    port map (
            O => \N__44505\,
            I => \N__44478\
        );

    \I__10391\ : InMux
    port map (
            O => \N__44502\,
            I => \N__44455\
        );

    \I__10390\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44455\
        );

    \I__10389\ : InMux
    port map (
            O => \N__44496\,
            I => \N__44455\
        );

    \I__10388\ : InMux
    port map (
            O => \N__44493\,
            I => \N__44455\
        );

    \I__10387\ : InMux
    port map (
            O => \N__44492\,
            I => \N__44455\
        );

    \I__10386\ : InMux
    port map (
            O => \N__44491\,
            I => \N__44455\
        );

    \I__10385\ : InMux
    port map (
            O => \N__44490\,
            I => \N__44455\
        );

    \I__10384\ : InMux
    port map (
            O => \N__44489\,
            I => \N__44455\
        );

    \I__10383\ : InMux
    port map (
            O => \N__44486\,
            I => \N__44446\
        );

    \I__10382\ : InMux
    port map (
            O => \N__44483\,
            I => \N__44446\
        );

    \I__10381\ : InMux
    port map (
            O => \N__44482\,
            I => \N__44446\
        );

    \I__10380\ : InMux
    port map (
            O => \N__44481\,
            I => \N__44446\
        );

    \I__10379\ : InMux
    port map (
            O => \N__44478\,
            I => \N__44441\
        );

    \I__10378\ : InMux
    port map (
            O => \N__44477\,
            I => \N__44434\
        );

    \I__10377\ : InMux
    port map (
            O => \N__44476\,
            I => \N__44434\
        );

    \I__10376\ : InMux
    port map (
            O => \N__44475\,
            I => \N__44434\
        );

    \I__10375\ : CascadeMux
    port map (
            O => \N__44474\,
            I => \N__44430\
        );

    \I__10374\ : InMux
    port map (
            O => \N__44473\,
            I => \N__44423\
        );

    \I__10373\ : InMux
    port map (
            O => \N__44472\,
            I => \N__44423\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__44455\,
            I => \N__44418\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__44446\,
            I => \N__44418\
        );

    \I__10370\ : InMux
    port map (
            O => \N__44445\,
            I => \N__44413\
        );

    \I__10369\ : InMux
    port map (
            O => \N__44444\,
            I => \N__44413\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__44441\,
            I => \N__44410\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__44434\,
            I => \N__44407\
        );

    \I__10366\ : InMux
    port map (
            O => \N__44433\,
            I => \N__44404\
        );

    \I__10365\ : InMux
    port map (
            O => \N__44430\,
            I => \N__44397\
        );

    \I__10364\ : InMux
    port map (
            O => \N__44429\,
            I => \N__44397\
        );

    \I__10363\ : InMux
    port map (
            O => \N__44428\,
            I => \N__44397\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__44423\,
            I => \N__44394\
        );

    \I__10361\ : Span4Mux_v
    port map (
            O => \N__44418\,
            I => \N__44391\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__44413\,
            I => \N__44380\
        );

    \I__10359\ : Span4Mux_v
    port map (
            O => \N__44410\,
            I => \N__44380\
        );

    \I__10358\ : Span4Mux_h
    port map (
            O => \N__44407\,
            I => \N__44380\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__44404\,
            I => \N__44380\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__44397\,
            I => \N__44380\
        );

    \I__10355\ : Odrv4
    port map (
            O => \N__44394\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__10354\ : Odrv4
    port map (
            O => \N__44391\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__10353\ : Odrv4
    port map (
            O => \N__44380\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__10352\ : CascadeMux
    port map (
            O => \N__44373\,
            I => \N__44370\
        );

    \I__10351\ : InMux
    port map (
            O => \N__44370\,
            I => \N__44367\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__44367\,
            I => \N__44364\
        );

    \I__10349\ : Span4Mux_v
    port map (
            O => \N__44364\,
            I => \N__44361\
        );

    \I__10348\ : Odrv4
    port map (
            O => \N__44361\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2\
        );

    \I__10347\ : CascadeMux
    port map (
            O => \N__44358\,
            I => \N__44354\
        );

    \I__10346\ : InMux
    port map (
            O => \N__44357\,
            I => \N__44334\
        );

    \I__10345\ : InMux
    port map (
            O => \N__44354\,
            I => \N__44331\
        );

    \I__10344\ : InMux
    port map (
            O => \N__44353\,
            I => \N__44314\
        );

    \I__10343\ : InMux
    port map (
            O => \N__44352\,
            I => \N__44314\
        );

    \I__10342\ : InMux
    port map (
            O => \N__44351\,
            I => \N__44314\
        );

    \I__10341\ : InMux
    port map (
            O => \N__44350\,
            I => \N__44314\
        );

    \I__10340\ : InMux
    port map (
            O => \N__44349\,
            I => \N__44314\
        );

    \I__10339\ : InMux
    port map (
            O => \N__44348\,
            I => \N__44314\
        );

    \I__10338\ : InMux
    port map (
            O => \N__44347\,
            I => \N__44314\
        );

    \I__10337\ : InMux
    port map (
            O => \N__44346\,
            I => \N__44314\
        );

    \I__10336\ : InMux
    port map (
            O => \N__44345\,
            I => \N__44303\
        );

    \I__10335\ : InMux
    port map (
            O => \N__44344\,
            I => \N__44303\
        );

    \I__10334\ : InMux
    port map (
            O => \N__44343\,
            I => \N__44303\
        );

    \I__10333\ : InMux
    port map (
            O => \N__44342\,
            I => \N__44303\
        );

    \I__10332\ : InMux
    port map (
            O => \N__44341\,
            I => \N__44303\
        );

    \I__10331\ : CascadeMux
    port map (
            O => \N__44340\,
            I => \N__44295\
        );

    \I__10330\ : InMux
    port map (
            O => \N__44339\,
            I => \N__44288\
        );

    \I__10329\ : InMux
    port map (
            O => \N__44338\,
            I => \N__44288\
        );

    \I__10328\ : InMux
    port map (
            O => \N__44337\,
            I => \N__44288\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__44334\,
            I => \N__44283\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__44331\,
            I => \N__44283\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__44314\,
            I => \N__44278\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__44303\,
            I => \N__44278\
        );

    \I__10323\ : InMux
    port map (
            O => \N__44302\,
            I => \N__44275\
        );

    \I__10322\ : InMux
    port map (
            O => \N__44301\,
            I => \N__44268\
        );

    \I__10321\ : InMux
    port map (
            O => \N__44300\,
            I => \N__44268\
        );

    \I__10320\ : InMux
    port map (
            O => \N__44299\,
            I => \N__44268\
        );

    \I__10319\ : InMux
    port map (
            O => \N__44298\,
            I => \N__44263\
        );

    \I__10318\ : InMux
    port map (
            O => \N__44295\,
            I => \N__44263\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__44288\,
            I => \N__44252\
        );

    \I__10316\ : Span4Mux_v
    port map (
            O => \N__44283\,
            I => \N__44252\
        );

    \I__10315\ : Span4Mux_v
    port map (
            O => \N__44278\,
            I => \N__44252\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__44275\,
            I => \N__44252\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__44268\,
            I => \N__44252\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__44263\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10311\ : Odrv4
    port map (
            O => \N__44252\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10310\ : CascadeMux
    port map (
            O => \N__44247\,
            I => \N__44244\
        );

    \I__10309\ : InMux
    port map (
            O => \N__44244\,
            I => \N__44241\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__44241\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_0\
        );

    \I__10307\ : CascadeMux
    port map (
            O => \N__44238\,
            I => \N__44235\
        );

    \I__10306\ : InMux
    port map (
            O => \N__44235\,
            I => \N__44232\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__44232\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__10304\ : CascadeMux
    port map (
            O => \N__44229\,
            I => \N__44225\
        );

    \I__10303\ : InMux
    port map (
            O => \N__44228\,
            I => \N__44222\
        );

    \I__10302\ : InMux
    port map (
            O => \N__44225\,
            I => \N__44218\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__44222\,
            I => \N__44215\
        );

    \I__10300\ : InMux
    port map (
            O => \N__44221\,
            I => \N__44212\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__44218\,
            I => \N__44207\
        );

    \I__10298\ : Span12Mux_v
    port map (
            O => \N__44215\,
            I => \N__44207\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__44212\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10296\ : Odrv12
    port map (
            O => \N__44207\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10295\ : InMux
    port map (
            O => \N__44202\,
            I => \N__44199\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__44199\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__10293\ : CascadeMux
    port map (
            O => \N__44196\,
            I => \N__44193\
        );

    \I__10292\ : InMux
    port map (
            O => \N__44193\,
            I => \N__44190\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__44190\,
            I => \N__44187\
        );

    \I__10290\ : Odrv4
    port map (
            O => \N__44187\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__10289\ : InMux
    port map (
            O => \N__44184\,
            I => \N__44181\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__44181\,
            I => \N__44177\
        );

    \I__10287\ : InMux
    port map (
            O => \N__44180\,
            I => \N__44174\
        );

    \I__10286\ : Odrv12
    port map (
            O => \N__44177\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__44174\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__10284\ : InMux
    port map (
            O => \N__44169\,
            I => \N__44166\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__44166\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__10282\ : CascadeMux
    port map (
            O => \N__44163\,
            I => \N__44160\
        );

    \I__10281\ : InMux
    port map (
            O => \N__44160\,
            I => \N__44157\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__44157\,
            I => \N__44153\
        );

    \I__10279\ : InMux
    port map (
            O => \N__44156\,
            I => \N__44150\
        );

    \I__10278\ : Odrv4
    port map (
            O => \N__44153\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__44150\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__10276\ : CascadeMux
    port map (
            O => \N__44145\,
            I => \N__44142\
        );

    \I__10275\ : InMux
    port map (
            O => \N__44142\,
            I => \N__44139\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__44139\,
            I => \N__44136\
        );

    \I__10273\ : Span4Mux_h
    port map (
            O => \N__44136\,
            I => \N__44133\
        );

    \I__10272\ : Odrv4
    port map (
            O => \N__44133\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__10271\ : InMux
    port map (
            O => \N__44130\,
            I => \N__44127\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__44127\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__10269\ : CascadeMux
    port map (
            O => \N__44124\,
            I => \N__44121\
        );

    \I__10268\ : InMux
    port map (
            O => \N__44121\,
            I => \N__44118\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__44118\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__10266\ : InMux
    port map (
            O => \N__44115\,
            I => \N__44112\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__44112\,
            I => \N__44108\
        );

    \I__10264\ : InMux
    port map (
            O => \N__44111\,
            I => \N__44105\
        );

    \I__10263\ : Odrv12
    port map (
            O => \N__44108\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__44105\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__10261\ : InMux
    port map (
            O => \N__44100\,
            I => \N__44097\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__44097\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__10259\ : InMux
    port map (
            O => \N__44094\,
            I => \N__44091\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__44091\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17\
        );

    \I__10257\ : InMux
    port map (
            O => \N__44088\,
            I => \bfn_18_15_0_\
        );

    \I__10256\ : InMux
    port map (
            O => \N__44085\,
            I => \N__44082\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__44082\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18\
        );

    \I__10254\ : InMux
    port map (
            O => \N__44079\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44076\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__10252\ : InMux
    port map (
            O => \N__44073\,
            I => \N__44070\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__44070\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19\
        );

    \I__10250\ : InMux
    port map (
            O => \N__44067\,
            I => \N__44064\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__44064\,
            I => \N__44061\
        );

    \I__10248\ : Odrv4
    port map (
            O => \N__44061\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3\
        );

    \I__10247\ : CascadeMux
    port map (
            O => \N__44058\,
            I => \N__44055\
        );

    \I__10246\ : InMux
    port map (
            O => \N__44055\,
            I => \N__44052\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__44052\,
            I => \N__44049\
        );

    \I__10244\ : Odrv4
    port map (
            O => \N__44049\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44046\,
            I => \N__44043\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__44043\,
            I => \N__44040\
        );

    \I__10241\ : Odrv4
    port map (
            O => \N__44040\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6\
        );

    \I__10240\ : InMux
    port map (
            O => \N__44037\,
            I => \N__44034\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__44034\,
            I => \N__44031\
        );

    \I__10238\ : Odrv4
    port map (
            O => \N__44031\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12\
        );

    \I__10237\ : InMux
    port map (
            O => \N__44028\,
            I => \N__44025\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__44025\,
            I => \N__44022\
        );

    \I__10235\ : Odrv4
    port map (
            O => \N__44022\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4\
        );

    \I__10234\ : InMux
    port map (
            O => \N__44019\,
            I => \N__44016\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__44016\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44013\,
            I => \bfn_18_14_0_\
        );

    \I__10231\ : InMux
    port map (
            O => \N__44010\,
            I => \N__44007\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__44007\,
            I => \N__44004\
        );

    \I__10229\ : Odrv12
    port map (
            O => \N__44004\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10\
        );

    \I__10228\ : InMux
    port map (
            O => \N__44001\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__10227\ : InMux
    port map (
            O => \N__43998\,
            I => \N__43995\
        );

    \I__10226\ : LocalMux
    port map (
            O => \N__43995\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11\
        );

    \I__10225\ : InMux
    port map (
            O => \N__43992\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__10224\ : InMux
    port map (
            O => \N__43989\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__10223\ : InMux
    port map (
            O => \N__43986\,
            I => \N__43983\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__43983\,
            I => \N__43980\
        );

    \I__10221\ : Odrv4
    port map (
            O => \N__43980\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13\
        );

    \I__10220\ : InMux
    port map (
            O => \N__43977\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__10219\ : InMux
    port map (
            O => \N__43974\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__10218\ : InMux
    port map (
            O => \N__43971\,
            I => \N__43968\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__43968\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15\
        );

    \I__10216\ : InMux
    port map (
            O => \N__43965\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__10215\ : InMux
    port map (
            O => \N__43962\,
            I => \N__43959\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__43959\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16\
        );

    \I__10213\ : InMux
    port map (
            O => \N__43956\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__10212\ : InMux
    port map (
            O => \N__43953\,
            I => \N__43949\
        );

    \I__10211\ : CascadeMux
    port map (
            O => \N__43952\,
            I => \N__43946\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__43949\,
            I => \N__43941\
        );

    \I__10209\ : InMux
    port map (
            O => \N__43946\,
            I => \N__43936\
        );

    \I__10208\ : InMux
    port map (
            O => \N__43945\,
            I => \N__43936\
        );

    \I__10207\ : InMux
    port map (
            O => \N__43944\,
            I => \N__43933\
        );

    \I__10206\ : Span4Mux_v
    port map (
            O => \N__43941\,
            I => \N__43928\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__43936\,
            I => \N__43928\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__43933\,
            I => \phase_controller_inst2.stoper_hc.time_passed11\
        );

    \I__10203\ : Odrv4
    port map (
            O => \N__43928\,
            I => \phase_controller_inst2.stoper_hc.time_passed11\
        );

    \I__10202\ : InMux
    port map (
            O => \N__43923\,
            I => \N__43920\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__43920\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__10200\ : InMux
    port map (
            O => \N__43917\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__10199\ : InMux
    port map (
            O => \N__43914\,
            I => \N__43911\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__43911\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0\
        );

    \I__10197\ : InMux
    port map (
            O => \N__43908\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__10196\ : InMux
    port map (
            O => \N__43905\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__10195\ : InMux
    port map (
            O => \N__43902\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__10194\ : InMux
    port map (
            O => \N__43899\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__10193\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43893\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__43893\,
            I => \N__43890\
        );

    \I__10191\ : Odrv4
    port map (
            O => \N__43890\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7\
        );

    \I__10190\ : InMux
    port map (
            O => \N__43887\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__10189\ : InMux
    port map (
            O => \N__43884\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__10188\ : InMux
    port map (
            O => \N__43881\,
            I => \N__43877\
        );

    \I__10187\ : InMux
    port map (
            O => \N__43880\,
            I => \N__43874\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__43877\,
            I => \N__43871\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__43874\,
            I => \N__43867\
        );

    \I__10184\ : Span4Mux_v
    port map (
            O => \N__43871\,
            I => \N__43864\
        );

    \I__10183\ : InMux
    port map (
            O => \N__43870\,
            I => \N__43861\
        );

    \I__10182\ : Odrv4
    port map (
            O => \N__43867\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10181\ : Odrv4
    port map (
            O => \N__43864\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__43861\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10179\ : InMux
    port map (
            O => \N__43854\,
            I => \N__43851\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__43851\,
            I => \N__43847\
        );

    \I__10177\ : CascadeMux
    port map (
            O => \N__43850\,
            I => \N__43844\
        );

    \I__10176\ : Span4Mux_v
    port map (
            O => \N__43847\,
            I => \N__43841\
        );

    \I__10175\ : InMux
    port map (
            O => \N__43844\,
            I => \N__43838\
        );

    \I__10174\ : Span4Mux_v
    port map (
            O => \N__43841\,
            I => \N__43833\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__43838\,
            I => \N__43833\
        );

    \I__10172\ : Odrv4
    port map (
            O => \N__43833\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__10171\ : CEMux
    port map (
            O => \N__43830\,
            I => \N__43812\
        );

    \I__10170\ : CEMux
    port map (
            O => \N__43829\,
            I => \N__43812\
        );

    \I__10169\ : CEMux
    port map (
            O => \N__43828\,
            I => \N__43812\
        );

    \I__10168\ : CEMux
    port map (
            O => \N__43827\,
            I => \N__43812\
        );

    \I__10167\ : CEMux
    port map (
            O => \N__43826\,
            I => \N__43812\
        );

    \I__10166\ : CEMux
    port map (
            O => \N__43825\,
            I => \N__43812\
        );

    \I__10165\ : GlobalMux
    port map (
            O => \N__43812\,
            I => \N__43809\
        );

    \I__10164\ : gio2CtrlBuf
    port map (
            O => \N__43809\,
            I => \delay_measurement_inst.delay_tr_timer.N_463_i_g\
        );

    \I__10163\ : CascadeMux
    port map (
            O => \N__43806\,
            I => \N__43802\
        );

    \I__10162\ : InMux
    port map (
            O => \N__43805\,
            I => \N__43798\
        );

    \I__10161\ : InMux
    port map (
            O => \N__43802\,
            I => \N__43793\
        );

    \I__10160\ : InMux
    port map (
            O => \N__43801\,
            I => \N__43793\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__43798\,
            I => \N__43790\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__43793\,
            I => \N__43787\
        );

    \I__10157\ : Span4Mux_h
    port map (
            O => \N__43790\,
            I => \N__43784\
        );

    \I__10156\ : Span4Mux_h
    port map (
            O => \N__43787\,
            I => \N__43781\
        );

    \I__10155\ : Odrv4
    port map (
            O => \N__43784\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__10154\ : Odrv4
    port map (
            O => \N__43781\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__10153\ : InMux
    port map (
            O => \N__43776\,
            I => \N__43772\
        );

    \I__10152\ : InMux
    port map (
            O => \N__43775\,
            I => \N__43769\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__43772\,
            I => \N__43766\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__43769\,
            I => \N__43763\
        );

    \I__10149\ : Span4Mux_v
    port map (
            O => \N__43766\,
            I => \N__43758\
        );

    \I__10148\ : Span4Mux_v
    port map (
            O => \N__43763\,
            I => \N__43755\
        );

    \I__10147\ : InMux
    port map (
            O => \N__43762\,
            I => \N__43750\
        );

    \I__10146\ : InMux
    port map (
            O => \N__43761\,
            I => \N__43750\
        );

    \I__10145\ : Span4Mux_h
    port map (
            O => \N__43758\,
            I => \N__43747\
        );

    \I__10144\ : Span4Mux_h
    port map (
            O => \N__43755\,
            I => \N__43742\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__43750\,
            I => \N__43742\
        );

    \I__10142\ : Sp12to4
    port map (
            O => \N__43747\,
            I => \N__43739\
        );

    \I__10141\ : Span4Mux_h
    port map (
            O => \N__43742\,
            I => \N__43736\
        );

    \I__10140\ : Odrv12
    port map (
            O => \N__43739\,
            I => measured_delay_tr_17
        );

    \I__10139\ : Odrv4
    port map (
            O => \N__43736\,
            I => measured_delay_tr_17
        );

    \I__10138\ : InMux
    port map (
            O => \N__43731\,
            I => \N__43723\
        );

    \I__10137\ : InMux
    port map (
            O => \N__43730\,
            I => \N__43723\
        );

    \I__10136\ : InMux
    port map (
            O => \N__43729\,
            I => \N__43716\
        );

    \I__10135\ : InMux
    port map (
            O => \N__43728\,
            I => \N__43716\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__43723\,
            I => \N__43713\
        );

    \I__10133\ : InMux
    port map (
            O => \N__43722\,
            I => \N__43708\
        );

    \I__10132\ : InMux
    port map (
            O => \N__43721\,
            I => \N__43708\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__43716\,
            I => \N__43702\
        );

    \I__10130\ : Span4Mux_h
    port map (
            O => \N__43713\,
            I => \N__43699\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__43708\,
            I => \N__43696\
        );

    \I__10128\ : InMux
    port map (
            O => \N__43707\,
            I => \N__43691\
        );

    \I__10127\ : InMux
    port map (
            O => \N__43706\,
            I => \N__43691\
        );

    \I__10126\ : InMux
    port map (
            O => \N__43705\,
            I => \N__43688\
        );

    \I__10125\ : Odrv4
    port map (
            O => \N__43702\,
            I => \delay_measurement_inst.N_498\
        );

    \I__10124\ : Odrv4
    port map (
            O => \N__43699\,
            I => \delay_measurement_inst.N_498\
        );

    \I__10123\ : Odrv4
    port map (
            O => \N__43696\,
            I => \delay_measurement_inst.N_498\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__43691\,
            I => \delay_measurement_inst.N_498\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__43688\,
            I => \delay_measurement_inst.N_498\
        );

    \I__10120\ : CascadeMux
    port map (
            O => \N__43677\,
            I => \N__43667\
        );

    \I__10119\ : CascadeMux
    port map (
            O => \N__43676\,
            I => \N__43662\
        );

    \I__10118\ : CascadeMux
    port map (
            O => \N__43675\,
            I => \N__43657\
        );

    \I__10117\ : CascadeMux
    port map (
            O => \N__43674\,
            I => \N__43654\
        );

    \I__10116\ : InMux
    port map (
            O => \N__43673\,
            I => \N__43649\
        );

    \I__10115\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43649\
        );

    \I__10114\ : InMux
    port map (
            O => \N__43671\,
            I => \N__43636\
        );

    \I__10113\ : InMux
    port map (
            O => \N__43670\,
            I => \N__43636\
        );

    \I__10112\ : InMux
    port map (
            O => \N__43667\,
            I => \N__43636\
        );

    \I__10111\ : InMux
    port map (
            O => \N__43666\,
            I => \N__43636\
        );

    \I__10110\ : InMux
    port map (
            O => \N__43665\,
            I => \N__43636\
        );

    \I__10109\ : InMux
    port map (
            O => \N__43662\,
            I => \N__43629\
        );

    \I__10108\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43629\
        );

    \I__10107\ : InMux
    port map (
            O => \N__43660\,
            I => \N__43629\
        );

    \I__10106\ : InMux
    port map (
            O => \N__43657\,
            I => \N__43626\
        );

    \I__10105\ : InMux
    port map (
            O => \N__43654\,
            I => \N__43623\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__43649\,
            I => \N__43620\
        );

    \I__10103\ : InMux
    port map (
            O => \N__43648\,
            I => \N__43615\
        );

    \I__10102\ : InMux
    port map (
            O => \N__43647\,
            I => \N__43615\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__43636\,
            I => \N__43610\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__43629\,
            I => \N__43610\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__43626\,
            I => \N__43607\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__43623\,
            I => \N__43604\
        );

    \I__10097\ : Span4Mux_v
    port map (
            O => \N__43620\,
            I => \N__43601\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__43615\,
            I => \N__43598\
        );

    \I__10095\ : Span4Mux_h
    port map (
            O => \N__43610\,
            I => \N__43595\
        );

    \I__10094\ : Span4Mux_v
    port map (
            O => \N__43607\,
            I => \N__43590\
        );

    \I__10093\ : Span4Mux_v
    port map (
            O => \N__43604\,
            I => \N__43590\
        );

    \I__10092\ : Odrv4
    port map (
            O => \N__43601\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__10091\ : Odrv12
    port map (
            O => \N__43598\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__10090\ : Odrv4
    port map (
            O => \N__43595\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__10089\ : Odrv4
    port map (
            O => \N__43590\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__10088\ : InMux
    port map (
            O => \N__43581\,
            I => \N__43578\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__43578\,
            I => \N__43573\
        );

    \I__10086\ : InMux
    port map (
            O => \N__43577\,
            I => \N__43568\
        );

    \I__10085\ : InMux
    port map (
            O => \N__43576\,
            I => \N__43568\
        );

    \I__10084\ : Span4Mux_h
    port map (
            O => \N__43573\,
            I => \N__43565\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__43568\,
            I => \N__43562\
        );

    \I__10082\ : Odrv4
    port map (
            O => \N__43565\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__10081\ : Odrv4
    port map (
            O => \N__43562\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__10080\ : InMux
    port map (
            O => \N__43557\,
            I => \N__43553\
        );

    \I__10079\ : InMux
    port map (
            O => \N__43556\,
            I => \N__43550\
        );

    \I__10078\ : LocalMux
    port map (
            O => \N__43553\,
            I => \N__43547\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__43550\,
            I => \N__43544\
        );

    \I__10076\ : Span4Mux_v
    port map (
            O => \N__43547\,
            I => \N__43539\
        );

    \I__10075\ : Span4Mux_v
    port map (
            O => \N__43544\,
            I => \N__43536\
        );

    \I__10074\ : InMux
    port map (
            O => \N__43543\,
            I => \N__43531\
        );

    \I__10073\ : InMux
    port map (
            O => \N__43542\,
            I => \N__43531\
        );

    \I__10072\ : Sp12to4
    port map (
            O => \N__43539\,
            I => \N__43524\
        );

    \I__10071\ : Sp12to4
    port map (
            O => \N__43536\,
            I => \N__43524\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__43531\,
            I => \N__43524\
        );

    \I__10069\ : Odrv12
    port map (
            O => \N__43524\,
            I => measured_delay_tr_18
        );

    \I__10068\ : CEMux
    port map (
            O => \N__43521\,
            I => \N__43516\
        );

    \I__10067\ : CEMux
    port map (
            O => \N__43520\,
            I => \N__43512\
        );

    \I__10066\ : CEMux
    port map (
            O => \N__43519\,
            I => \N__43508\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__43516\,
            I => \N__43505\
        );

    \I__10064\ : CEMux
    port map (
            O => \N__43515\,
            I => \N__43502\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__43512\,
            I => \N__43499\
        );

    \I__10062\ : CEMux
    port map (
            O => \N__43511\,
            I => \N__43496\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__43508\,
            I => \N__43493\
        );

    \I__10060\ : Span4Mux_h
    port map (
            O => \N__43505\,
            I => \N__43490\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__43502\,
            I => \N__43487\
        );

    \I__10058\ : Span4Mux_h
    port map (
            O => \N__43499\,
            I => \N__43480\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__43496\,
            I => \N__43480\
        );

    \I__10056\ : Span4Mux_h
    port map (
            O => \N__43493\,
            I => \N__43480\
        );

    \I__10055\ : Odrv4
    port map (
            O => \N__43490\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__10054\ : Odrv12
    port map (
            O => \N__43487\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__10053\ : Odrv4
    port map (
            O => \N__43480\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__10052\ : InMux
    port map (
            O => \N__43473\,
            I => \N__43455\
        );

    \I__10051\ : InMux
    port map (
            O => \N__43472\,
            I => \N__43455\
        );

    \I__10050\ : InMux
    port map (
            O => \N__43471\,
            I => \N__43455\
        );

    \I__10049\ : InMux
    port map (
            O => \N__43470\,
            I => \N__43455\
        );

    \I__10048\ : InMux
    port map (
            O => \N__43469\,
            I => \N__43455\
        );

    \I__10047\ : InMux
    port map (
            O => \N__43468\,
            I => \N__43455\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__43455\,
            I => \N__43439\
        );

    \I__10045\ : InMux
    port map (
            O => \N__43454\,
            I => \N__43430\
        );

    \I__10044\ : InMux
    port map (
            O => \N__43453\,
            I => \N__43430\
        );

    \I__10043\ : InMux
    port map (
            O => \N__43452\,
            I => \N__43430\
        );

    \I__10042\ : InMux
    port map (
            O => \N__43451\,
            I => \N__43430\
        );

    \I__10041\ : InMux
    port map (
            O => \N__43450\,
            I => \N__43425\
        );

    \I__10040\ : InMux
    port map (
            O => \N__43449\,
            I => \N__43412\
        );

    \I__10039\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43412\
        );

    \I__10038\ : InMux
    port map (
            O => \N__43447\,
            I => \N__43412\
        );

    \I__10037\ : InMux
    port map (
            O => \N__43446\,
            I => \N__43412\
        );

    \I__10036\ : InMux
    port map (
            O => \N__43445\,
            I => \N__43412\
        );

    \I__10035\ : InMux
    port map (
            O => \N__43444\,
            I => \N__43412\
        );

    \I__10034\ : InMux
    port map (
            O => \N__43443\,
            I => \N__43407\
        );

    \I__10033\ : InMux
    port map (
            O => \N__43442\,
            I => \N__43407\
        );

    \I__10032\ : Span4Mux_v
    port map (
            O => \N__43439\,
            I => \N__43402\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__43430\,
            I => \N__43402\
        );

    \I__10030\ : InMux
    port map (
            O => \N__43429\,
            I => \N__43398\
        );

    \I__10029\ : InMux
    port map (
            O => \N__43428\,
            I => \N__43393\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__43425\,
            I => \N__43390\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__43412\,
            I => \N__43387\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__43407\,
            I => \N__43382\
        );

    \I__10025\ : Span4Mux_h
    port map (
            O => \N__43402\,
            I => \N__43382\
        );

    \I__10024\ : InMux
    port map (
            O => \N__43401\,
            I => \N__43379\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__43398\,
            I => \N__43376\
        );

    \I__10022\ : InMux
    port map (
            O => \N__43397\,
            I => \N__43373\
        );

    \I__10021\ : InMux
    port map (
            O => \N__43396\,
            I => \N__43370\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__43393\,
            I => \N__43363\
        );

    \I__10019\ : Span4Mux_v
    port map (
            O => \N__43390\,
            I => \N__43363\
        );

    \I__10018\ : Span4Mux_v
    port map (
            O => \N__43387\,
            I => \N__43363\
        );

    \I__10017\ : Span4Mux_v
    port map (
            O => \N__43382\,
            I => \N__43358\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__43379\,
            I => \N__43358\
        );

    \I__10015\ : Span4Mux_h
    port map (
            O => \N__43376\,
            I => \N__43355\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__43373\,
            I => \N__43352\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__43370\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10012\ : Odrv4
    port map (
            O => \N__43363\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__43358\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10010\ : Odrv4
    port map (
            O => \N__43355\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10009\ : Odrv12
    port map (
            O => \N__43352\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10008\ : CascadeMux
    port map (
            O => \N__43341\,
            I => \N__43327\
        );

    \I__10007\ : CascadeMux
    port map (
            O => \N__43340\,
            I => \N__43324\
        );

    \I__10006\ : CascadeMux
    port map (
            O => \N__43339\,
            I => \N__43321\
        );

    \I__10005\ : CascadeMux
    port map (
            O => \N__43338\,
            I => \N__43318\
        );

    \I__10004\ : CascadeMux
    port map (
            O => \N__43337\,
            I => \N__43312\
        );

    \I__10003\ : CascadeMux
    port map (
            O => \N__43336\,
            I => \N__43308\
        );

    \I__10002\ : CascadeMux
    port map (
            O => \N__43335\,
            I => \N__43305\
        );

    \I__10001\ : CascadeMux
    port map (
            O => \N__43334\,
            I => \N__43302\
        );

    \I__10000\ : CascadeMux
    port map (
            O => \N__43333\,
            I => \N__43299\
        );

    \I__9999\ : CascadeMux
    port map (
            O => \N__43332\,
            I => \N__43296\
        );

    \I__9998\ : CascadeMux
    port map (
            O => \N__43331\,
            I => \N__43293\
        );

    \I__9997\ : InMux
    port map (
            O => \N__43330\,
            I => \N__43287\
        );

    \I__9996\ : InMux
    port map (
            O => \N__43327\,
            I => \N__43270\
        );

    \I__9995\ : InMux
    port map (
            O => \N__43324\,
            I => \N__43270\
        );

    \I__9994\ : InMux
    port map (
            O => \N__43321\,
            I => \N__43270\
        );

    \I__9993\ : InMux
    port map (
            O => \N__43318\,
            I => \N__43270\
        );

    \I__9992\ : InMux
    port map (
            O => \N__43317\,
            I => \N__43270\
        );

    \I__9991\ : InMux
    port map (
            O => \N__43316\,
            I => \N__43270\
        );

    \I__9990\ : InMux
    port map (
            O => \N__43315\,
            I => \N__43265\
        );

    \I__9989\ : InMux
    port map (
            O => \N__43312\,
            I => \N__43265\
        );

    \I__9988\ : InMux
    port map (
            O => \N__43311\,
            I => \N__43256\
        );

    \I__9987\ : InMux
    port map (
            O => \N__43308\,
            I => \N__43256\
        );

    \I__9986\ : InMux
    port map (
            O => \N__43305\,
            I => \N__43256\
        );

    \I__9985\ : InMux
    port map (
            O => \N__43302\,
            I => \N__43256\
        );

    \I__9984\ : InMux
    port map (
            O => \N__43299\,
            I => \N__43243\
        );

    \I__9983\ : InMux
    port map (
            O => \N__43296\,
            I => \N__43243\
        );

    \I__9982\ : InMux
    port map (
            O => \N__43293\,
            I => \N__43243\
        );

    \I__9981\ : InMux
    port map (
            O => \N__43292\,
            I => \N__43243\
        );

    \I__9980\ : InMux
    port map (
            O => \N__43291\,
            I => \N__43243\
        );

    \I__9979\ : InMux
    port map (
            O => \N__43290\,
            I => \N__43243\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__43287\,
            I => \N__43240\
        );

    \I__9977\ : InMux
    port map (
            O => \N__43286\,
            I => \N__43237\
        );

    \I__9976\ : InMux
    port map (
            O => \N__43285\,
            I => \N__43234\
        );

    \I__9975\ : CascadeMux
    port map (
            O => \N__43284\,
            I => \N__43231\
        );

    \I__9974\ : CascadeMux
    port map (
            O => \N__43283\,
            I => \N__43228\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__43270\,
            I => \N__43224\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__43265\,
            I => \N__43221\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__43256\,
            I => \N__43216\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__43243\,
            I => \N__43216\
        );

    \I__9969\ : Span4Mux_v
    port map (
            O => \N__43240\,
            I => \N__43211\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__43237\,
            I => \N__43211\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__43234\,
            I => \N__43208\
        );

    \I__9966\ : InMux
    port map (
            O => \N__43231\,
            I => \N__43205\
        );

    \I__9965\ : InMux
    port map (
            O => \N__43228\,
            I => \N__43200\
        );

    \I__9964\ : InMux
    port map (
            O => \N__43227\,
            I => \N__43200\
        );

    \I__9963\ : Span4Mux_v
    port map (
            O => \N__43224\,
            I => \N__43197\
        );

    \I__9962\ : Span4Mux_v
    port map (
            O => \N__43221\,
            I => \N__43194\
        );

    \I__9961\ : Span4Mux_v
    port map (
            O => \N__43216\,
            I => \N__43187\
        );

    \I__9960\ : Span4Mux_h
    port map (
            O => \N__43211\,
            I => \N__43187\
        );

    \I__9959\ : Span4Mux_h
    port map (
            O => \N__43208\,
            I => \N__43187\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__43205\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__43200\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__9956\ : Odrv4
    port map (
            O => \N__43197\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__9955\ : Odrv4
    port map (
            O => \N__43194\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__9954\ : Odrv4
    port map (
            O => \N__43187\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__9953\ : InMux
    port map (
            O => \N__43176\,
            I => \N__43173\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__43173\,
            I => \N__43169\
        );

    \I__9951\ : InMux
    port map (
            O => \N__43172\,
            I => \N__43166\
        );

    \I__9950\ : Span4Mux_v
    port map (
            O => \N__43169\,
            I => \N__43160\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__43166\,
            I => \N__43160\
        );

    \I__9948\ : InMux
    port map (
            O => \N__43165\,
            I => \N__43157\
        );

    \I__9947\ : Span4Mux_h
    port map (
            O => \N__43160\,
            I => \N__43152\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__43157\,
            I => \N__43149\
        );

    \I__9945\ : InMux
    port map (
            O => \N__43156\,
            I => \N__43146\
        );

    \I__9944\ : InMux
    port map (
            O => \N__43155\,
            I => \N__43143\
        );

    \I__9943\ : Span4Mux_v
    port map (
            O => \N__43152\,
            I => \N__43140\
        );

    \I__9942\ : Span4Mux_v
    port map (
            O => \N__43149\,
            I => \N__43133\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__43146\,
            I => \N__43133\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__43143\,
            I => \N__43133\
        );

    \I__9939\ : Odrv4
    port map (
            O => \N__43140\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9938\ : Odrv4
    port map (
            O => \N__43133\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9937\ : CascadeMux
    port map (
            O => \N__43128\,
            I => \N__43121\
        );

    \I__9936\ : CascadeMux
    port map (
            O => \N__43127\,
            I => \N__43118\
        );

    \I__9935\ : CascadeMux
    port map (
            O => \N__43126\,
            I => \N__43111\
        );

    \I__9934\ : CascadeMux
    port map (
            O => \N__43125\,
            I => \N__43105\
        );

    \I__9933\ : CascadeMux
    port map (
            O => \N__43124\,
            I => \N__43102\
        );

    \I__9932\ : InMux
    port map (
            O => \N__43121\,
            I => \N__43093\
        );

    \I__9931\ : InMux
    port map (
            O => \N__43118\,
            I => \N__43093\
        );

    \I__9930\ : InMux
    port map (
            O => \N__43117\,
            I => \N__43084\
        );

    \I__9929\ : InMux
    port map (
            O => \N__43116\,
            I => \N__43084\
        );

    \I__9928\ : InMux
    port map (
            O => \N__43115\,
            I => \N__43084\
        );

    \I__9927\ : InMux
    port map (
            O => \N__43114\,
            I => \N__43084\
        );

    \I__9926\ : InMux
    port map (
            O => \N__43111\,
            I => \N__43080\
        );

    \I__9925\ : InMux
    port map (
            O => \N__43110\,
            I => \N__43073\
        );

    \I__9924\ : InMux
    port map (
            O => \N__43109\,
            I => \N__43073\
        );

    \I__9923\ : InMux
    port map (
            O => \N__43108\,
            I => \N__43073\
        );

    \I__9922\ : InMux
    port map (
            O => \N__43105\,
            I => \N__43062\
        );

    \I__9921\ : InMux
    port map (
            O => \N__43102\,
            I => \N__43062\
        );

    \I__9920\ : InMux
    port map (
            O => \N__43101\,
            I => \N__43062\
        );

    \I__9919\ : InMux
    port map (
            O => \N__43100\,
            I => \N__43055\
        );

    \I__9918\ : InMux
    port map (
            O => \N__43099\,
            I => \N__43055\
        );

    \I__9917\ : InMux
    port map (
            O => \N__43098\,
            I => \N__43055\
        );

    \I__9916\ : LocalMux
    port map (
            O => \N__43093\,
            I => \N__43050\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__43084\,
            I => \N__43050\
        );

    \I__9914\ : InMux
    port map (
            O => \N__43083\,
            I => \N__43047\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__43080\,
            I => \N__43043\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__43073\,
            I => \N__43040\
        );

    \I__9911\ : InMux
    port map (
            O => \N__43072\,
            I => \N__43035\
        );

    \I__9910\ : InMux
    port map (
            O => \N__43071\,
            I => \N__43035\
        );

    \I__9909\ : InMux
    port map (
            O => \N__43070\,
            I => \N__43032\
        );

    \I__9908\ : InMux
    port map (
            O => \N__43069\,
            I => \N__43028\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__43062\,
            I => \N__43023\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__43055\,
            I => \N__43023\
        );

    \I__9905\ : Span4Mux_v
    port map (
            O => \N__43050\,
            I => \N__43018\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__43047\,
            I => \N__43018\
        );

    \I__9903\ : InMux
    port map (
            O => \N__43046\,
            I => \N__43015\
        );

    \I__9902\ : Span4Mux_h
    port map (
            O => \N__43043\,
            I => \N__43006\
        );

    \I__9901\ : Span4Mux_h
    port map (
            O => \N__43040\,
            I => \N__43006\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__43035\,
            I => \N__43006\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__43032\,
            I => \N__43006\
        );

    \I__9898\ : CascadeMux
    port map (
            O => \N__43031\,
            I => \N__43003\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__43028\,
            I => \N__43000\
        );

    \I__9896\ : Span4Mux_h
    port map (
            O => \N__43023\,
            I => \N__42997\
        );

    \I__9895\ : Span4Mux_v
    port map (
            O => \N__43018\,
            I => \N__42993\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__43015\,
            I => \N__42988\
        );

    \I__9893\ : Span4Mux_v
    port map (
            O => \N__43006\,
            I => \N__42988\
        );

    \I__9892\ : InMux
    port map (
            O => \N__43003\,
            I => \N__42985\
        );

    \I__9891\ : Span4Mux_v
    port map (
            O => \N__43000\,
            I => \N__42982\
        );

    \I__9890\ : Span4Mux_v
    port map (
            O => \N__42997\,
            I => \N__42979\
        );

    \I__9889\ : InMux
    port map (
            O => \N__42996\,
            I => \N__42976\
        );

    \I__9888\ : Span4Mux_h
    port map (
            O => \N__42993\,
            I => \N__42971\
        );

    \I__9887\ : Span4Mux_v
    port map (
            O => \N__42988\,
            I => \N__42971\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__42985\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9885\ : Odrv4
    port map (
            O => \N__42982\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9884\ : Odrv4
    port map (
            O => \N__42979\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__42976\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__42971\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9881\ : CascadeMux
    port map (
            O => \N__42960\,
            I => \N__42944\
        );

    \I__9880\ : CascadeMux
    port map (
            O => \N__42959\,
            I => \N__42940\
        );

    \I__9879\ : CascadeMux
    port map (
            O => \N__42958\,
            I => \N__42931\
        );

    \I__9878\ : CascadeMux
    port map (
            O => \N__42957\,
            I => \N__42928\
        );

    \I__9877\ : CascadeMux
    port map (
            O => \N__42956\,
            I => \N__42925\
        );

    \I__9876\ : CascadeMux
    port map (
            O => \N__42955\,
            I => \N__42922\
        );

    \I__9875\ : CascadeMux
    port map (
            O => \N__42954\,
            I => \N__42919\
        );

    \I__9874\ : InMux
    port map (
            O => \N__42953\,
            I => \N__42905\
        );

    \I__9873\ : InMux
    port map (
            O => \N__42952\,
            I => \N__42905\
        );

    \I__9872\ : InMux
    port map (
            O => \N__42951\,
            I => \N__42905\
        );

    \I__9871\ : InMux
    port map (
            O => \N__42950\,
            I => \N__42905\
        );

    \I__9870\ : InMux
    port map (
            O => \N__42949\,
            I => \N__42905\
        );

    \I__9869\ : InMux
    port map (
            O => \N__42948\,
            I => \N__42905\
        );

    \I__9868\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42902\
        );

    \I__9867\ : InMux
    port map (
            O => \N__42944\,
            I => \N__42899\
        );

    \I__9866\ : InMux
    port map (
            O => \N__42943\,
            I => \N__42896\
        );

    \I__9865\ : InMux
    port map (
            O => \N__42940\,
            I => \N__42889\
        );

    \I__9864\ : InMux
    port map (
            O => \N__42939\,
            I => \N__42889\
        );

    \I__9863\ : InMux
    port map (
            O => \N__42938\,
            I => \N__42889\
        );

    \I__9862\ : InMux
    port map (
            O => \N__42937\,
            I => \N__42872\
        );

    \I__9861\ : InMux
    port map (
            O => \N__42936\,
            I => \N__42872\
        );

    \I__9860\ : InMux
    port map (
            O => \N__42935\,
            I => \N__42872\
        );

    \I__9859\ : InMux
    port map (
            O => \N__42934\,
            I => \N__42872\
        );

    \I__9858\ : InMux
    port map (
            O => \N__42931\,
            I => \N__42872\
        );

    \I__9857\ : InMux
    port map (
            O => \N__42928\,
            I => \N__42872\
        );

    \I__9856\ : InMux
    port map (
            O => \N__42925\,
            I => \N__42872\
        );

    \I__9855\ : InMux
    port map (
            O => \N__42922\,
            I => \N__42872\
        );

    \I__9854\ : InMux
    port map (
            O => \N__42919\,
            I => \N__42867\
        );

    \I__9853\ : InMux
    port map (
            O => \N__42918\,
            I => \N__42867\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__42905\,
            I => \N__42864\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__42902\,
            I => \N__42859\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__42899\,
            I => \N__42859\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__42896\,
            I => \N__42856\
        );

    \I__9848\ : LocalMux
    port map (
            O => \N__42889\,
            I => \N__42853\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__42872\,
            I => \N__42850\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__42867\,
            I => \N__42839\
        );

    \I__9845\ : Span4Mux_h
    port map (
            O => \N__42864\,
            I => \N__42839\
        );

    \I__9844\ : Span4Mux_v
    port map (
            O => \N__42859\,
            I => \N__42839\
        );

    \I__9843\ : Span4Mux_v
    port map (
            O => \N__42856\,
            I => \N__42839\
        );

    \I__9842\ : Span4Mux_h
    port map (
            O => \N__42853\,
            I => \N__42834\
        );

    \I__9841\ : Span4Mux_h
    port map (
            O => \N__42850\,
            I => \N__42834\
        );

    \I__9840\ : InMux
    port map (
            O => \N__42849\,
            I => \N__42831\
        );

    \I__9839\ : InMux
    port map (
            O => \N__42848\,
            I => \N__42828\
        );

    \I__9838\ : Odrv4
    port map (
            O => \N__42839\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9837\ : Odrv4
    port map (
            O => \N__42834\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__42831\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__42828\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__42819\,
            I => \N__42816\
        );

    \I__9833\ : InMux
    port map (
            O => \N__42816\,
            I => \N__42809\
        );

    \I__9832\ : InMux
    port map (
            O => \N__42815\,
            I => \N__42798\
        );

    \I__9831\ : InMux
    port map (
            O => \N__42814\,
            I => \N__42798\
        );

    \I__9830\ : InMux
    port map (
            O => \N__42813\,
            I => \N__42798\
        );

    \I__9829\ : InMux
    port map (
            O => \N__42812\,
            I => \N__42794\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__42809\,
            I => \N__42782\
        );

    \I__9827\ : CascadeMux
    port map (
            O => \N__42808\,
            I => \N__42777\
        );

    \I__9826\ : CascadeMux
    port map (
            O => \N__42807\,
            I => \N__42772\
        );

    \I__9825\ : CascadeMux
    port map (
            O => \N__42806\,
            I => \N__42769\
        );

    \I__9824\ : CascadeMux
    port map (
            O => \N__42805\,
            I => \N__42766\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__42798\,
            I => \N__42763\
        );

    \I__9822\ : InMux
    port map (
            O => \N__42797\,
            I => \N__42760\
        );

    \I__9821\ : LocalMux
    port map (
            O => \N__42794\,
            I => \N__42757\
        );

    \I__9820\ : InMux
    port map (
            O => \N__42793\,
            I => \N__42754\
        );

    \I__9819\ : InMux
    port map (
            O => \N__42792\,
            I => \N__42736\
        );

    \I__9818\ : InMux
    port map (
            O => \N__42791\,
            I => \N__42736\
        );

    \I__9817\ : InMux
    port map (
            O => \N__42790\,
            I => \N__42736\
        );

    \I__9816\ : InMux
    port map (
            O => \N__42789\,
            I => \N__42736\
        );

    \I__9815\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42736\
        );

    \I__9814\ : InMux
    port map (
            O => \N__42787\,
            I => \N__42736\
        );

    \I__9813\ : InMux
    port map (
            O => \N__42786\,
            I => \N__42736\
        );

    \I__9812\ : InMux
    port map (
            O => \N__42785\,
            I => \N__42736\
        );

    \I__9811\ : Span4Mux_v
    port map (
            O => \N__42782\,
            I => \N__42733\
        );

    \I__9810\ : InMux
    port map (
            O => \N__42781\,
            I => \N__42730\
        );

    \I__9809\ : InMux
    port map (
            O => \N__42780\,
            I => \N__42725\
        );

    \I__9808\ : InMux
    port map (
            O => \N__42777\,
            I => \N__42725\
        );

    \I__9807\ : InMux
    port map (
            O => \N__42776\,
            I => \N__42714\
        );

    \I__9806\ : InMux
    port map (
            O => \N__42775\,
            I => \N__42714\
        );

    \I__9805\ : InMux
    port map (
            O => \N__42772\,
            I => \N__42714\
        );

    \I__9804\ : InMux
    port map (
            O => \N__42769\,
            I => \N__42714\
        );

    \I__9803\ : InMux
    port map (
            O => \N__42766\,
            I => \N__42714\
        );

    \I__9802\ : Span4Mux_v
    port map (
            O => \N__42763\,
            I => \N__42711\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__42760\,
            I => \N__42704\
        );

    \I__9800\ : Span4Mux_v
    port map (
            O => \N__42757\,
            I => \N__42704\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__42754\,
            I => \N__42704\
        );

    \I__9798\ : InMux
    port map (
            O => \N__42753\,
            I => \N__42701\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__42736\,
            I => \N__42694\
        );

    \I__9796\ : Span4Mux_h
    port map (
            O => \N__42733\,
            I => \N__42694\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__42730\,
            I => \N__42694\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__42725\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__42714\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9792\ : Odrv4
    port map (
            O => \N__42711\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9791\ : Odrv4
    port map (
            O => \N__42704\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__42701\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9789\ : Odrv4
    port map (
            O => \N__42694\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9788\ : InMux
    port map (
            O => \N__42681\,
            I => \N__42677\
        );

    \I__9787\ : InMux
    port map (
            O => \N__42680\,
            I => \N__42674\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__42677\,
            I => \N__42669\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__42674\,
            I => \N__42666\
        );

    \I__9784\ : InMux
    port map (
            O => \N__42673\,
            I => \N__42663\
        );

    \I__9783\ : InMux
    port map (
            O => \N__42672\,
            I => \N__42660\
        );

    \I__9782\ : Span4Mux_v
    port map (
            O => \N__42669\,
            I => \N__42655\
        );

    \I__9781\ : Span12Mux_v
    port map (
            O => \N__42666\,
            I => \N__42652\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__42663\,
            I => \N__42649\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__42660\,
            I => \N__42646\
        );

    \I__9778\ : InMux
    port map (
            O => \N__42659\,
            I => \N__42641\
        );

    \I__9777\ : InMux
    port map (
            O => \N__42658\,
            I => \N__42641\
        );

    \I__9776\ : Odrv4
    port map (
            O => \N__42655\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9775\ : Odrv12
    port map (
            O => \N__42652\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9774\ : Odrv4
    port map (
            O => \N__42649\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9773\ : Odrv4
    port map (
            O => \N__42646\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__42641\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9771\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42614\
        );

    \I__9770\ : InMux
    port map (
            O => \N__42629\,
            I => \N__42611\
        );

    \I__9769\ : InMux
    port map (
            O => \N__42628\,
            I => \N__42600\
        );

    \I__9768\ : InMux
    port map (
            O => \N__42627\,
            I => \N__42585\
        );

    \I__9767\ : InMux
    port map (
            O => \N__42626\,
            I => \N__42585\
        );

    \I__9766\ : InMux
    port map (
            O => \N__42625\,
            I => \N__42585\
        );

    \I__9765\ : InMux
    port map (
            O => \N__42624\,
            I => \N__42585\
        );

    \I__9764\ : InMux
    port map (
            O => \N__42623\,
            I => \N__42585\
        );

    \I__9763\ : InMux
    port map (
            O => \N__42622\,
            I => \N__42585\
        );

    \I__9762\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42585\
        );

    \I__9761\ : InMux
    port map (
            O => \N__42620\,
            I => \N__42582\
        );

    \I__9760\ : InMux
    port map (
            O => \N__42619\,
            I => \N__42574\
        );

    \I__9759\ : InMux
    port map (
            O => \N__42618\,
            I => \N__42574\
        );

    \I__9758\ : InMux
    port map (
            O => \N__42617\,
            I => \N__42574\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__42614\,
            I => \N__42569\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__42611\,
            I => \N__42569\
        );

    \I__9755\ : InMux
    port map (
            O => \N__42610\,
            I => \N__42552\
        );

    \I__9754\ : InMux
    port map (
            O => \N__42609\,
            I => \N__42552\
        );

    \I__9753\ : InMux
    port map (
            O => \N__42608\,
            I => \N__42552\
        );

    \I__9752\ : InMux
    port map (
            O => \N__42607\,
            I => \N__42552\
        );

    \I__9751\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42552\
        );

    \I__9750\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42552\
        );

    \I__9749\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42552\
        );

    \I__9748\ : InMux
    port map (
            O => \N__42603\,
            I => \N__42552\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__42600\,
            I => \N__42549\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__42585\,
            I => \N__42544\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__42582\,
            I => \N__42544\
        );

    \I__9744\ : InMux
    port map (
            O => \N__42581\,
            I => \N__42541\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__42574\,
            I => \N__42535\
        );

    \I__9742\ : Span4Mux_h
    port map (
            O => \N__42569\,
            I => \N__42535\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__42552\,
            I => \N__42526\
        );

    \I__9740\ : Span4Mux_h
    port map (
            O => \N__42549\,
            I => \N__42526\
        );

    \I__9739\ : Span4Mux_v
    port map (
            O => \N__42544\,
            I => \N__42526\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__42541\,
            I => \N__42526\
        );

    \I__9737\ : InMux
    port map (
            O => \N__42540\,
            I => \N__42523\
        );

    \I__9736\ : Span4Mux_v
    port map (
            O => \N__42535\,
            I => \N__42520\
        );

    \I__9735\ : Span4Mux_v
    port map (
            O => \N__42526\,
            I => \N__42517\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__42523\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__9733\ : Odrv4
    port map (
            O => \N__42520\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__9732\ : Odrv4
    port map (
            O => \N__42517\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__9731\ : CEMux
    port map (
            O => \N__42510\,
            I => \N__42503\
        );

    \I__9730\ : CEMux
    port map (
            O => \N__42509\,
            I => \N__42499\
        );

    \I__9729\ : CEMux
    port map (
            O => \N__42508\,
            I => \N__42496\
        );

    \I__9728\ : CEMux
    port map (
            O => \N__42507\,
            I => \N__42493\
        );

    \I__9727\ : IoInMux
    port map (
            O => \N__42506\,
            I => \N__42490\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__42503\,
            I => \N__42487\
        );

    \I__9725\ : CEMux
    port map (
            O => \N__42502\,
            I => \N__42484\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__42499\,
            I => \N__42481\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__42496\,
            I => \N__42478\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__42493\,
            I => \N__42475\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__42490\,
            I => \N__42472\
        );

    \I__9720\ : Span4Mux_v
    port map (
            O => \N__42487\,
            I => \N__42469\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__42484\,
            I => \N__42466\
        );

    \I__9718\ : Span12Mux_h
    port map (
            O => \N__42481\,
            I => \N__42463\
        );

    \I__9717\ : Span12Mux_s10_v
    port map (
            O => \N__42478\,
            I => \N__42458\
        );

    \I__9716\ : Sp12to4
    port map (
            O => \N__42475\,
            I => \N__42458\
        );

    \I__9715\ : Span4Mux_s3_v
    port map (
            O => \N__42472\,
            I => \N__42455\
        );

    \I__9714\ : Span4Mux_v
    port map (
            O => \N__42469\,
            I => \N__42452\
        );

    \I__9713\ : Span4Mux_v
    port map (
            O => \N__42466\,
            I => \N__42449\
        );

    \I__9712\ : Span12Mux_v
    port map (
            O => \N__42463\,
            I => \N__42446\
        );

    \I__9711\ : Span12Mux_v
    port map (
            O => \N__42458\,
            I => \N__42443\
        );

    \I__9710\ : Span4Mux_v
    port map (
            O => \N__42455\,
            I => \N__42440\
        );

    \I__9709\ : Span4Mux_v
    port map (
            O => \N__42452\,
            I => \N__42437\
        );

    \I__9708\ : Span4Mux_v
    port map (
            O => \N__42449\,
            I => \N__42434\
        );

    \I__9707\ : Odrv12
    port map (
            O => \N__42446\,
            I => red_c_i
        );

    \I__9706\ : Odrv12
    port map (
            O => \N__42443\,
            I => red_c_i
        );

    \I__9705\ : Odrv4
    port map (
            O => \N__42440\,
            I => red_c_i
        );

    \I__9704\ : Odrv4
    port map (
            O => \N__42437\,
            I => red_c_i
        );

    \I__9703\ : Odrv4
    port map (
            O => \N__42434\,
            I => red_c_i
        );

    \I__9702\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42419\
        );

    \I__9701\ : InMux
    port map (
            O => \N__42422\,
            I => \N__42416\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__42419\,
            I => \N__42411\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__42416\,
            I => \N__42411\
        );

    \I__9698\ : Span4Mux_v
    port map (
            O => \N__42411\,
            I => \N__42408\
        );

    \I__9697\ : Odrv4
    port map (
            O => \N__42408\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__9696\ : CascadeMux
    port map (
            O => \N__42405\,
            I => \N__42402\
        );

    \I__9695\ : InMux
    port map (
            O => \N__42402\,
            I => \N__42397\
        );

    \I__9694\ : InMux
    port map (
            O => \N__42401\,
            I => \N__42394\
        );

    \I__9693\ : CascadeMux
    port map (
            O => \N__42400\,
            I => \N__42391\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__42397\,
            I => \N__42388\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__42394\,
            I => \N__42385\
        );

    \I__9690\ : InMux
    port map (
            O => \N__42391\,
            I => \N__42382\
        );

    \I__9689\ : Span4Mux_h
    port map (
            O => \N__42388\,
            I => \N__42379\
        );

    \I__9688\ : Odrv4
    port map (
            O => \N__42385\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__42382\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__9686\ : Odrv4
    port map (
            O => \N__42379\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__9685\ : InMux
    port map (
            O => \N__42372\,
            I => \N__42368\
        );

    \I__9684\ : InMux
    port map (
            O => \N__42371\,
            I => \N__42365\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__42368\,
            I => \N__42362\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__42365\,
            I => \N__42359\
        );

    \I__9681\ : Span4Mux_v
    port map (
            O => \N__42362\,
            I => \N__42353\
        );

    \I__9680\ : Span4Mux_h
    port map (
            O => \N__42359\,
            I => \N__42353\
        );

    \I__9679\ : InMux
    port map (
            O => \N__42358\,
            I => \N__42350\
        );

    \I__9678\ : Odrv4
    port map (
            O => \N__42353\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__42350\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__9676\ : InMux
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__42342\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_3\
        );

    \I__9674\ : InMux
    port map (
            O => \N__42339\,
            I => \N__42336\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__42336\,
            I => \N__42332\
        );

    \I__9672\ : InMux
    port map (
            O => \N__42335\,
            I => \N__42329\
        );

    \I__9671\ : Span4Mux_v
    port map (
            O => \N__42332\,
            I => \N__42326\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__42329\,
            I => \N__42323\
        );

    \I__9669\ : Odrv4
    port map (
            O => \N__42326\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__9668\ : Odrv4
    port map (
            O => \N__42323\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__9667\ : InMux
    port map (
            O => \N__42318\,
            I => \N__42314\
        );

    \I__9666\ : InMux
    port map (
            O => \N__42317\,
            I => \N__42311\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__42314\,
            I => \delay_measurement_inst.N_332\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__42311\,
            I => \delay_measurement_inst.N_332\
        );

    \I__9663\ : InMux
    port map (
            O => \N__42306\,
            I => \N__42302\
        );

    \I__9662\ : InMux
    port map (
            O => \N__42305\,
            I => \N__42299\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__42302\,
            I => \delay_measurement_inst.N_318\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__42299\,
            I => \delay_measurement_inst.N_318\
        );

    \I__9659\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42291\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__42291\,
            I => \N__42288\
        );

    \I__9657\ : Odrv12
    port map (
            O => \N__42288\,
            I => \delay_measurement_inst.N_295\
        );

    \I__9656\ : InMux
    port map (
            O => \N__42285\,
            I => \N__42282\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__42282\,
            I => \N__42279\
        );

    \I__9654\ : Span4Mux_h
    port map (
            O => \N__42279\,
            I => \N__42273\
        );

    \I__9653\ : InMux
    port map (
            O => \N__42278\,
            I => \N__42266\
        );

    \I__9652\ : InMux
    port map (
            O => \N__42277\,
            I => \N__42266\
        );

    \I__9651\ : InMux
    port map (
            O => \N__42276\,
            I => \N__42266\
        );

    \I__9650\ : Odrv4
    port map (
            O => \N__42273\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__42266\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__9648\ : InMux
    port map (
            O => \N__42261\,
            I => \N__42253\
        );

    \I__9647\ : InMux
    port map (
            O => \N__42260\,
            I => \N__42250\
        );

    \I__9646\ : InMux
    port map (
            O => \N__42259\,
            I => \N__42247\
        );

    \I__9645\ : InMux
    port map (
            O => \N__42258\,
            I => \N__42242\
        );

    \I__9644\ : InMux
    port map (
            O => \N__42257\,
            I => \N__42242\
        );

    \I__9643\ : CascadeMux
    port map (
            O => \N__42256\,
            I => \N__42239\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__42253\,
            I => \N__42232\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__42250\,
            I => \N__42232\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__42247\,
            I => \N__42232\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__42242\,
            I => \N__42229\
        );

    \I__9638\ : InMux
    port map (
            O => \N__42239\,
            I => \N__42226\
        );

    \I__9637\ : Sp12to4
    port map (
            O => \N__42232\,
            I => \N__42223\
        );

    \I__9636\ : Span4Mux_h
    port map (
            O => \N__42229\,
            I => \N__42220\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__42226\,
            I => measured_delay_hc_15
        );

    \I__9634\ : Odrv12
    port map (
            O => \N__42223\,
            I => measured_delay_hc_15
        );

    \I__9633\ : Odrv4
    port map (
            O => \N__42220\,
            I => measured_delay_hc_15
        );

    \I__9632\ : CascadeMux
    port map (
            O => \N__42213\,
            I => \N__42210\
        );

    \I__9631\ : InMux
    port map (
            O => \N__42210\,
            I => \N__42207\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__42207\,
            I => \N__42204\
        );

    \I__9629\ : Span4Mux_h
    port map (
            O => \N__42204\,
            I => \N__42201\
        );

    \I__9628\ : Odrv4
    port map (
            O => \N__42201\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\
        );

    \I__9627\ : InMux
    port map (
            O => \N__42198\,
            I => \N__42194\
        );

    \I__9626\ : InMux
    port map (
            O => \N__42197\,
            I => \N__42191\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__42194\,
            I => \N__42188\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__42191\,
            I => \N__42185\
        );

    \I__9623\ : Span4Mux_v
    port map (
            O => \N__42188\,
            I => \N__42182\
        );

    \I__9622\ : Span4Mux_v
    port map (
            O => \N__42185\,
            I => \N__42179\
        );

    \I__9621\ : Span4Mux_h
    port map (
            O => \N__42182\,
            I => \N__42176\
        );

    \I__9620\ : Span4Mux_h
    port map (
            O => \N__42179\,
            I => \N__42173\
        );

    \I__9619\ : Odrv4
    port map (
            O => \N__42176\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__9618\ : Odrv4
    port map (
            O => \N__42173\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__9617\ : InMux
    port map (
            O => \N__42168\,
            I => \N__42165\
        );

    \I__9616\ : LocalMux
    port map (
            O => \N__42165\,
            I => \N__42162\
        );

    \I__9615\ : Span4Mux_h
    port map (
            O => \N__42162\,
            I => \N__42159\
        );

    \I__9614\ : Odrv4
    port map (
            O => \N__42159\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\
        );

    \I__9613\ : InMux
    port map (
            O => \N__42156\,
            I => \N__42152\
        );

    \I__9612\ : InMux
    port map (
            O => \N__42155\,
            I => \N__42149\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__42152\,
            I => \N__42146\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__42149\,
            I => \N__42143\
        );

    \I__9609\ : Span4Mux_v
    port map (
            O => \N__42146\,
            I => \N__42140\
        );

    \I__9608\ : Span12Mux_s8_v
    port map (
            O => \N__42143\,
            I => \N__42137\
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__42140\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__9606\ : Odrv12
    port map (
            O => \N__42137\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__42132\,
            I => \N__42129\
        );

    \I__9604\ : InMux
    port map (
            O => \N__42129\,
            I => \N__42126\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__42126\,
            I => \N__42123\
        );

    \I__9602\ : Odrv12
    port map (
            O => \N__42123\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\
        );

    \I__9601\ : InMux
    port map (
            O => \N__42120\,
            I => \N__42116\
        );

    \I__9600\ : InMux
    port map (
            O => \N__42119\,
            I => \N__42113\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__42116\,
            I => \N__42108\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__42113\,
            I => \N__42108\
        );

    \I__9597\ : Odrv12
    port map (
            O => \N__42108\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__9596\ : CascadeMux
    port map (
            O => \N__42105\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__9595\ : InMux
    port map (
            O => \N__42102\,
            I => \N__42098\
        );

    \I__9594\ : InMux
    port map (
            O => \N__42101\,
            I => \N__42095\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__42098\,
            I => measured_delay_hc_27
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__42095\,
            I => measured_delay_hc_27
        );

    \I__9591\ : InMux
    port map (
            O => \N__42090\,
            I => \N__42086\
        );

    \I__9590\ : InMux
    port map (
            O => \N__42089\,
            I => \N__42083\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__42086\,
            I => measured_delay_hc_28
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__42083\,
            I => measured_delay_hc_28
        );

    \I__9587\ : InMux
    port map (
            O => \N__42078\,
            I => \N__42073\
        );

    \I__9586\ : InMux
    port map (
            O => \N__42077\,
            I => \N__42070\
        );

    \I__9585\ : InMux
    port map (
            O => \N__42076\,
            I => \N__42067\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__42073\,
            I => \N__42063\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__42070\,
            I => \N__42058\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__42067\,
            I => \N__42058\
        );

    \I__9581\ : InMux
    port map (
            O => \N__42066\,
            I => \N__42055\
        );

    \I__9580\ : Span4Mux_h
    port map (
            O => \N__42063\,
            I => \N__42050\
        );

    \I__9579\ : Span4Mux_v
    port map (
            O => \N__42058\,
            I => \N__42050\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__42055\,
            I => measured_delay_hc_0
        );

    \I__9577\ : Odrv4
    port map (
            O => \N__42050\,
            I => measured_delay_hc_0
        );

    \I__9576\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42041\
        );

    \I__9575\ : CascadeMux
    port map (
            O => \N__42044\,
            I => \N__42037\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__42041\,
            I => \N__42034\
        );

    \I__9573\ : InMux
    port map (
            O => \N__42040\,
            I => \N__42031\
        );

    \I__9572\ : InMux
    port map (
            O => \N__42037\,
            I => \N__42028\
        );

    \I__9571\ : Span4Mux_v
    port map (
            O => \N__42034\,
            I => \N__42025\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__42031\,
            I => \N__42022\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__42028\,
            I => \N__42019\
        );

    \I__9568\ : Span4Mux_h
    port map (
            O => \N__42025\,
            I => \N__42014\
        );

    \I__9567\ : Span4Mux_v
    port map (
            O => \N__42022\,
            I => \N__42014\
        );

    \I__9566\ : Span4Mux_h
    port map (
            O => \N__42019\,
            I => \N__42011\
        );

    \I__9565\ : Odrv4
    port map (
            O => \N__42014\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__9564\ : Odrv4
    port map (
            O => \N__42011\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__9563\ : CascadeMux
    port map (
            O => \N__42006\,
            I => \N__42002\
        );

    \I__9562\ : CascadeMux
    port map (
            O => \N__42005\,
            I => \N__41999\
        );

    \I__9561\ : InMux
    port map (
            O => \N__42002\,
            I => \N__41994\
        );

    \I__9560\ : InMux
    port map (
            O => \N__41999\,
            I => \N__41991\
        );

    \I__9559\ : CascadeMux
    port map (
            O => \N__41998\,
            I => \N__41987\
        );

    \I__9558\ : InMux
    port map (
            O => \N__41997\,
            I => \N__41984\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__41994\,
            I => \N__41981\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__41991\,
            I => \N__41978\
        );

    \I__9555\ : InMux
    port map (
            O => \N__41990\,
            I => \N__41975\
        );

    \I__9554\ : InMux
    port map (
            O => \N__41987\,
            I => \N__41972\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__41984\,
            I => measured_delay_hc_19
        );

    \I__9552\ : Odrv12
    port map (
            O => \N__41981\,
            I => measured_delay_hc_19
        );

    \I__9551\ : Odrv4
    port map (
            O => \N__41978\,
            I => measured_delay_hc_19
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__41975\,
            I => measured_delay_hc_19
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__41972\,
            I => measured_delay_hc_19
        );

    \I__9548\ : InMux
    port map (
            O => \N__41961\,
            I => \N__41958\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__41958\,
            I => \N__41955\
        );

    \I__9546\ : Span4Mux_h
    port map (
            O => \N__41955\,
            I => \N__41950\
        );

    \I__9545\ : InMux
    port map (
            O => \N__41954\,
            I => \N__41945\
        );

    \I__9544\ : InMux
    port map (
            O => \N__41953\,
            I => \N__41945\
        );

    \I__9543\ : Odrv4
    port map (
            O => \N__41950\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__41945\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__9541\ : InMux
    port map (
            O => \N__41940\,
            I => \N__41937\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__41937\,
            I => \N__41931\
        );

    \I__9539\ : InMux
    port map (
            O => \N__41936\,
            I => \N__41928\
        );

    \I__9538\ : InMux
    port map (
            O => \N__41935\,
            I => \N__41925\
        );

    \I__9537\ : InMux
    port map (
            O => \N__41934\,
            I => \N__41922\
        );

    \I__9536\ : Span4Mux_h
    port map (
            O => \N__41931\,
            I => \N__41918\
        );

    \I__9535\ : LocalMux
    port map (
            O => \N__41928\,
            I => \N__41911\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__41925\,
            I => \N__41911\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__41922\,
            I => \N__41911\
        );

    \I__9532\ : InMux
    port map (
            O => \N__41921\,
            I => \N__41908\
        );

    \I__9531\ : Span4Mux_v
    port map (
            O => \N__41918\,
            I => \N__41905\
        );

    \I__9530\ : Span4Mux_v
    port map (
            O => \N__41911\,
            I => \N__41902\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__41908\,
            I => measured_delay_hc_1
        );

    \I__9528\ : Odrv4
    port map (
            O => \N__41905\,
            I => measured_delay_hc_1
        );

    \I__9527\ : Odrv4
    port map (
            O => \N__41902\,
            I => measured_delay_hc_1
        );

    \I__9526\ : CascadeMux
    port map (
            O => \N__41895\,
            I => \N__41892\
        );

    \I__9525\ : InMux
    port map (
            O => \N__41892\,
            I => \N__41889\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__41889\,
            I => \N__41886\
        );

    \I__9523\ : Span4Mux_h
    port map (
            O => \N__41886\,
            I => \N__41881\
        );

    \I__9522\ : InMux
    port map (
            O => \N__41885\,
            I => \N__41878\
        );

    \I__9521\ : InMux
    port map (
            O => \N__41884\,
            I => \N__41875\
        );

    \I__9520\ : Odrv4
    port map (
            O => \N__41881\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__41878\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__41875\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__9517\ : InMux
    port map (
            O => \N__41868\,
            I => \N__41863\
        );

    \I__9516\ : InMux
    port map (
            O => \N__41867\,
            I => \N__41860\
        );

    \I__9515\ : InMux
    port map (
            O => \N__41866\,
            I => \N__41855\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__41863\,
            I => \N__41850\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__41860\,
            I => \N__41850\
        );

    \I__9512\ : InMux
    port map (
            O => \N__41859\,
            I => \N__41847\
        );

    \I__9511\ : InMux
    port map (
            O => \N__41858\,
            I => \N__41844\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__41855\,
            I => \N__41841\
        );

    \I__9509\ : Span4Mux_v
    port map (
            O => \N__41850\,
            I => \N__41836\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__41847\,
            I => \N__41836\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__41844\,
            I => measured_delay_hc_18
        );

    \I__9506\ : Odrv4
    port map (
            O => \N__41841\,
            I => measured_delay_hc_18
        );

    \I__9505\ : Odrv4
    port map (
            O => \N__41836\,
            I => measured_delay_hc_18
        );

    \I__9504\ : InMux
    port map (
            O => \N__41829\,
            I => \N__41824\
        );

    \I__9503\ : InMux
    port map (
            O => \N__41828\,
            I => \N__41821\
        );

    \I__9502\ : CascadeMux
    port map (
            O => \N__41827\,
            I => \N__41818\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__41824\,
            I => \N__41811\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__41821\,
            I => \N__41811\
        );

    \I__9499\ : InMux
    port map (
            O => \N__41818\,
            I => \N__41808\
        );

    \I__9498\ : CascadeMux
    port map (
            O => \N__41817\,
            I => \N__41805\
        );

    \I__9497\ : InMux
    port map (
            O => \N__41816\,
            I => \N__41802\
        );

    \I__9496\ : Span4Mux_v
    port map (
            O => \N__41811\,
            I => \N__41797\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__41808\,
            I => \N__41797\
        );

    \I__9494\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41794\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__41802\,
            I => \N__41791\
        );

    \I__9492\ : Span4Mux_h
    port map (
            O => \N__41797\,
            I => \N__41788\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__41794\,
            I => measured_delay_hc_13
        );

    \I__9490\ : Odrv4
    port map (
            O => \N__41791\,
            I => measured_delay_hc_13
        );

    \I__9489\ : Odrv4
    port map (
            O => \N__41788\,
            I => measured_delay_hc_13
        );

    \I__9488\ : CascadeMux
    port map (
            O => \N__41781\,
            I => \N__41775\
        );

    \I__9487\ : CascadeMux
    port map (
            O => \N__41780\,
            I => \N__41772\
        );

    \I__9486\ : CascadeMux
    port map (
            O => \N__41779\,
            I => \N__41765\
        );

    \I__9485\ : InMux
    port map (
            O => \N__41778\,
            I => \N__41754\
        );

    \I__9484\ : InMux
    port map (
            O => \N__41775\,
            I => \N__41754\
        );

    \I__9483\ : InMux
    port map (
            O => \N__41772\,
            I => \N__41754\
        );

    \I__9482\ : InMux
    port map (
            O => \N__41771\,
            I => \N__41754\
        );

    \I__9481\ : CascadeMux
    port map (
            O => \N__41770\,
            I => \N__41743\
        );

    \I__9480\ : CascadeMux
    port map (
            O => \N__41769\,
            I => \N__41740\
        );

    \I__9479\ : CascadeMux
    port map (
            O => \N__41768\,
            I => \N__41737\
        );

    \I__9478\ : InMux
    port map (
            O => \N__41765\,
            I => \N__41726\
        );

    \I__9477\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41726\
        );

    \I__9476\ : InMux
    port map (
            O => \N__41763\,
            I => \N__41726\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__41754\,
            I => \N__41723\
        );

    \I__9474\ : InMux
    port map (
            O => \N__41753\,
            I => \N__41708\
        );

    \I__9473\ : InMux
    port map (
            O => \N__41752\,
            I => \N__41708\
        );

    \I__9472\ : InMux
    port map (
            O => \N__41751\,
            I => \N__41708\
        );

    \I__9471\ : InMux
    port map (
            O => \N__41750\,
            I => \N__41708\
        );

    \I__9470\ : InMux
    port map (
            O => \N__41749\,
            I => \N__41708\
        );

    \I__9469\ : InMux
    port map (
            O => \N__41748\,
            I => \N__41708\
        );

    \I__9468\ : InMux
    port map (
            O => \N__41747\,
            I => \N__41708\
        );

    \I__9467\ : InMux
    port map (
            O => \N__41746\,
            I => \N__41699\
        );

    \I__9466\ : InMux
    port map (
            O => \N__41743\,
            I => \N__41699\
        );

    \I__9465\ : InMux
    port map (
            O => \N__41740\,
            I => \N__41699\
        );

    \I__9464\ : InMux
    port map (
            O => \N__41737\,
            I => \N__41699\
        );

    \I__9463\ : InMux
    port map (
            O => \N__41736\,
            I => \N__41690\
        );

    \I__9462\ : InMux
    port map (
            O => \N__41735\,
            I => \N__41690\
        );

    \I__9461\ : InMux
    port map (
            O => \N__41734\,
            I => \N__41690\
        );

    \I__9460\ : InMux
    port map (
            O => \N__41733\,
            I => \N__41690\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__41726\,
            I => \N__41687\
        );

    \I__9458\ : Span4Mux_h
    port map (
            O => \N__41723\,
            I => \N__41684\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__41708\,
            I => \N__41681\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__41699\,
            I => \phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__41690\,
            I => \phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0\
        );

    \I__9454\ : Odrv4
    port map (
            O => \N__41687\,
            I => \phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0\
        );

    \I__9453\ : Odrv4
    port map (
            O => \N__41684\,
            I => \phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0\
        );

    \I__9452\ : Odrv12
    port map (
            O => \N__41681\,
            I => \phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0\
        );

    \I__9451\ : InMux
    port map (
            O => \N__41670\,
            I => \N__41665\
        );

    \I__9450\ : InMux
    port map (
            O => \N__41669\,
            I => \N__41660\
        );

    \I__9449\ : InMux
    port map (
            O => \N__41668\,
            I => \N__41660\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__41665\,
            I => \phase_controller_inst1.stoper_hc.N_459\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__41660\,
            I => \phase_controller_inst1.stoper_hc.N_459\
        );

    \I__9446\ : CascadeMux
    port map (
            O => \N__41655\,
            I => \N__41652\
        );

    \I__9445\ : InMux
    port map (
            O => \N__41652\,
            I => \N__41649\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__41649\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3\
        );

    \I__9443\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41641\
        );

    \I__9442\ : InMux
    port map (
            O => \N__41645\,
            I => \N__41638\
        );

    \I__9441\ : InMux
    port map (
            O => \N__41644\,
            I => \N__41634\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__41641\,
            I => \N__41629\
        );

    \I__9439\ : LocalMux
    port map (
            O => \N__41638\,
            I => \N__41629\
        );

    \I__9438\ : InMux
    port map (
            O => \N__41637\,
            I => \N__41626\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__41634\,
            I => \N__41623\
        );

    \I__9436\ : Span4Mux_v
    port map (
            O => \N__41629\,
            I => \N__41617\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__41626\,
            I => \N__41617\
        );

    \I__9434\ : Span4Mux_v
    port map (
            O => \N__41623\,
            I => \N__41614\
        );

    \I__9433\ : InMux
    port map (
            O => \N__41622\,
            I => \N__41611\
        );

    \I__9432\ : Span4Mux_h
    port map (
            O => \N__41617\,
            I => \N__41608\
        );

    \I__9431\ : Span4Mux_h
    port map (
            O => \N__41614\,
            I => \N__41605\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__41611\,
            I => measured_delay_hc_3
        );

    \I__9429\ : Odrv4
    port map (
            O => \N__41608\,
            I => measured_delay_hc_3
        );

    \I__9428\ : Odrv4
    port map (
            O => \N__41605\,
            I => measured_delay_hc_3
        );

    \I__9427\ : CascadeMux
    port map (
            O => \N__41598\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3_cascade_\
        );

    \I__9426\ : CascadeMux
    port map (
            O => \N__41595\,
            I => \N__41589\
        );

    \I__9425\ : CascadeMux
    port map (
            O => \N__41594\,
            I => \N__41586\
        );

    \I__9424\ : CascadeMux
    port map (
            O => \N__41593\,
            I => \N__41583\
        );

    \I__9423\ : CascadeMux
    port map (
            O => \N__41592\,
            I => \N__41579\
        );

    \I__9422\ : InMux
    port map (
            O => \N__41589\,
            I => \N__41576\
        );

    \I__9421\ : InMux
    port map (
            O => \N__41586\,
            I => \N__41573\
        );

    \I__9420\ : InMux
    port map (
            O => \N__41583\,
            I => \N__41570\
        );

    \I__9419\ : InMux
    port map (
            O => \N__41582\,
            I => \N__41567\
        );

    \I__9418\ : InMux
    port map (
            O => \N__41579\,
            I => \N__41564\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__41576\,
            I => \N__41557\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__41573\,
            I => \N__41557\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__41570\,
            I => \N__41557\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__41567\,
            I => \N__41554\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__41564\,
            I => \N__41549\
        );

    \I__9412\ : Span4Mux_v
    port map (
            O => \N__41557\,
            I => \N__41549\
        );

    \I__9411\ : Span4Mux_h
    port map (
            O => \N__41554\,
            I => \N__41546\
        );

    \I__9410\ : Odrv4
    port map (
            O => \N__41549\,
            I => measured_delay_hc_14
        );

    \I__9409\ : Odrv4
    port map (
            O => \N__41546\,
            I => measured_delay_hc_14
        );

    \I__9408\ : CascadeMux
    port map (
            O => \N__41541\,
            I => \N__41535\
        );

    \I__9407\ : CascadeMux
    port map (
            O => \N__41540\,
            I => \N__41532\
        );

    \I__9406\ : CascadeMux
    port map (
            O => \N__41539\,
            I => \N__41529\
        );

    \I__9405\ : CascadeMux
    port map (
            O => \N__41538\,
            I => \N__41526\
        );

    \I__9404\ : InMux
    port map (
            O => \N__41535\,
            I => \N__41518\
        );

    \I__9403\ : InMux
    port map (
            O => \N__41532\,
            I => \N__41501\
        );

    \I__9402\ : InMux
    port map (
            O => \N__41529\,
            I => \N__41501\
        );

    \I__9401\ : InMux
    port map (
            O => \N__41526\,
            I => \N__41501\
        );

    \I__9400\ : InMux
    port map (
            O => \N__41525\,
            I => \N__41501\
        );

    \I__9399\ : InMux
    port map (
            O => \N__41524\,
            I => \N__41501\
        );

    \I__9398\ : InMux
    port map (
            O => \N__41523\,
            I => \N__41501\
        );

    \I__9397\ : InMux
    port map (
            O => \N__41522\,
            I => \N__41501\
        );

    \I__9396\ : InMux
    port map (
            O => \N__41521\,
            I => \N__41501\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__41518\,
            I => \N__41489\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__41501\,
            I => \N__41486\
        );

    \I__9393\ : CascadeMux
    port map (
            O => \N__41500\,
            I => \N__41483\
        );

    \I__9392\ : CascadeMux
    port map (
            O => \N__41499\,
            I => \N__41480\
        );

    \I__9391\ : CascadeMux
    port map (
            O => \N__41498\,
            I => \N__41477\
        );

    \I__9390\ : CascadeMux
    port map (
            O => \N__41497\,
            I => \N__41472\
        );

    \I__9389\ : CascadeMux
    port map (
            O => \N__41496\,
            I => \N__41469\
        );

    \I__9388\ : CascadeMux
    port map (
            O => \N__41495\,
            I => \N__41466\
        );

    \I__9387\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41452\
        );

    \I__9386\ : InMux
    port map (
            O => \N__41493\,
            I => \N__41447\
        );

    \I__9385\ : InMux
    port map (
            O => \N__41492\,
            I => \N__41447\
        );

    \I__9384\ : Span4Mux_v
    port map (
            O => \N__41489\,
            I => \N__41442\
        );

    \I__9383\ : Span4Mux_h
    port map (
            O => \N__41486\,
            I => \N__41442\
        );

    \I__9382\ : InMux
    port map (
            O => \N__41483\,
            I => \N__41439\
        );

    \I__9381\ : InMux
    port map (
            O => \N__41480\,
            I => \N__41430\
        );

    \I__9380\ : InMux
    port map (
            O => \N__41477\,
            I => \N__41430\
        );

    \I__9379\ : InMux
    port map (
            O => \N__41476\,
            I => \N__41430\
        );

    \I__9378\ : InMux
    port map (
            O => \N__41475\,
            I => \N__41430\
        );

    \I__9377\ : InMux
    port map (
            O => \N__41472\,
            I => \N__41417\
        );

    \I__9376\ : InMux
    port map (
            O => \N__41469\,
            I => \N__41417\
        );

    \I__9375\ : InMux
    port map (
            O => \N__41466\,
            I => \N__41417\
        );

    \I__9374\ : InMux
    port map (
            O => \N__41465\,
            I => \N__41417\
        );

    \I__9373\ : InMux
    port map (
            O => \N__41464\,
            I => \N__41417\
        );

    \I__9372\ : InMux
    port map (
            O => \N__41463\,
            I => \N__41417\
        );

    \I__9371\ : InMux
    port map (
            O => \N__41462\,
            I => \N__41412\
        );

    \I__9370\ : InMux
    port map (
            O => \N__41461\,
            I => \N__41412\
        );

    \I__9369\ : InMux
    port map (
            O => \N__41460\,
            I => \N__41399\
        );

    \I__9368\ : InMux
    port map (
            O => \N__41459\,
            I => \N__41399\
        );

    \I__9367\ : InMux
    port map (
            O => \N__41458\,
            I => \N__41399\
        );

    \I__9366\ : InMux
    port map (
            O => \N__41457\,
            I => \N__41399\
        );

    \I__9365\ : InMux
    port map (
            O => \N__41456\,
            I => \N__41399\
        );

    \I__9364\ : InMux
    port map (
            O => \N__41455\,
            I => \N__41399\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__41452\,
            I => \N__41396\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__41447\,
            I => \N__41391\
        );

    \I__9361\ : Span4Mux_h
    port map (
            O => \N__41442\,
            I => \N__41391\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__41439\,
            I => \phase_controller_inst1.stoper_hc.N_405\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__41430\,
            I => \phase_controller_inst1.stoper_hc.N_405\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__41417\,
            I => \phase_controller_inst1.stoper_hc.N_405\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__41412\,
            I => \phase_controller_inst1.stoper_hc.N_405\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__41399\,
            I => \phase_controller_inst1.stoper_hc.N_405\
        );

    \I__9355\ : Odrv4
    port map (
            O => \N__41396\,
            I => \phase_controller_inst1.stoper_hc.N_405\
        );

    \I__9354\ : Odrv4
    port map (
            O => \N__41391\,
            I => \phase_controller_inst1.stoper_hc.N_405\
        );

    \I__9353\ : CascadeMux
    port map (
            O => \N__41376\,
            I => \N__41370\
        );

    \I__9352\ : InMux
    port map (
            O => \N__41375\,
            I => \N__41367\
        );

    \I__9351\ : InMux
    port map (
            O => \N__41374\,
            I => \N__41364\
        );

    \I__9350\ : InMux
    port map (
            O => \N__41373\,
            I => \N__41361\
        );

    \I__9349\ : InMux
    port map (
            O => \N__41370\,
            I => \N__41357\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__41367\,
            I => \N__41354\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__41364\,
            I => \N__41349\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__41361\,
            I => \N__41349\
        );

    \I__9345\ : InMux
    port map (
            O => \N__41360\,
            I => \N__41346\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__41357\,
            I => \N__41343\
        );

    \I__9343\ : Span4Mux_h
    port map (
            O => \N__41354\,
            I => \N__41340\
        );

    \I__9342\ : Span12Mux_s11_h
    port map (
            O => \N__41349\,
            I => \N__41337\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__41346\,
            I => measured_delay_hc_9
        );

    \I__9340\ : Odrv4
    port map (
            O => \N__41343\,
            I => measured_delay_hc_9
        );

    \I__9339\ : Odrv4
    port map (
            O => \N__41340\,
            I => measured_delay_hc_9
        );

    \I__9338\ : Odrv12
    port map (
            O => \N__41337\,
            I => measured_delay_hc_9
        );

    \I__9337\ : CascadeMux
    port map (
            O => \N__41328\,
            I => \N__41325\
        );

    \I__9336\ : InMux
    port map (
            O => \N__41325\,
            I => \N__41322\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__41322\,
            I => \N__41318\
        );

    \I__9334\ : InMux
    port map (
            O => \N__41321\,
            I => \N__41315\
        );

    \I__9333\ : Span4Mux_h
    port map (
            O => \N__41318\,
            I => \N__41312\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__41315\,
            I => \N__41307\
        );

    \I__9331\ : Span4Mux_v
    port map (
            O => \N__41312\,
            I => \N__41307\
        );

    \I__9330\ : Odrv4
    port map (
            O => \N__41307\,
            I => measured_delay_hc_30
        );

    \I__9329\ : InMux
    port map (
            O => \N__41304\,
            I => \N__41301\
        );

    \I__9328\ : LocalMux
    port map (
            O => \N__41301\,
            I => \N__41298\
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__41298\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6Z0Z_19\
        );

    \I__9326\ : CascadeMux
    port map (
            O => \N__41295\,
            I => \N__41289\
        );

    \I__9325\ : InMux
    port map (
            O => \N__41294\,
            I => \N__41286\
        );

    \I__9324\ : InMux
    port map (
            O => \N__41293\,
            I => \N__41283\
        );

    \I__9323\ : CascadeMux
    port map (
            O => \N__41292\,
            I => \N__41279\
        );

    \I__9322\ : InMux
    port map (
            O => \N__41289\,
            I => \N__41276\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__41286\,
            I => \N__41271\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__41283\,
            I => \N__41271\
        );

    \I__9319\ : InMux
    port map (
            O => \N__41282\,
            I => \N__41268\
        );

    \I__9318\ : InMux
    port map (
            O => \N__41279\,
            I => \N__41265\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__41276\,
            I => \N__41258\
        );

    \I__9316\ : Span4Mux_v
    port map (
            O => \N__41271\,
            I => \N__41258\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__41268\,
            I => \N__41258\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__41265\,
            I => measured_delay_hc_6
        );

    \I__9313\ : Odrv4
    port map (
            O => \N__41258\,
            I => measured_delay_hc_6
        );

    \I__9312\ : InMux
    port map (
            O => \N__41253\,
            I => \N__41249\
        );

    \I__9311\ : InMux
    port map (
            O => \N__41252\,
            I => \N__41246\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__41249\,
            I => measured_delay_hc_29
        );

    \I__9309\ : LocalMux
    port map (
            O => \N__41246\,
            I => measured_delay_hc_29
        );

    \I__9308\ : InMux
    port map (
            O => \N__41241\,
            I => \N__41235\
        );

    \I__9307\ : InMux
    port map (
            O => \N__41240\,
            I => \N__41232\
        );

    \I__9306\ : InMux
    port map (
            O => \N__41239\,
            I => \N__41229\
        );

    \I__9305\ : CascadeMux
    port map (
            O => \N__41238\,
            I => \N__41226\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__41235\,
            I => \N__41219\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__41232\,
            I => \N__41219\
        );

    \I__9302\ : LocalMux
    port map (
            O => \N__41229\,
            I => \N__41216\
        );

    \I__9301\ : InMux
    port map (
            O => \N__41226\,
            I => \N__41213\
        );

    \I__9300\ : InMux
    port map (
            O => \N__41225\,
            I => \N__41208\
        );

    \I__9299\ : InMux
    port map (
            O => \N__41224\,
            I => \N__41208\
        );

    \I__9298\ : Span4Mux_v
    port map (
            O => \N__41219\,
            I => \N__41203\
        );

    \I__9297\ : Span4Mux_v
    port map (
            O => \N__41216\,
            I => \N__41203\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__41213\,
            I => measured_delay_hc_7
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__41208\,
            I => measured_delay_hc_7
        );

    \I__9294\ : Odrv4
    port map (
            O => \N__41203\,
            I => measured_delay_hc_7
        );

    \I__9293\ : InMux
    port map (
            O => \N__41196\,
            I => \N__41192\
        );

    \I__9292\ : InMux
    port map (
            O => \N__41195\,
            I => \N__41188\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__41192\,
            I => \N__41183\
        );

    \I__9290\ : InMux
    port map (
            O => \N__41191\,
            I => \N__41180\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__41188\,
            I => \N__41177\
        );

    \I__9288\ : CascadeMux
    port map (
            O => \N__41187\,
            I => \N__41174\
        );

    \I__9287\ : InMux
    port map (
            O => \N__41186\,
            I => \N__41171\
        );

    \I__9286\ : Span4Mux_h
    port map (
            O => \N__41183\,
            I => \N__41168\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__41180\,
            I => \N__41163\
        );

    \I__9284\ : Span4Mux_v
    port map (
            O => \N__41177\,
            I => \N__41163\
        );

    \I__9283\ : InMux
    port map (
            O => \N__41174\,
            I => \N__41160\
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__41171\,
            I => measured_delay_hc_5
        );

    \I__9281\ : Odrv4
    port map (
            O => \N__41168\,
            I => measured_delay_hc_5
        );

    \I__9280\ : Odrv4
    port map (
            O => \N__41163\,
            I => measured_delay_hc_5
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__41160\,
            I => measured_delay_hc_5
        );

    \I__9278\ : InMux
    port map (
            O => \N__41151\,
            I => \N__41148\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__41148\,
            I => \N__41145\
        );

    \I__9276\ : Odrv4
    port map (
            O => \N__41145\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3Z0Z_18\
        );

    \I__9275\ : CascadeMux
    port map (
            O => \N__41142\,
            I => \N__41139\
        );

    \I__9274\ : InMux
    port map (
            O => \N__41139\,
            I => \N__41136\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__41136\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3Z0Z_2\
        );

    \I__9272\ : InMux
    port map (
            O => \N__41133\,
            I => \N__41130\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__41130\,
            I => \phase_controller_inst1.stoper_hc.N_388\
        );

    \I__9270\ : CascadeMux
    port map (
            O => \N__41127\,
            I => \phase_controller_inst1.stoper_hc.N_405_cascade_\
        );

    \I__9269\ : InMux
    port map (
            O => \N__41124\,
            I => \N__41120\
        );

    \I__9268\ : InMux
    port map (
            O => \N__41123\,
            I => \N__41115\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__41120\,
            I => \N__41112\
        );

    \I__9266\ : InMux
    port map (
            O => \N__41119\,
            I => \N__41109\
        );

    \I__9265\ : InMux
    port map (
            O => \N__41118\,
            I => \N__41106\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__41115\,
            I => \N__41103\
        );

    \I__9263\ : Span4Mux_h
    port map (
            O => \N__41112\,
            I => \N__41098\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__41109\,
            I => \N__41098\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__41106\,
            I => \N__41092\
        );

    \I__9260\ : Span4Mux_v
    port map (
            O => \N__41103\,
            I => \N__41092\
        );

    \I__9259\ : Span4Mux_v
    port map (
            O => \N__41098\,
            I => \N__41089\
        );

    \I__9258\ : InMux
    port map (
            O => \N__41097\,
            I => \N__41086\
        );

    \I__9257\ : Odrv4
    port map (
            O => \N__41092\,
            I => measured_delay_hc_4
        );

    \I__9256\ : Odrv4
    port map (
            O => \N__41089\,
            I => measured_delay_hc_4
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__41086\,
            I => measured_delay_hc_4
        );

    \I__9254\ : CascadeMux
    port map (
            O => \N__41079\,
            I => \N__41076\
        );

    \I__9253\ : InMux
    port map (
            O => \N__41076\,
            I => \N__41072\
        );

    \I__9252\ : CascadeMux
    port map (
            O => \N__41075\,
            I => \N__41066\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__41072\,
            I => \N__41063\
        );

    \I__9250\ : InMux
    port map (
            O => \N__41071\,
            I => \N__41060\
        );

    \I__9249\ : InMux
    port map (
            O => \N__41070\,
            I => \N__41057\
        );

    \I__9248\ : InMux
    port map (
            O => \N__41069\,
            I => \N__41054\
        );

    \I__9247\ : InMux
    port map (
            O => \N__41066\,
            I => \N__41051\
        );

    \I__9246\ : Span4Mux_v
    port map (
            O => \N__41063\,
            I => \N__41046\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__41060\,
            I => \N__41046\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__41057\,
            I => \N__41041\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__41054\,
            I => \N__41041\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__41051\,
            I => measured_delay_hc_10
        );

    \I__9241\ : Odrv4
    port map (
            O => \N__41046\,
            I => measured_delay_hc_10
        );

    \I__9240\ : Odrv4
    port map (
            O => \N__41041\,
            I => measured_delay_hc_10
        );

    \I__9239\ : InMux
    port map (
            O => \N__41034\,
            I => \N__41031\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__41031\,
            I => \N__41025\
        );

    \I__9237\ : CascadeMux
    port map (
            O => \N__41030\,
            I => \N__41022\
        );

    \I__9236\ : CascadeMux
    port map (
            O => \N__41029\,
            I => \N__41019\
        );

    \I__9235\ : InMux
    port map (
            O => \N__41028\,
            I => \N__41015\
        );

    \I__9234\ : Span4Mux_h
    port map (
            O => \N__41025\,
            I => \N__41012\
        );

    \I__9233\ : InMux
    port map (
            O => \N__41022\,
            I => \N__41009\
        );

    \I__9232\ : InMux
    port map (
            O => \N__41019\,
            I => \N__41004\
        );

    \I__9231\ : InMux
    port map (
            O => \N__41018\,
            I => \N__41004\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__41015\,
            I => \N__41001\
        );

    \I__9229\ : Odrv4
    port map (
            O => \N__41012\,
            I => measured_delay_hc_11
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__41009\,
            I => measured_delay_hc_11
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__41004\,
            I => measured_delay_hc_11
        );

    \I__9226\ : Odrv4
    port map (
            O => \N__41001\,
            I => measured_delay_hc_11
        );

    \I__9225\ : CascadeMux
    port map (
            O => \N__40992\,
            I => \N__40987\
        );

    \I__9224\ : InMux
    port map (
            O => \N__40991\,
            I => \N__40984\
        );

    \I__9223\ : CascadeMux
    port map (
            O => \N__40990\,
            I => \N__40981\
        );

    \I__9222\ : InMux
    port map (
            O => \N__40987\,
            I => \N__40978\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__40984\,
            I => \N__40975\
        );

    \I__9220\ : InMux
    port map (
            O => \N__40981\,
            I => \N__40972\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__40978\,
            I => \N__40967\
        );

    \I__9218\ : Span4Mux_h
    port map (
            O => \N__40975\,
            I => \N__40962\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__40972\,
            I => \N__40962\
        );

    \I__9216\ : InMux
    port map (
            O => \N__40971\,
            I => \N__40957\
        );

    \I__9215\ : InMux
    port map (
            O => \N__40970\,
            I => \N__40957\
        );

    \I__9214\ : Odrv4
    port map (
            O => \N__40967\,
            I => measured_delay_hc_12
        );

    \I__9213\ : Odrv4
    port map (
            O => \N__40962\,
            I => measured_delay_hc_12
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__40957\,
            I => measured_delay_hc_12
        );

    \I__9211\ : InMux
    port map (
            O => \N__40950\,
            I => \N__40947\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__40947\,
            I => \N__40942\
        );

    \I__9209\ : InMux
    port map (
            O => \N__40946\,
            I => \N__40939\
        );

    \I__9208\ : InMux
    port map (
            O => \N__40945\,
            I => \N__40934\
        );

    \I__9207\ : Span4Mux_h
    port map (
            O => \N__40942\,
            I => \N__40929\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__40939\,
            I => \N__40929\
        );

    \I__9205\ : InMux
    port map (
            O => \N__40938\,
            I => \N__40926\
        );

    \I__9204\ : CascadeMux
    port map (
            O => \N__40937\,
            I => \N__40923\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__40934\,
            I => \N__40918\
        );

    \I__9202\ : Span4Mux_h
    port map (
            O => \N__40929\,
            I => \N__40918\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__40926\,
            I => \N__40915\
        );

    \I__9200\ : InMux
    port map (
            O => \N__40923\,
            I => \N__40912\
        );

    \I__9199\ : Span4Mux_v
    port map (
            O => \N__40918\,
            I => \N__40907\
        );

    \I__9198\ : Span4Mux_h
    port map (
            O => \N__40915\,
            I => \N__40907\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__40912\,
            I => measured_delay_hc_8
        );

    \I__9196\ : Odrv4
    port map (
            O => \N__40907\,
            I => measured_delay_hc_8
        );

    \I__9195\ : InMux
    port map (
            O => \N__40902\,
            I => \N__40899\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__40899\,
            I => \N__40895\
        );

    \I__9193\ : InMux
    port map (
            O => \N__40898\,
            I => \N__40892\
        );

    \I__9192\ : Span4Mux_h
    port map (
            O => \N__40895\,
            I => \N__40889\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__40892\,
            I => \N__40886\
        );

    \I__9190\ : Odrv4
    port map (
            O => \N__40889\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_1\
        );

    \I__9189\ : Odrv4
    port map (
            O => \N__40886\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_1\
        );

    \I__9188\ : CascadeMux
    port map (
            O => \N__40881\,
            I => \N__40878\
        );

    \I__9187\ : InMux
    port map (
            O => \N__40878\,
            I => \N__40875\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__40875\,
            I => \N__40872\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__40872\,
            I => \N__40869\
        );

    \I__9184\ : Odrv4
    port map (
            O => \N__40869\,
            I => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__9183\ : InMux
    port map (
            O => \N__40866\,
            I => \N__40862\
        );

    \I__9182\ : InMux
    port map (
            O => \N__40865\,
            I => \N__40859\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__40862\,
            I => \N__40855\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__40859\,
            I => \N__40852\
        );

    \I__9179\ : InMux
    port map (
            O => \N__40858\,
            I => \N__40849\
        );

    \I__9178\ : Odrv4
    port map (
            O => \N__40855\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__9177\ : Odrv4
    port map (
            O => \N__40852\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__40849\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__9175\ : InMux
    port map (
            O => \N__40842\,
            I => \N__40839\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__40839\,
            I => \N__40834\
        );

    \I__9173\ : InMux
    port map (
            O => \N__40838\,
            I => \N__40831\
        );

    \I__9172\ : InMux
    port map (
            O => \N__40837\,
            I => \N__40828\
        );

    \I__9171\ : Span4Mux_h
    port map (
            O => \N__40834\,
            I => \N__40825\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__40831\,
            I => \N__40822\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__40828\,
            I => \N__40819\
        );

    \I__9168\ : Sp12to4
    port map (
            O => \N__40825\,
            I => \N__40816\
        );

    \I__9167\ : Sp12to4
    port map (
            O => \N__40822\,
            I => \N__40813\
        );

    \I__9166\ : Span4Mux_h
    port map (
            O => \N__40819\,
            I => \N__40810\
        );

    \I__9165\ : Span12Mux_v
    port map (
            O => \N__40816\,
            I => \N__40807\
        );

    \I__9164\ : Span12Mux_s10_v
    port map (
            O => \N__40813\,
            I => \N__40804\
        );

    \I__9163\ : Odrv4
    port map (
            O => \N__40810\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__9162\ : Odrv12
    port map (
            O => \N__40807\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__9161\ : Odrv12
    port map (
            O => \N__40804\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__9160\ : CascadeMux
    port map (
            O => \N__40797\,
            I => \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa_cascade_\
        );

    \I__9159\ : InMux
    port map (
            O => \N__40794\,
            I => \N__40789\
        );

    \I__9158\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40786\
        );

    \I__9157\ : InMux
    port map (
            O => \N__40792\,
            I => \N__40783\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__40789\,
            I => \N__40777\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__40786\,
            I => \N__40777\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__40783\,
            I => \N__40774\
        );

    \I__9153\ : InMux
    port map (
            O => \N__40782\,
            I => \N__40771\
        );

    \I__9152\ : Span12Mux_h
    port map (
            O => \N__40777\,
            I => \N__40768\
        );

    \I__9151\ : Odrv12
    port map (
            O => \N__40774\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__40771\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__9149\ : Odrv12
    port map (
            O => \N__40768\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__9148\ : InMux
    port map (
            O => \N__40761\,
            I => \N__40756\
        );

    \I__9147\ : InMux
    port map (
            O => \N__40760\,
            I => \N__40753\
        );

    \I__9146\ : InMux
    port map (
            O => \N__40759\,
            I => \N__40750\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__40756\,
            I => \N__40744\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__40753\,
            I => \N__40744\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__40750\,
            I => \N__40741\
        );

    \I__9142\ : InMux
    port map (
            O => \N__40749\,
            I => \N__40738\
        );

    \I__9141\ : Span4Mux_v
    port map (
            O => \N__40744\,
            I => \N__40733\
        );

    \I__9140\ : Span4Mux_h
    port map (
            O => \N__40741\,
            I => \N__40733\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__40738\,
            I => \N__40730\
        );

    \I__9138\ : Span4Mux_v
    port map (
            O => \N__40733\,
            I => \N__40727\
        );

    \I__9137\ : Span4Mux_v
    port map (
            O => \N__40730\,
            I => \N__40724\
        );

    \I__9136\ : Odrv4
    port map (
            O => \N__40727\,
            I => delay_hc_d2
        );

    \I__9135\ : Odrv4
    port map (
            O => \N__40724\,
            I => delay_hc_d2
        );

    \I__9134\ : InMux
    port map (
            O => \N__40719\,
            I => \N__40716\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__40716\,
            I => \N__40712\
        );

    \I__9132\ : InMux
    port map (
            O => \N__40715\,
            I => \N__40709\
        );

    \I__9131\ : Span12Mux_h
    port map (
            O => \N__40712\,
            I => \N__40705\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__40709\,
            I => \N__40702\
        );

    \I__9129\ : InMux
    port map (
            O => \N__40708\,
            I => \N__40699\
        );

    \I__9128\ : Odrv12
    port map (
            O => \N__40705\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__9127\ : Odrv4
    port map (
            O => \N__40702\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__40699\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__9125\ : CascadeMux
    port map (
            O => \N__40692\,
            I => \N__40688\
        );

    \I__9124\ : CascadeMux
    port map (
            O => \N__40691\,
            I => \N__40685\
        );

    \I__9123\ : InMux
    port map (
            O => \N__40688\,
            I => \N__40679\
        );

    \I__9122\ : InMux
    port map (
            O => \N__40685\,
            I => \N__40679\
        );

    \I__9121\ : InMux
    port map (
            O => \N__40684\,
            I => \N__40676\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__40679\,
            I => \N__40673\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__40676\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__9118\ : Odrv4
    port map (
            O => \N__40673\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__9117\ : InMux
    port map (
            O => \N__40668\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__9116\ : InMux
    port map (
            O => \N__40665\,
            I => \N__40661\
        );

    \I__9115\ : CascadeMux
    port map (
            O => \N__40664\,
            I => \N__40658\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__40661\,
            I => \N__40654\
        );

    \I__9113\ : InMux
    port map (
            O => \N__40658\,
            I => \N__40651\
        );

    \I__9112\ : InMux
    port map (
            O => \N__40657\,
            I => \N__40648\
        );

    \I__9111\ : Span4Mux_v
    port map (
            O => \N__40654\,
            I => \N__40643\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__40651\,
            I => \N__40643\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__40648\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__9108\ : Odrv4
    port map (
            O => \N__40643\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__9107\ : InMux
    port map (
            O => \N__40638\,
            I => \bfn_17_11_0_\
        );

    \I__9106\ : CascadeMux
    port map (
            O => \N__40635\,
            I => \N__40632\
        );

    \I__9105\ : InMux
    port map (
            O => \N__40632\,
            I => \N__40629\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__40629\,
            I => \N__40624\
        );

    \I__9103\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40621\
        );

    \I__9102\ : InMux
    port map (
            O => \N__40627\,
            I => \N__40618\
        );

    \I__9101\ : Span4Mux_v
    port map (
            O => \N__40624\,
            I => \N__40615\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__40621\,
            I => \N__40612\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__40618\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__9098\ : Odrv4
    port map (
            O => \N__40615\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__9097\ : Odrv4
    port map (
            O => \N__40612\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__9096\ : InMux
    port map (
            O => \N__40605\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__9095\ : CascadeMux
    port map (
            O => \N__40602\,
            I => \N__40598\
        );

    \I__9094\ : CascadeMux
    port map (
            O => \N__40601\,
            I => \N__40595\
        );

    \I__9093\ : InMux
    port map (
            O => \N__40598\,
            I => \N__40589\
        );

    \I__9092\ : InMux
    port map (
            O => \N__40595\,
            I => \N__40589\
        );

    \I__9091\ : InMux
    port map (
            O => \N__40594\,
            I => \N__40586\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__40589\,
            I => \N__40583\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__40586\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__9088\ : Odrv4
    port map (
            O => \N__40583\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__9087\ : InMux
    port map (
            O => \N__40578\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__9086\ : InMux
    port map (
            O => \N__40575\,
            I => \N__40568\
        );

    \I__9085\ : InMux
    port map (
            O => \N__40574\,
            I => \N__40568\
        );

    \I__9084\ : InMux
    port map (
            O => \N__40573\,
            I => \N__40565\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__40568\,
            I => \N__40562\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__40565\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__9081\ : Odrv4
    port map (
            O => \N__40562\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__9080\ : InMux
    port map (
            O => \N__40557\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__9079\ : InMux
    port map (
            O => \N__40554\,
            I => \N__40551\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__40551\,
            I => \N__40547\
        );

    \I__9077\ : InMux
    port map (
            O => \N__40550\,
            I => \N__40544\
        );

    \I__9076\ : Span4Mux_h
    port map (
            O => \N__40547\,
            I => \N__40541\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__40544\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__9074\ : Odrv4
    port map (
            O => \N__40541\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__9073\ : InMux
    port map (
            O => \N__40536\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__9072\ : InMux
    port map (
            O => \N__40533\,
            I => \N__40513\
        );

    \I__9071\ : InMux
    port map (
            O => \N__40532\,
            I => \N__40513\
        );

    \I__9070\ : InMux
    port map (
            O => \N__40531\,
            I => \N__40513\
        );

    \I__9069\ : InMux
    port map (
            O => \N__40530\,
            I => \N__40513\
        );

    \I__9068\ : InMux
    port map (
            O => \N__40529\,
            I => \N__40504\
        );

    \I__9067\ : InMux
    port map (
            O => \N__40528\,
            I => \N__40504\
        );

    \I__9066\ : InMux
    port map (
            O => \N__40527\,
            I => \N__40504\
        );

    \I__9065\ : InMux
    port map (
            O => \N__40526\,
            I => \N__40504\
        );

    \I__9064\ : InMux
    port map (
            O => \N__40525\,
            I => \N__40495\
        );

    \I__9063\ : InMux
    port map (
            O => \N__40524\,
            I => \N__40495\
        );

    \I__9062\ : InMux
    port map (
            O => \N__40523\,
            I => \N__40495\
        );

    \I__9061\ : InMux
    port map (
            O => \N__40522\,
            I => \N__40495\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__40513\,
            I => \N__40478\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__40504\,
            I => \N__40478\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__40495\,
            I => \N__40478\
        );

    \I__9057\ : InMux
    port map (
            O => \N__40494\,
            I => \N__40473\
        );

    \I__9056\ : InMux
    port map (
            O => \N__40493\,
            I => \N__40473\
        );

    \I__9055\ : InMux
    port map (
            O => \N__40492\,
            I => \N__40464\
        );

    \I__9054\ : InMux
    port map (
            O => \N__40491\,
            I => \N__40464\
        );

    \I__9053\ : InMux
    port map (
            O => \N__40490\,
            I => \N__40464\
        );

    \I__9052\ : InMux
    port map (
            O => \N__40489\,
            I => \N__40464\
        );

    \I__9051\ : InMux
    port map (
            O => \N__40488\,
            I => \N__40447\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40487\,
            I => \N__40447\
        );

    \I__9049\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40447\
        );

    \I__9048\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40447\
        );

    \I__9047\ : Span4Mux_v
    port map (
            O => \N__40478\,
            I => \N__40440\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__40473\,
            I => \N__40440\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__40464\,
            I => \N__40440\
        );

    \I__9044\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40431\
        );

    \I__9043\ : InMux
    port map (
            O => \N__40462\,
            I => \N__40431\
        );

    \I__9042\ : InMux
    port map (
            O => \N__40461\,
            I => \N__40431\
        );

    \I__9041\ : InMux
    port map (
            O => \N__40460\,
            I => \N__40431\
        );

    \I__9040\ : InMux
    port map (
            O => \N__40459\,
            I => \N__40422\
        );

    \I__9039\ : InMux
    port map (
            O => \N__40458\,
            I => \N__40422\
        );

    \I__9038\ : InMux
    port map (
            O => \N__40457\,
            I => \N__40422\
        );

    \I__9037\ : InMux
    port map (
            O => \N__40456\,
            I => \N__40422\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__40447\,
            I => \N__40417\
        );

    \I__9035\ : Span4Mux_v
    port map (
            O => \N__40440\,
            I => \N__40417\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__40431\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__40422\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9032\ : Odrv4
    port map (
            O => \N__40417\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9031\ : InMux
    port map (
            O => \N__40410\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__9030\ : CascadeMux
    port map (
            O => \N__40407\,
            I => \N__40404\
        );

    \I__9029\ : InMux
    port map (
            O => \N__40404\,
            I => \N__40401\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__40401\,
            I => \N__40397\
        );

    \I__9027\ : InMux
    port map (
            O => \N__40400\,
            I => \N__40394\
        );

    \I__9026\ : Span4Mux_h
    port map (
            O => \N__40397\,
            I => \N__40391\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__40394\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__9024\ : Odrv4
    port map (
            O => \N__40391\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__9023\ : CEMux
    port map (
            O => \N__40386\,
            I => \N__40382\
        );

    \I__9022\ : CEMux
    port map (
            O => \N__40385\,
            I => \N__40379\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__40382\,
            I => \N__40372\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__40379\,
            I => \N__40372\
        );

    \I__9019\ : CEMux
    port map (
            O => \N__40378\,
            I => \N__40369\
        );

    \I__9018\ : CEMux
    port map (
            O => \N__40377\,
            I => \N__40366\
        );

    \I__9017\ : Span4Mux_v
    port map (
            O => \N__40372\,
            I => \N__40363\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__40369\,
            I => \N__40358\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__40366\,
            I => \N__40358\
        );

    \I__9014\ : Span4Mux_h
    port map (
            O => \N__40363\,
            I => \N__40353\
        );

    \I__9013\ : Span4Mux_v
    port map (
            O => \N__40358\,
            I => \N__40353\
        );

    \I__9012\ : Span4Mux_h
    port map (
            O => \N__40353\,
            I => \N__40350\
        );

    \I__9011\ : Odrv4
    port map (
            O => \N__40350\,
            I => \delay_measurement_inst.delay_tr_timer.N_464_i\
        );

    \I__9010\ : InMux
    port map (
            O => \N__40347\,
            I => \N__40344\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__40344\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9008\ : InMux
    port map (
            O => \N__40341\,
            I => \N__40338\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__40338\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9006\ : InMux
    port map (
            O => \N__40335\,
            I => \N__40332\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__40332\,
            I => \N__40329\
        );

    \I__9004\ : Odrv4
    port map (
            O => \N__40329\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\
        );

    \I__9003\ : CascadeMux
    port map (
            O => \N__40326\,
            I => \N__40322\
        );

    \I__9002\ : CascadeMux
    port map (
            O => \N__40325\,
            I => \N__40319\
        );

    \I__9001\ : InMux
    port map (
            O => \N__40322\,
            I => \N__40314\
        );

    \I__9000\ : InMux
    port map (
            O => \N__40319\,
            I => \N__40314\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__40314\,
            I => \N__40310\
        );

    \I__8998\ : InMux
    port map (
            O => \N__40313\,
            I => \N__40307\
        );

    \I__8997\ : Span4Mux_h
    port map (
            O => \N__40310\,
            I => \N__40304\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__40307\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8995\ : Odrv4
    port map (
            O => \N__40304\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8994\ : InMux
    port map (
            O => \N__40299\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__8993\ : CascadeMux
    port map (
            O => \N__40296\,
            I => \N__40292\
        );

    \I__8992\ : CascadeMux
    port map (
            O => \N__40295\,
            I => \N__40289\
        );

    \I__8991\ : InMux
    port map (
            O => \N__40292\,
            I => \N__40283\
        );

    \I__8990\ : InMux
    port map (
            O => \N__40289\,
            I => \N__40283\
        );

    \I__8989\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40280\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__40283\,
            I => \N__40277\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__40280\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8986\ : Odrv4
    port map (
            O => \N__40277\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8985\ : InMux
    port map (
            O => \N__40272\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__8984\ : InMux
    port map (
            O => \N__40269\,
            I => \N__40265\
        );

    \I__8983\ : InMux
    port map (
            O => \N__40268\,
            I => \N__40262\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__40265\,
            I => \N__40259\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__40262\,
            I => \N__40255\
        );

    \I__8980\ : Span4Mux_v
    port map (
            O => \N__40259\,
            I => \N__40252\
        );

    \I__8979\ : InMux
    port map (
            O => \N__40258\,
            I => \N__40249\
        );

    \I__8978\ : Span4Mux_h
    port map (
            O => \N__40255\,
            I => \N__40246\
        );

    \I__8977\ : Odrv4
    port map (
            O => \N__40252\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__40249\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8975\ : Odrv4
    port map (
            O => \N__40246\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8974\ : InMux
    port map (
            O => \N__40239\,
            I => \bfn_17_10_0_\
        );

    \I__8973\ : InMux
    port map (
            O => \N__40236\,
            I => \N__40233\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__40233\,
            I => \N__40228\
        );

    \I__8971\ : InMux
    port map (
            O => \N__40232\,
            I => \N__40225\
        );

    \I__8970\ : InMux
    port map (
            O => \N__40231\,
            I => \N__40222\
        );

    \I__8969\ : Span4Mux_v
    port map (
            O => \N__40228\,
            I => \N__40217\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__40225\,
            I => \N__40217\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__40222\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8966\ : Odrv4
    port map (
            O => \N__40217\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8965\ : InMux
    port map (
            O => \N__40212\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__8964\ : CascadeMux
    port map (
            O => \N__40209\,
            I => \N__40205\
        );

    \I__8963\ : CascadeMux
    port map (
            O => \N__40208\,
            I => \N__40202\
        );

    \I__8962\ : InMux
    port map (
            O => \N__40205\,
            I => \N__40196\
        );

    \I__8961\ : InMux
    port map (
            O => \N__40202\,
            I => \N__40196\
        );

    \I__8960\ : InMux
    port map (
            O => \N__40201\,
            I => \N__40193\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__40196\,
            I => \N__40190\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__40193\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__8957\ : Odrv4
    port map (
            O => \N__40190\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__8956\ : InMux
    port map (
            O => \N__40185\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__8955\ : CascadeMux
    port map (
            O => \N__40182\,
            I => \N__40178\
        );

    \I__8954\ : CascadeMux
    port map (
            O => \N__40181\,
            I => \N__40175\
        );

    \I__8953\ : InMux
    port map (
            O => \N__40178\,
            I => \N__40170\
        );

    \I__8952\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40170\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__40170\,
            I => \N__40166\
        );

    \I__8950\ : InMux
    port map (
            O => \N__40169\,
            I => \N__40163\
        );

    \I__8949\ : Span4Mux_h
    port map (
            O => \N__40166\,
            I => \N__40160\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__40163\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8947\ : Odrv4
    port map (
            O => \N__40160\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8946\ : InMux
    port map (
            O => \N__40155\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__8945\ : CascadeMux
    port map (
            O => \N__40152\,
            I => \N__40148\
        );

    \I__8944\ : InMux
    port map (
            O => \N__40151\,
            I => \N__40145\
        );

    \I__8943\ : InMux
    port map (
            O => \N__40148\,
            I => \N__40141\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__40145\,
            I => \N__40138\
        );

    \I__8941\ : InMux
    port map (
            O => \N__40144\,
            I => \N__40135\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__40141\,
            I => \N__40130\
        );

    \I__8939\ : Span4Mux_h
    port map (
            O => \N__40138\,
            I => \N__40130\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__40135\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__8937\ : Odrv4
    port map (
            O => \N__40130\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__8936\ : InMux
    port map (
            O => \N__40125\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__8935\ : InMux
    port map (
            O => \N__40122\,
            I => \N__40115\
        );

    \I__8934\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40115\
        );

    \I__8933\ : InMux
    port map (
            O => \N__40120\,
            I => \N__40112\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__40115\,
            I => \N__40109\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__40112\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8930\ : Odrv4
    port map (
            O => \N__40109\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8929\ : InMux
    port map (
            O => \N__40104\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__8928\ : InMux
    port map (
            O => \N__40101\,
            I => \N__40094\
        );

    \I__8927\ : InMux
    port map (
            O => \N__40100\,
            I => \N__40094\
        );

    \I__8926\ : InMux
    port map (
            O => \N__40099\,
            I => \N__40091\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__40094\,
            I => \N__40088\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__40091\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8923\ : Odrv4
    port map (
            O => \N__40088\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8922\ : InMux
    port map (
            O => \N__40083\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__8921\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40073\
        );

    \I__8920\ : InMux
    port map (
            O => \N__40079\,
            I => \N__40073\
        );

    \I__8919\ : InMux
    port map (
            O => \N__40078\,
            I => \N__40070\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__40073\,
            I => \N__40067\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__40070\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8916\ : Odrv4
    port map (
            O => \N__40067\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8915\ : InMux
    port map (
            O => \N__40062\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__8914\ : CascadeMux
    port map (
            O => \N__40059\,
            I => \N__40055\
        );

    \I__8913\ : CascadeMux
    port map (
            O => \N__40058\,
            I => \N__40052\
        );

    \I__8912\ : InMux
    port map (
            O => \N__40055\,
            I => \N__40047\
        );

    \I__8911\ : InMux
    port map (
            O => \N__40052\,
            I => \N__40047\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__40047\,
            I => \N__40043\
        );

    \I__8909\ : InMux
    port map (
            O => \N__40046\,
            I => \N__40040\
        );

    \I__8908\ : Span4Mux_h
    port map (
            O => \N__40043\,
            I => \N__40037\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__40040\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8906\ : Odrv4
    port map (
            O => \N__40037\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8905\ : InMux
    port map (
            O => \N__40032\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__8904\ : InMux
    port map (
            O => \N__40029\,
            I => \N__40025\
        );

    \I__8903\ : CascadeMux
    port map (
            O => \N__40028\,
            I => \N__40022\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__40025\,
            I => \N__40018\
        );

    \I__8901\ : InMux
    port map (
            O => \N__40022\,
            I => \N__40015\
        );

    \I__8900\ : InMux
    port map (
            O => \N__40021\,
            I => \N__40012\
        );

    \I__8899\ : Span4Mux_v
    port map (
            O => \N__40018\,
            I => \N__40007\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__40015\,
            I => \N__40007\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__40012\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8896\ : Odrv4
    port map (
            O => \N__40007\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8895\ : InMux
    port map (
            O => \N__40002\,
            I => \bfn_17_9_0_\
        );

    \I__8894\ : CascadeMux
    port map (
            O => \N__39999\,
            I => \N__39996\
        );

    \I__8893\ : InMux
    port map (
            O => \N__39996\,
            I => \N__39992\
        );

    \I__8892\ : InMux
    port map (
            O => \N__39995\,
            I => \N__39988\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__39992\,
            I => \N__39985\
        );

    \I__8890\ : InMux
    port map (
            O => \N__39991\,
            I => \N__39982\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__39988\,
            I => \N__39977\
        );

    \I__8888\ : Span4Mux_v
    port map (
            O => \N__39985\,
            I => \N__39977\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__39982\,
            I => \N__39974\
        );

    \I__8886\ : Odrv4
    port map (
            O => \N__39977\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8885\ : Odrv4
    port map (
            O => \N__39974\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8884\ : InMux
    port map (
            O => \N__39969\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__8883\ : CascadeMux
    port map (
            O => \N__39966\,
            I => \N__39962\
        );

    \I__8882\ : CascadeMux
    port map (
            O => \N__39965\,
            I => \N__39959\
        );

    \I__8881\ : InMux
    port map (
            O => \N__39962\,
            I => \N__39953\
        );

    \I__8880\ : InMux
    port map (
            O => \N__39959\,
            I => \N__39953\
        );

    \I__8879\ : InMux
    port map (
            O => \N__39958\,
            I => \N__39950\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__39953\,
            I => \N__39947\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__39950\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__8876\ : Odrv4
    port map (
            O => \N__39947\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__8875\ : InMux
    port map (
            O => \N__39942\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__8874\ : InMux
    port map (
            O => \N__39939\,
            I => \N__39932\
        );

    \I__8873\ : InMux
    port map (
            O => \N__39938\,
            I => \N__39932\
        );

    \I__8872\ : InMux
    port map (
            O => \N__39937\,
            I => \N__39929\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__39932\,
            I => \N__39926\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__39929\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__8869\ : Odrv4
    port map (
            O => \N__39926\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__8868\ : InMux
    port map (
            O => \N__39921\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__8867\ : InMux
    port map (
            O => \N__39918\,
            I => \N__39912\
        );

    \I__8866\ : InMux
    port map (
            O => \N__39917\,
            I => \N__39912\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__39912\,
            I => \N__39908\
        );

    \I__8864\ : InMux
    port map (
            O => \N__39911\,
            I => \N__39905\
        );

    \I__8863\ : Span4Mux_h
    port map (
            O => \N__39908\,
            I => \N__39902\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__39905\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__8861\ : Odrv4
    port map (
            O => \N__39902\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__8860\ : InMux
    port map (
            O => \N__39897\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__8859\ : CascadeMux
    port map (
            O => \N__39894\,
            I => \N__39891\
        );

    \I__8858\ : InMux
    port map (
            O => \N__39891\,
            I => \N__39887\
        );

    \I__8857\ : InMux
    port map (
            O => \N__39890\,
            I => \N__39883\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__39887\,
            I => \N__39880\
        );

    \I__8855\ : InMux
    port map (
            O => \N__39886\,
            I => \N__39877\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__39883\,
            I => \N__39872\
        );

    \I__8853\ : Span4Mux_h
    port map (
            O => \N__39880\,
            I => \N__39872\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__39877\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8851\ : Odrv4
    port map (
            O => \N__39872\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8850\ : InMux
    port map (
            O => \N__39867\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__8849\ : InMux
    port map (
            O => \N__39864\,
            I => \N__39860\
        );

    \I__8848\ : InMux
    port map (
            O => \N__39863\,
            I => \N__39857\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__39860\,
            I => \N__39851\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__39857\,
            I => \N__39851\
        );

    \I__8845\ : InMux
    port map (
            O => \N__39856\,
            I => \N__39848\
        );

    \I__8844\ : Sp12to4
    port map (
            O => \N__39851\,
            I => \N__39842\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__39848\,
            I => \N__39842\
        );

    \I__8842\ : InMux
    port map (
            O => \N__39847\,
            I => \N__39839\
        );

    \I__8841\ : Span12Mux_v
    port map (
            O => \N__39842\,
            I => \N__39836\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__39839\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__8839\ : Odrv12
    port map (
            O => \N__39836\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__8838\ : IoInMux
    port map (
            O => \N__39831\,
            I => \N__39828\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__39828\,
            I => \N__39825\
        );

    \I__8836\ : IoSpan4Mux
    port map (
            O => \N__39825\,
            I => \N__39822\
        );

    \I__8835\ : IoSpan4Mux
    port map (
            O => \N__39822\,
            I => \N__39819\
        );

    \I__8834\ : IoSpan4Mux
    port map (
            O => \N__39819\,
            I => \N__39816\
        );

    \I__8833\ : Odrv4
    port map (
            O => \N__39816\,
            I => \delay_measurement_inst.delay_hc_timer.N_461_i\
        );

    \I__8832\ : InMux
    port map (
            O => \N__39813\,
            I => \N__39810\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__39810\,
            I => \N__39807\
        );

    \I__8830\ : Odrv12
    port map (
            O => \N__39807\,
            I => delay_hc_input_c
        );

    \I__8829\ : InMux
    port map (
            O => \N__39804\,
            I => \N__39801\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__39801\,
            I => delay_hc_d1
        );

    \I__8827\ : InMux
    port map (
            O => \N__39798\,
            I => \bfn_17_8_0_\
        );

    \I__8826\ : CascadeMux
    port map (
            O => \N__39795\,
            I => \N__39792\
        );

    \I__8825\ : InMux
    port map (
            O => \N__39792\,
            I => \N__39789\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__39789\,
            I => \N__39785\
        );

    \I__8823\ : InMux
    port map (
            O => \N__39788\,
            I => \N__39782\
        );

    \I__8822\ : Span4Mux_v
    port map (
            O => \N__39785\,
            I => \N__39778\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__39782\,
            I => \N__39775\
        );

    \I__8820\ : InMux
    port map (
            O => \N__39781\,
            I => \N__39772\
        );

    \I__8819\ : Span4Mux_h
    port map (
            O => \N__39778\,
            I => \N__39769\
        );

    \I__8818\ : Odrv4
    port map (
            O => \N__39775\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__39772\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8816\ : Odrv4
    port map (
            O => \N__39769\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8815\ : InMux
    port map (
            O => \N__39762\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__8814\ : CascadeMux
    port map (
            O => \N__39759\,
            I => \N__39755\
        );

    \I__8813\ : CascadeMux
    port map (
            O => \N__39758\,
            I => \N__39752\
        );

    \I__8812\ : InMux
    port map (
            O => \N__39755\,
            I => \N__39746\
        );

    \I__8811\ : InMux
    port map (
            O => \N__39752\,
            I => \N__39746\
        );

    \I__8810\ : InMux
    port map (
            O => \N__39751\,
            I => \N__39743\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__39746\,
            I => \N__39740\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__39743\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8807\ : Odrv4
    port map (
            O => \N__39740\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8806\ : InMux
    port map (
            O => \N__39735\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__8805\ : InMux
    port map (
            O => \N__39732\,
            I => \N__39725\
        );

    \I__8804\ : InMux
    port map (
            O => \N__39731\,
            I => \N__39725\
        );

    \I__8803\ : InMux
    port map (
            O => \N__39730\,
            I => \N__39722\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__39725\,
            I => \N__39719\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__39722\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8800\ : Odrv4
    port map (
            O => \N__39719\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8799\ : InMux
    port map (
            O => \N__39714\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__8798\ : CascadeMux
    port map (
            O => \N__39711\,
            I => \N__39707\
        );

    \I__8797\ : InMux
    port map (
            O => \N__39710\,
            I => \N__39704\
        );

    \I__8796\ : InMux
    port map (
            O => \N__39707\,
            I => \N__39700\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__39704\,
            I => \N__39697\
        );

    \I__8794\ : InMux
    port map (
            O => \N__39703\,
            I => \N__39694\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__39700\,
            I => \N__39689\
        );

    \I__8792\ : Span4Mux_h
    port map (
            O => \N__39697\,
            I => \N__39689\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__39694\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__8790\ : Odrv4
    port map (
            O => \N__39689\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__8789\ : InMux
    port map (
            O => \N__39684\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__8788\ : CascadeMux
    port map (
            O => \N__39681\,
            I => \N__39678\
        );

    \I__8787\ : InMux
    port map (
            O => \N__39678\,
            I => \N__39674\
        );

    \I__8786\ : InMux
    port map (
            O => \N__39677\,
            I => \N__39670\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__39674\,
            I => \N__39667\
        );

    \I__8784\ : InMux
    port map (
            O => \N__39673\,
            I => \N__39664\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__39670\,
            I => \N__39659\
        );

    \I__8782\ : Span4Mux_h
    port map (
            O => \N__39667\,
            I => \N__39659\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__39664\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8780\ : Odrv4
    port map (
            O => \N__39659\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8779\ : InMux
    port map (
            O => \N__39654\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__8778\ : InMux
    port map (
            O => \N__39651\,
            I => \N__39648\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__39648\,
            I => \N__39644\
        );

    \I__8776\ : InMux
    port map (
            O => \N__39647\,
            I => \N__39641\
        );

    \I__8775\ : Span4Mux_h
    port map (
            O => \N__39644\,
            I => \N__39638\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__39641\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__8773\ : Odrv4
    port map (
            O => \N__39638\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__8772\ : InMux
    port map (
            O => \N__39633\,
            I => \N__39630\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__39630\,
            I => \delay_measurement_inst.delay_hc_timer.N_319\
        );

    \I__8770\ : CascadeMux
    port map (
            O => \N__39627\,
            I => \delay_measurement_inst.N_318_cascade_\
        );

    \I__8769\ : InMux
    port map (
            O => \N__39624\,
            I => \N__39621\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__39621\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__8767\ : InMux
    port map (
            O => \N__39618\,
            I => \N__39615\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__39615\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8765\ : CascadeMux
    port map (
            O => \N__39612\,
            I => \N__39609\
        );

    \I__8764\ : InMux
    port map (
            O => \N__39609\,
            I => \N__39606\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__39606\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__8762\ : InMux
    port map (
            O => \N__39603\,
            I => \N__39600\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__39600\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__8760\ : InMux
    port map (
            O => \N__39597\,
            I => \N__39594\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__39594\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_6_6\
        );

    \I__8758\ : InMux
    port map (
            O => \N__39591\,
            I => \N__39588\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__39588\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__8756\ : InMux
    port map (
            O => \N__39585\,
            I => \N__39582\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__39582\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__8754\ : CascadeMux
    port map (
            O => \N__39579\,
            I => \N__39576\
        );

    \I__8753\ : InMux
    port map (
            O => \N__39576\,
            I => \N__39573\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__39573\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__8751\ : InMux
    port map (
            O => \N__39570\,
            I => \N__39567\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__39567\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__8749\ : InMux
    port map (
            O => \N__39564\,
            I => \N__39561\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__39561\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_7_6\
        );

    \I__8747\ : InMux
    port map (
            O => \N__39558\,
            I => \N__39555\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__39555\,
            I => \N__39551\
        );

    \I__8745\ : InMux
    port map (
            O => \N__39554\,
            I => \N__39548\
        );

    \I__8744\ : Span4Mux_h
    port map (
            O => \N__39551\,
            I => \N__39545\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__39548\,
            I => measured_delay_hc_21
        );

    \I__8742\ : Odrv4
    port map (
            O => \N__39545\,
            I => measured_delay_hc_21
        );

    \I__8741\ : InMux
    port map (
            O => \N__39540\,
            I => \N__39537\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__39537\,
            I => \N__39534\
        );

    \I__8739\ : Odrv4
    port map (
            O => \N__39534\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0Z0Z_19\
        );

    \I__8738\ : InMux
    port map (
            O => \N__39531\,
            I => \N__39527\
        );

    \I__8737\ : InMux
    port map (
            O => \N__39530\,
            I => \N__39524\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__39527\,
            I => \N__39520\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__39524\,
            I => \N__39517\
        );

    \I__8734\ : InMux
    port map (
            O => \N__39523\,
            I => \N__39514\
        );

    \I__8733\ : Span4Mux_h
    port map (
            O => \N__39520\,
            I => \N__39511\
        );

    \I__8732\ : Odrv4
    port map (
            O => \N__39517\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__39514\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__8730\ : Odrv4
    port map (
            O => \N__39511\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__8729\ : CascadeMux
    port map (
            O => \N__39504\,
            I => \N__39500\
        );

    \I__8728\ : InMux
    port map (
            O => \N__39503\,
            I => \N__39497\
        );

    \I__8727\ : InMux
    port map (
            O => \N__39500\,
            I => \N__39494\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__39497\,
            I => \N__39491\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__39494\,
            I => \delay_measurement_inst.delay_hc_timer.N_408\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__39491\,
            I => \delay_measurement_inst.delay_hc_timer.N_408\
        );

    \I__8723\ : CascadeMux
    port map (
            O => \N__39486\,
            I => \N__39483\
        );

    \I__8722\ : InMux
    port map (
            O => \N__39483\,
            I => \N__39480\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__39480\,
            I => \N__39476\
        );

    \I__8720\ : InMux
    port map (
            O => \N__39479\,
            I => \N__39473\
        );

    \I__8719\ : Span4Mux_h
    port map (
            O => \N__39476\,
            I => \N__39470\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__39473\,
            I => measured_delay_hc_26
        );

    \I__8717\ : Odrv4
    port map (
            O => \N__39470\,
            I => measured_delay_hc_26
        );

    \I__8716\ : InMux
    port map (
            O => \N__39465\,
            I => \N__39461\
        );

    \I__8715\ : CascadeMux
    port map (
            O => \N__39464\,
            I => \N__39457\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__39461\,
            I => \N__39454\
        );

    \I__8713\ : InMux
    port map (
            O => \N__39460\,
            I => \N__39451\
        );

    \I__8712\ : InMux
    port map (
            O => \N__39457\,
            I => \N__39448\
        );

    \I__8711\ : Odrv4
    port map (
            O => \N__39454\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__39451\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__39448\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__8708\ : InMux
    port map (
            O => \N__39441\,
            I => \N__39437\
        );

    \I__8707\ : InMux
    port map (
            O => \N__39440\,
            I => \N__39434\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__39437\,
            I => measured_delay_hc_20
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__39434\,
            I => measured_delay_hc_20
        );

    \I__8704\ : InMux
    port map (
            O => \N__39429\,
            I => \N__39426\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__39426\,
            I => \N__39421\
        );

    \I__8702\ : InMux
    port map (
            O => \N__39425\,
            I => \N__39418\
        );

    \I__8701\ : InMux
    port map (
            O => \N__39424\,
            I => \N__39415\
        );

    \I__8700\ : Odrv12
    port map (
            O => \N__39421\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__39418\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__39415\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__8697\ : InMux
    port map (
            O => \N__39408\,
            I => \N__39405\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__39405\,
            I => \N__39401\
        );

    \I__8695\ : CascadeMux
    port map (
            O => \N__39404\,
            I => \N__39398\
        );

    \I__8694\ : Span4Mux_v
    port map (
            O => \N__39401\,
            I => \N__39394\
        );

    \I__8693\ : InMux
    port map (
            O => \N__39398\,
            I => \N__39389\
        );

    \I__8692\ : InMux
    port map (
            O => \N__39397\,
            I => \N__39389\
        );

    \I__8691\ : Odrv4
    port map (
            O => \N__39394\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__39389\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__8689\ : CascadeMux
    port map (
            O => \N__39384\,
            I => \delay_measurement_inst.delay_hc_timer.N_318_1_cascade_\
        );

    \I__8688\ : InMux
    port map (
            O => \N__39381\,
            I => \N__39378\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__39378\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_6\
        );

    \I__8686\ : InMux
    port map (
            O => \N__39375\,
            I => \N__39372\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__39372\,
            I => \N__39369\
        );

    \I__8684\ : Odrv4
    port map (
            O => \N__39369\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_5\
        );

    \I__8683\ : CascadeMux
    port map (
            O => \N__39366\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_9_cascade_\
        );

    \I__8682\ : InMux
    port map (
            O => \N__39363\,
            I => \N__39360\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__39360\,
            I => \delay_measurement_inst.delay_hc_timer.N_440\
        );

    \I__8680\ : InMux
    port map (
            O => \N__39357\,
            I => \N__39354\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__39354\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__8678\ : InMux
    port map (
            O => \N__39351\,
            I => \N__39348\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__39348\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__8676\ : InMux
    port map (
            O => \N__39345\,
            I => \N__39342\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__39342\,
            I => \N__39339\
        );

    \I__8674\ : Odrv4
    port map (
            O => \N__39339\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__8673\ : CascadeMux
    port map (
            O => \N__39336\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_0_6_cascade_\
        );

    \I__8672\ : CascadeMux
    port map (
            O => \N__39333\,
            I => \delay_measurement_inst.delay_hc_timer.N_328_cascade_\
        );

    \I__8671\ : InMux
    port map (
            O => \N__39330\,
            I => \N__39327\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__39327\,
            I => \N__39324\
        );

    \I__8669\ : Odrv4
    port map (
            O => \N__39324\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_4\
        );

    \I__8668\ : InMux
    port map (
            O => \N__39321\,
            I => \N__39318\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__39318\,
            I => \delay_measurement_inst.delay_hc_timer.N_318_1\
        );

    \I__8666\ : InMux
    port map (
            O => \N__39315\,
            I => \N__39309\
        );

    \I__8665\ : InMux
    port map (
            O => \N__39314\,
            I => \N__39309\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__39309\,
            I => \N__39304\
        );

    \I__8663\ : InMux
    port map (
            O => \N__39308\,
            I => \N__39299\
        );

    \I__8662\ : InMux
    port map (
            O => \N__39307\,
            I => \N__39299\
        );

    \I__8661\ : Odrv4
    port map (
            O => \N__39304\,
            I => \delay_measurement_inst.delay_hc_timer.N_331\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__39299\,
            I => \delay_measurement_inst.delay_hc_timer.N_331\
        );

    \I__8659\ : InMux
    port map (
            O => \N__39294\,
            I => \N__39290\
        );

    \I__8658\ : InMux
    port map (
            O => \N__39293\,
            I => \N__39287\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__39290\,
            I => \delay_measurement_inst.delay_hc_timer.N_328\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__39287\,
            I => \delay_measurement_inst.delay_hc_timer.N_328\
        );

    \I__8655\ : InMux
    port map (
            O => \N__39282\,
            I => \N__39279\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__39279\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2Z0Z_18\
        );

    \I__8653\ : InMux
    port map (
            O => \N__39276\,
            I => \N__39273\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__39273\,
            I => \N__39270\
        );

    \I__8651\ : Span4Mux_v
    port map (
            O => \N__39270\,
            I => \N__39266\
        );

    \I__8650\ : InMux
    port map (
            O => \N__39269\,
            I => \N__39263\
        );

    \I__8649\ : Odrv4
    port map (
            O => \N__39266\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__39263\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__8647\ : InMux
    port map (
            O => \N__39258\,
            I => \N__39255\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__39255\,
            I => \N__39252\
        );

    \I__8645\ : Span4Mux_v
    port map (
            O => \N__39252\,
            I => \N__39248\
        );

    \I__8644\ : InMux
    port map (
            O => \N__39251\,
            I => \N__39245\
        );

    \I__8643\ : Odrv4
    port map (
            O => \N__39248\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__39245\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__8641\ : InMux
    port map (
            O => \N__39240\,
            I => \N__39237\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__39237\,
            I => \N__39233\
        );

    \I__8639\ : CascadeMux
    port map (
            O => \N__39236\,
            I => \N__39230\
        );

    \I__8638\ : Span4Mux_h
    port map (
            O => \N__39233\,
            I => \N__39227\
        );

    \I__8637\ : InMux
    port map (
            O => \N__39230\,
            I => \N__39224\
        );

    \I__8636\ : Odrv4
    port map (
            O => \N__39227\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__39224\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__8634\ : InMux
    port map (
            O => \N__39219\,
            I => \N__39216\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__39216\,
            I => \N__39212\
        );

    \I__8632\ : InMux
    port map (
            O => \N__39215\,
            I => \N__39209\
        );

    \I__8631\ : Odrv4
    port map (
            O => \N__39212\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__39209\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__8629\ : InMux
    port map (
            O => \N__39204\,
            I => \N__39200\
        );

    \I__8628\ : InMux
    port map (
            O => \N__39203\,
            I => \N__39197\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__39200\,
            I => \N__39194\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__39197\,
            I => measured_delay_hc_24
        );

    \I__8625\ : Odrv4
    port map (
            O => \N__39194\,
            I => measured_delay_hc_24
        );

    \I__8624\ : InMux
    port map (
            O => \N__39189\,
            I => \N__39185\
        );

    \I__8623\ : InMux
    port map (
            O => \N__39188\,
            I => \N__39182\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__39185\,
            I => \N__39179\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__39182\,
            I => measured_delay_hc_23
        );

    \I__8620\ : Odrv12
    port map (
            O => \N__39179\,
            I => measured_delay_hc_23
        );

    \I__8619\ : InMux
    port map (
            O => \N__39174\,
            I => \N__39170\
        );

    \I__8618\ : InMux
    port map (
            O => \N__39173\,
            I => \N__39167\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__39170\,
            I => \N__39164\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__39167\,
            I => measured_delay_hc_22
        );

    \I__8615\ : Odrv12
    port map (
            O => \N__39164\,
            I => measured_delay_hc_22
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__39159\,
            I => \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7Z0Z_19_cascade_\
        );

    \I__8613\ : InMux
    port map (
            O => \N__39156\,
            I => \N__39151\
        );

    \I__8612\ : InMux
    port map (
            O => \N__39155\,
            I => \N__39148\
        );

    \I__8611\ : InMux
    port map (
            O => \N__39154\,
            I => \N__39145\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__39151\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__39148\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__39145\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__8607\ : InMux
    port map (
            O => \N__39138\,
            I => \N__39133\
        );

    \I__8606\ : InMux
    port map (
            O => \N__39137\,
            I => \N__39130\
        );

    \I__8605\ : InMux
    port map (
            O => \N__39136\,
            I => \N__39127\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__39133\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__39130\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__39127\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__8601\ : CascadeMux
    port map (
            O => \N__39120\,
            I => \delay_measurement_inst.delay_hc_timer.N_299_cascade_\
        );

    \I__8600\ : InMux
    port map (
            O => \N__39117\,
            I => \N__39114\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__39114\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_2_6\
        );

    \I__8598\ : CascadeMux
    port map (
            O => \N__39111\,
            I => \delay_measurement_inst.N_332_cascade_\
        );

    \I__8597\ : InMux
    port map (
            O => \N__39108\,
            I => \N__39105\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__39105\,
            I => \phase_controller_inst1.stoper_hc.N_406\
        );

    \I__8595\ : CascadeMux
    port map (
            O => \N__39102\,
            I => \phase_controller_inst1.stoper_hc.N_406_cascade_\
        );

    \I__8594\ : InMux
    port map (
            O => \N__39099\,
            I => \N__39094\
        );

    \I__8593\ : InMux
    port map (
            O => \N__39098\,
            I => \N__39091\
        );

    \I__8592\ : InMux
    port map (
            O => \N__39097\,
            I => \N__39088\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__39094\,
            I => \N__39085\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__39091\,
            I => \N__39082\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__39088\,
            I => \N__39079\
        );

    \I__8588\ : Span4Mux_v
    port map (
            O => \N__39085\,
            I => \N__39075\
        );

    \I__8587\ : Span4Mux_v
    port map (
            O => \N__39082\,
            I => \N__39070\
        );

    \I__8586\ : Span4Mux_v
    port map (
            O => \N__39079\,
            I => \N__39070\
        );

    \I__8585\ : InMux
    port map (
            O => \N__39078\,
            I => \N__39067\
        );

    \I__8584\ : Odrv4
    port map (
            O => \N__39075\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__8583\ : Odrv4
    port map (
            O => \N__39070\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__39067\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__8581\ : InMux
    port map (
            O => \N__39060\,
            I => \N__39057\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__39057\,
            I => \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_8\
        );

    \I__8579\ : CascadeMux
    port map (
            O => \N__39054\,
            I => \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_7_cascade_\
        );

    \I__8578\ : InMux
    port map (
            O => \N__39051\,
            I => \N__39048\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__39048\,
            I => \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_5\
        );

    \I__8576\ : InMux
    port map (
            O => \N__39045\,
            I => \N__39042\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__39042\,
            I => \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_6\
        );

    \I__8574\ : CascadeMux
    port map (
            O => \N__39039\,
            I => \N__39036\
        );

    \I__8573\ : InMux
    port map (
            O => \N__39036\,
            I => \N__39033\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__39033\,
            I => \N__39030\
        );

    \I__8571\ : Odrv4
    port map (
            O => \N__39030\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__8570\ : CascadeMux
    port map (
            O => \N__39027\,
            I => \N__39024\
        );

    \I__8569\ : InMux
    port map (
            O => \N__39024\,
            I => \N__39021\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__39021\,
            I => \N__39018\
        );

    \I__8567\ : Span4Mux_h
    port map (
            O => \N__39018\,
            I => \N__39015\
        );

    \I__8566\ : Odrv4
    port map (
            O => \N__39015\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__8565\ : CascadeMux
    port map (
            O => \N__39012\,
            I => \N__39009\
        );

    \I__8564\ : InMux
    port map (
            O => \N__39009\,
            I => \N__39006\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__39006\,
            I => \N__39003\
        );

    \I__8562\ : Span4Mux_h
    port map (
            O => \N__39003\,
            I => \N__39000\
        );

    \I__8561\ : Span4Mux_h
    port map (
            O => \N__39000\,
            I => \N__38997\
        );

    \I__8560\ : Odrv4
    port map (
            O => \N__38997\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__8559\ : CascadeMux
    port map (
            O => \N__38994\,
            I => \N__38991\
        );

    \I__8558\ : InMux
    port map (
            O => \N__38991\,
            I => \N__38988\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__38988\,
            I => \N__38985\
        );

    \I__8556\ : Span4Mux_h
    port map (
            O => \N__38985\,
            I => \N__38982\
        );

    \I__8555\ : Odrv4
    port map (
            O => \N__38982\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__8554\ : CascadeMux
    port map (
            O => \N__38979\,
            I => \N__38976\
        );

    \I__8553\ : InMux
    port map (
            O => \N__38976\,
            I => \N__38973\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__38973\,
            I => \N__38970\
        );

    \I__8551\ : Odrv12
    port map (
            O => \N__38970\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__8550\ : CascadeMux
    port map (
            O => \N__38967\,
            I => \N__38964\
        );

    \I__8549\ : InMux
    port map (
            O => \N__38964\,
            I => \N__38961\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__38961\,
            I => \N__38958\
        );

    \I__8547\ : Span4Mux_h
    port map (
            O => \N__38958\,
            I => \N__38955\
        );

    \I__8546\ : Odrv4
    port map (
            O => \N__38955\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__8545\ : CascadeMux
    port map (
            O => \N__38952\,
            I => \N__38949\
        );

    \I__8544\ : InMux
    port map (
            O => \N__38949\,
            I => \N__38946\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__38946\,
            I => \N__38943\
        );

    \I__8542\ : Span4Mux_h
    port map (
            O => \N__38943\,
            I => \N__38940\
        );

    \I__8541\ : Odrv4
    port map (
            O => \N__38940\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__8540\ : CEMux
    port map (
            O => \N__38937\,
            I => \N__38934\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__38934\,
            I => \N__38929\
        );

    \I__8538\ : CEMux
    port map (
            O => \N__38933\,
            I => \N__38926\
        );

    \I__8537\ : CEMux
    port map (
            O => \N__38932\,
            I => \N__38922\
        );

    \I__8536\ : Span4Mux_h
    port map (
            O => \N__38929\,
            I => \N__38917\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__38926\,
            I => \N__38917\
        );

    \I__8534\ : CEMux
    port map (
            O => \N__38925\,
            I => \N__38914\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__38922\,
            I => \N__38911\
        );

    \I__8532\ : Span4Mux_v
    port map (
            O => \N__38917\,
            I => \N__38906\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__38914\,
            I => \N__38906\
        );

    \I__8530\ : Span4Mux_v
    port map (
            O => \N__38911\,
            I => \N__38903\
        );

    \I__8529\ : Span4Mux_h
    port map (
            O => \N__38906\,
            I => \N__38900\
        );

    \I__8528\ : Span4Mux_v
    port map (
            O => \N__38903\,
            I => \N__38897\
        );

    \I__8527\ : Span4Mux_v
    port map (
            O => \N__38900\,
            I => \N__38894\
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__38897\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__8525\ : Odrv4
    port map (
            O => \N__38894\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__8524\ : CascadeMux
    port map (
            O => \N__38889\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0Z0Z_3_cascade_\
        );

    \I__8523\ : CascadeMux
    port map (
            O => \N__38886\,
            I => \phase_controller_inst1.stoper_hc.N_316_cascade_\
        );

    \I__8522\ : CascadeMux
    port map (
            O => \N__38883\,
            I => \N__38880\
        );

    \I__8521\ : InMux
    port map (
            O => \N__38880\,
            I => \N__38877\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__38877\,
            I => \N__38874\
        );

    \I__8519\ : Odrv4
    port map (
            O => \N__38874\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\
        );

    \I__8518\ : InMux
    port map (
            O => \N__38871\,
            I => \N__38867\
        );

    \I__8517\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38864\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__38867\,
            I => \N__38861\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__38864\,
            I => \N__38856\
        );

    \I__8514\ : Span4Mux_h
    port map (
            O => \N__38861\,
            I => \N__38856\
        );

    \I__8513\ : Odrv4
    port map (
            O => \N__38856\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__8512\ : InMux
    port map (
            O => \N__38853\,
            I => \N__38850\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__38850\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\
        );

    \I__8510\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38844\
        );

    \I__8509\ : LocalMux
    port map (
            O => \N__38844\,
            I => \N__38840\
        );

    \I__8508\ : InMux
    port map (
            O => \N__38843\,
            I => \N__38837\
        );

    \I__8507\ : Span4Mux_h
    port map (
            O => \N__38840\,
            I => \N__38834\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__38837\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__8505\ : Odrv4
    port map (
            O => \N__38834\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__8504\ : CascadeMux
    port map (
            O => \N__38829\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31_5_cascade_\
        );

    \I__8503\ : InMux
    port map (
            O => \N__38826\,
            I => \N__38823\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__38823\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__8501\ : InMux
    port map (
            O => \N__38820\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__8500\ : InMux
    port map (
            O => \N__38817\,
            I => \N__38814\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__38814\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__8498\ : InMux
    port map (
            O => \N__38811\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__8497\ : CascadeMux
    port map (
            O => \N__38808\,
            I => \N__38805\
        );

    \I__8496\ : InMux
    port map (
            O => \N__38805\,
            I => \N__38802\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__38802\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__8494\ : InMux
    port map (
            O => \N__38799\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__8493\ : InMux
    port map (
            O => \N__38796\,
            I => \N__38793\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__38793\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__8491\ : InMux
    port map (
            O => \N__38790\,
            I => \bfn_16_14_0_\
        );

    \I__8490\ : InMux
    port map (
            O => \N__38787\,
            I => \N__38784\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__38784\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__8488\ : InMux
    port map (
            O => \N__38781\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__8487\ : InMux
    port map (
            O => \N__38778\,
            I => \N__38775\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__38775\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__8485\ : InMux
    port map (
            O => \N__38772\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__8484\ : CascadeMux
    port map (
            O => \N__38769\,
            I => \N__38766\
        );

    \I__8483\ : InMux
    port map (
            O => \N__38766\,
            I => \N__38763\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__38763\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\
        );

    \I__8481\ : InMux
    port map (
            O => \N__38760\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__8480\ : InMux
    port map (
            O => \N__38757\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__8479\ : InMux
    port map (
            O => \N__38754\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__8478\ : InMux
    port map (
            O => \N__38751\,
            I => \N__38746\
        );

    \I__8477\ : InMux
    port map (
            O => \N__38750\,
            I => \N__38743\
        );

    \I__8476\ : InMux
    port map (
            O => \N__38749\,
            I => \N__38740\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__38746\,
            I => \N__38733\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__38743\,
            I => \N__38733\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__38740\,
            I => \N__38733\
        );

    \I__8472\ : Odrv4
    port map (
            O => \N__38733\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__8471\ : InMux
    port map (
            O => \N__38730\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__8470\ : InMux
    port map (
            O => \N__38727\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__8469\ : InMux
    port map (
            O => \N__38724\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__8468\ : CascadeMux
    port map (
            O => \N__38721\,
            I => \N__38716\
        );

    \I__8467\ : InMux
    port map (
            O => \N__38720\,
            I => \N__38713\
        );

    \I__8466\ : InMux
    port map (
            O => \N__38719\,
            I => \N__38708\
        );

    \I__8465\ : InMux
    port map (
            O => \N__38716\,
            I => \N__38708\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__38713\,
            I => \N__38705\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__38708\,
            I => \N__38702\
        );

    \I__8462\ : Odrv12
    port map (
            O => \N__38705\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__8461\ : Odrv12
    port map (
            O => \N__38702\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__8460\ : InMux
    port map (
            O => \N__38697\,
            I => \bfn_16_13_0_\
        );

    \I__8459\ : InMux
    port map (
            O => \N__38694\,
            I => \N__38691\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__38691\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__8457\ : InMux
    port map (
            O => \N__38688\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__8456\ : InMux
    port map (
            O => \N__38685\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__8455\ : InMux
    port map (
            O => \N__38682\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__8454\ : InMux
    port map (
            O => \N__38679\,
            I => \N__38676\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__38676\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__8452\ : InMux
    port map (
            O => \N__38673\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__8451\ : InMux
    port map (
            O => \N__38670\,
            I => \N__38667\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__38667\,
            I => \N__38664\
        );

    \I__8449\ : Span4Mux_h
    port map (
            O => \N__38664\,
            I => \N__38660\
        );

    \I__8448\ : InMux
    port map (
            O => \N__38663\,
            I => \N__38657\
        );

    \I__8447\ : Odrv4
    port map (
            O => \N__38660\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__38657\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__8445\ : InMux
    port map (
            O => \N__38652\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__8444\ : InMux
    port map (
            O => \N__38649\,
            I => \N__38646\
        );

    \I__8443\ : LocalMux
    port map (
            O => \N__38646\,
            I => \N__38643\
        );

    \I__8442\ : Span4Mux_h
    port map (
            O => \N__38643\,
            I => \N__38639\
        );

    \I__8441\ : InMux
    port map (
            O => \N__38642\,
            I => \N__38636\
        );

    \I__8440\ : Odrv4
    port map (
            O => \N__38639\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__38636\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__8438\ : InMux
    port map (
            O => \N__38631\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__8437\ : InMux
    port map (
            O => \N__38628\,
            I => \N__38624\
        );

    \I__8436\ : InMux
    port map (
            O => \N__38627\,
            I => \N__38621\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__38624\,
            I => \N__38616\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__38621\,
            I => \N__38616\
        );

    \I__8433\ : Span4Mux_h
    port map (
            O => \N__38616\,
            I => \N__38610\
        );

    \I__8432\ : InMux
    port map (
            O => \N__38615\,
            I => \N__38607\
        );

    \I__8431\ : InMux
    port map (
            O => \N__38614\,
            I => \N__38604\
        );

    \I__8430\ : InMux
    port map (
            O => \N__38613\,
            I => \N__38601\
        );

    \I__8429\ : Odrv4
    port map (
            O => \N__38610\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__38607\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__38604\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__38601\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__8425\ : InMux
    port map (
            O => \N__38592\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__8424\ : InMux
    port map (
            O => \N__38589\,
            I => \N__38586\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__38586\,
            I => \N__38583\
        );

    \I__8422\ : Span4Mux_v
    port map (
            O => \N__38583\,
            I => \N__38579\
        );

    \I__8421\ : InMux
    port map (
            O => \N__38582\,
            I => \N__38576\
        );

    \I__8420\ : Odrv4
    port map (
            O => \N__38579\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__38576\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__8418\ : InMux
    port map (
            O => \N__38571\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__8417\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38565\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__38565\,
            I => \N__38561\
        );

    \I__8415\ : InMux
    port map (
            O => \N__38564\,
            I => \N__38558\
        );

    \I__8414\ : Odrv4
    port map (
            O => \N__38561\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__38558\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__8412\ : InMux
    port map (
            O => \N__38553\,
            I => \bfn_16_12_0_\
        );

    \I__8411\ : InMux
    port map (
            O => \N__38550\,
            I => \N__38547\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__38547\,
            I => \N__38543\
        );

    \I__8409\ : InMux
    port map (
            O => \N__38546\,
            I => \N__38540\
        );

    \I__8408\ : Odrv4
    port map (
            O => \N__38543\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__38540\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__8406\ : InMux
    port map (
            O => \N__38535\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__8405\ : InMux
    port map (
            O => \N__38532\,
            I => \N__38528\
        );

    \I__8404\ : CascadeMux
    port map (
            O => \N__38531\,
            I => \N__38525\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__38528\,
            I => \N__38522\
        );

    \I__8402\ : InMux
    port map (
            O => \N__38525\,
            I => \N__38519\
        );

    \I__8401\ : Odrv4
    port map (
            O => \N__38522\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__38519\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__8399\ : InMux
    port map (
            O => \N__38514\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__8398\ : InMux
    port map (
            O => \N__38511\,
            I => \N__38505\
        );

    \I__8397\ : InMux
    port map (
            O => \N__38510\,
            I => \N__38502\
        );

    \I__8396\ : InMux
    port map (
            O => \N__38509\,
            I => \N__38498\
        );

    \I__8395\ : InMux
    port map (
            O => \N__38508\,
            I => \N__38495\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__38505\,
            I => \N__38490\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__38502\,
            I => \N__38490\
        );

    \I__8392\ : InMux
    port map (
            O => \N__38501\,
            I => \N__38487\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__38498\,
            I => \N__38484\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__38495\,
            I => \N__38481\
        );

    \I__8389\ : Odrv4
    port map (
            O => \N__38490\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__38487\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__8387\ : Odrv12
    port map (
            O => \N__38484\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__8386\ : Odrv4
    port map (
            O => \N__38481\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__8385\ : InMux
    port map (
            O => \N__38472\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__8384\ : CascadeMux
    port map (
            O => \N__38469\,
            I => \N__38465\
        );

    \I__8383\ : CascadeMux
    port map (
            O => \N__38468\,
            I => \N__38461\
        );

    \I__8382\ : InMux
    port map (
            O => \N__38465\,
            I => \N__38453\
        );

    \I__8381\ : InMux
    port map (
            O => \N__38464\,
            I => \N__38453\
        );

    \I__8380\ : InMux
    port map (
            O => \N__38461\,
            I => \N__38448\
        );

    \I__8379\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38443\
        );

    \I__8378\ : InMux
    port map (
            O => \N__38459\,
            I => \N__38443\
        );

    \I__8377\ : CascadeMux
    port map (
            O => \N__38458\,
            I => \N__38439\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__38453\,
            I => \N__38436\
        );

    \I__8375\ : InMux
    port map (
            O => \N__38452\,
            I => \N__38431\
        );

    \I__8374\ : InMux
    port map (
            O => \N__38451\,
            I => \N__38431\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__38448\,
            I => \N__38428\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__38443\,
            I => \N__38425\
        );

    \I__8371\ : InMux
    port map (
            O => \N__38442\,
            I => \N__38420\
        );

    \I__8370\ : InMux
    port map (
            O => \N__38439\,
            I => \N__38420\
        );

    \I__8369\ : Span4Mux_v
    port map (
            O => \N__38436\,
            I => \N__38415\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__38431\,
            I => \N__38415\
        );

    \I__8367\ : Span4Mux_h
    port map (
            O => \N__38428\,
            I => \N__38412\
        );

    \I__8366\ : Odrv4
    port map (
            O => \N__38425\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__38420\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__8364\ : Odrv4
    port map (
            O => \N__38415\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__8363\ : Odrv4
    port map (
            O => \N__38412\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__8362\ : InMux
    port map (
            O => \N__38403\,
            I => \N__38398\
        );

    \I__8361\ : InMux
    port map (
            O => \N__38402\,
            I => \N__38395\
        );

    \I__8360\ : InMux
    port map (
            O => \N__38401\,
            I => \N__38392\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__38398\,
            I => \N__38389\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__38395\,
            I => \N__38386\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__38392\,
            I => \N__38381\
        );

    \I__8356\ : Span4Mux_v
    port map (
            O => \N__38389\,
            I => \N__38381\
        );

    \I__8355\ : Odrv12
    port map (
            O => \N__38386\,
            I => \il_min_comp1_D2\
        );

    \I__8354\ : Odrv4
    port map (
            O => \N__38381\,
            I => \il_min_comp1_D2\
        );

    \I__8353\ : InMux
    port map (
            O => \N__38376\,
            I => \N__38373\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__38373\,
            I => \N__38370\
        );

    \I__8351\ : Odrv4
    port map (
            O => \N__38370\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__8350\ : InMux
    port map (
            O => \N__38367\,
            I => \N__38364\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__38364\,
            I => \N__38360\
        );

    \I__8348\ : InMux
    port map (
            O => \N__38363\,
            I => \N__38357\
        );

    \I__8347\ : Span4Mux_v
    port map (
            O => \N__38360\,
            I => \N__38351\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__38357\,
            I => \N__38351\
        );

    \I__8345\ : InMux
    port map (
            O => \N__38356\,
            I => \N__38348\
        );

    \I__8344\ : Span4Mux_v
    port map (
            O => \N__38351\,
            I => \N__38345\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__38348\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__8342\ : Odrv4
    port map (
            O => \N__38345\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__8341\ : CascadeMux
    port map (
            O => \N__38340\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\
        );

    \I__8340\ : InMux
    port map (
            O => \N__38337\,
            I => \N__38334\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__38334\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\
        );

    \I__8338\ : InMux
    port map (
            O => \N__38331\,
            I => \N__38325\
        );

    \I__8337\ : InMux
    port map (
            O => \N__38330\,
            I => \N__38325\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__38325\,
            I => \delay_measurement_inst.delay_tr_timer.N_373_4\
        );

    \I__8335\ : InMux
    port map (
            O => \N__38322\,
            I => \N__38319\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__38319\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\
        );

    \I__8333\ : InMux
    port map (
            O => \N__38316\,
            I => \N__38313\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__38313\,
            I => \N__38308\
        );

    \I__8331\ : InMux
    port map (
            O => \N__38312\,
            I => \N__38303\
        );

    \I__8330\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38303\
        );

    \I__8329\ : Odrv4
    port map (
            O => \N__38308\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__38303\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__8327\ : InMux
    port map (
            O => \N__38298\,
            I => \N__38295\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__38295\,
            I => \N__38291\
        );

    \I__8325\ : InMux
    port map (
            O => \N__38294\,
            I => \N__38288\
        );

    \I__8324\ : Odrv4
    port map (
            O => \N__38291\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__38288\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__8322\ : InMux
    port map (
            O => \N__38283\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__8321\ : InMux
    port map (
            O => \N__38280\,
            I => \N__38277\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__38277\,
            I => \N__38273\
        );

    \I__8319\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38270\
        );

    \I__8318\ : Odrv4
    port map (
            O => \N__38273\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__38270\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__8316\ : InMux
    port map (
            O => \N__38265\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__8315\ : InMux
    port map (
            O => \N__38262\,
            I => \N__38256\
        );

    \I__8314\ : InMux
    port map (
            O => \N__38261\,
            I => \N__38253\
        );

    \I__8313\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38250\
        );

    \I__8312\ : InMux
    port map (
            O => \N__38259\,
            I => \N__38247\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__38256\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__38253\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__38250\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__38247\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__8307\ : InMux
    port map (
            O => \N__38238\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__8306\ : CascadeMux
    port map (
            O => \N__38235\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_\
        );

    \I__8305\ : InMux
    port map (
            O => \N__38232\,
            I => \N__38227\
        );

    \I__8304\ : InMux
    port map (
            O => \N__38231\,
            I => \N__38224\
        );

    \I__8303\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38221\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__38227\,
            I => \N__38218\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__38224\,
            I => \N__38214\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__38221\,
            I => \N__38210\
        );

    \I__8299\ : Span4Mux_v
    port map (
            O => \N__38218\,
            I => \N__38207\
        );

    \I__8298\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38204\
        );

    \I__8297\ : Span4Mux_h
    port map (
            O => \N__38214\,
            I => \N__38201\
        );

    \I__8296\ : InMux
    port map (
            O => \N__38213\,
            I => \N__38198\
        );

    \I__8295\ : Span4Mux_v
    port map (
            O => \N__38210\,
            I => \N__38195\
        );

    \I__8294\ : Span4Mux_h
    port map (
            O => \N__38207\,
            I => \N__38190\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__38204\,
            I => \N__38190\
        );

    \I__8292\ : Span4Mux_h
    port map (
            O => \N__38201\,
            I => \N__38187\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__38198\,
            I => \N__38183\
        );

    \I__8290\ : Span4Mux_h
    port map (
            O => \N__38195\,
            I => \N__38178\
        );

    \I__8289\ : Span4Mux_v
    port map (
            O => \N__38190\,
            I => \N__38178\
        );

    \I__8288\ : Sp12to4
    port map (
            O => \N__38187\,
            I => \N__38175\
        );

    \I__8287\ : InMux
    port map (
            O => \N__38186\,
            I => \N__38172\
        );

    \I__8286\ : Span4Mux_v
    port map (
            O => \N__38183\,
            I => \N__38167\
        );

    \I__8285\ : Span4Mux_h
    port map (
            O => \N__38178\,
            I => \N__38167\
        );

    \I__8284\ : Odrv12
    port map (
            O => \N__38175\,
            I => phase_controller_inst1_state_4
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__38172\,
            I => phase_controller_inst1_state_4
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__38167\,
            I => phase_controller_inst1_state_4
        );

    \I__8281\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38157\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__38157\,
            I => \N__38153\
        );

    \I__8279\ : InMux
    port map (
            O => \N__38156\,
            I => \N__38150\
        );

    \I__8278\ : Span4Mux_h
    port map (
            O => \N__38153\,
            I => \N__38146\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__38150\,
            I => \N__38143\
        );

    \I__8276\ : InMux
    port map (
            O => \N__38149\,
            I => \N__38140\
        );

    \I__8275\ : Odrv4
    port map (
            O => \N__38146\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__8274\ : Odrv12
    port map (
            O => \N__38143\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__38140\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__8272\ : CascadeMux
    port map (
            O => \N__38133\,
            I => \N__38130\
        );

    \I__8271\ : InMux
    port map (
            O => \N__38130\,
            I => \N__38127\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__38127\,
            I => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__8269\ : InMux
    port map (
            O => \N__38124\,
            I => \N__38121\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__38121\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\
        );

    \I__8267\ : InMux
    port map (
            O => \N__38118\,
            I => \N__38115\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__38115\,
            I => \N__38111\
        );

    \I__8265\ : InMux
    port map (
            O => \N__38114\,
            I => \N__38108\
        );

    \I__8264\ : Span4Mux_v
    port map (
            O => \N__38111\,
            I => \N__38105\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__38108\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8262\ : Odrv4
    port map (
            O => \N__38105\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8261\ : CascadeMux
    port map (
            O => \N__38100\,
            I => \N__38096\
        );

    \I__8260\ : InMux
    port map (
            O => \N__38099\,
            I => \N__38088\
        );

    \I__8259\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38088\
        );

    \I__8258\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38088\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__38088\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__8256\ : InMux
    port map (
            O => \N__38085\,
            I => \N__38079\
        );

    \I__8255\ : InMux
    port map (
            O => \N__38084\,
            I => \N__38079\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__38079\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__8253\ : InMux
    port map (
            O => \N__38076\,
            I => \N__38070\
        );

    \I__8252\ : InMux
    port map (
            O => \N__38075\,
            I => \N__38067\
        );

    \I__8251\ : InMux
    port map (
            O => \N__38074\,
            I => \N__38062\
        );

    \I__8250\ : InMux
    port map (
            O => \N__38073\,
            I => \N__38062\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__38070\,
            I => \N__38059\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__38067\,
            I => \N__38054\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__38062\,
            I => \N__38054\
        );

    \I__8246\ : Span12Mux_h
    port map (
            O => \N__38059\,
            I => \N__38051\
        );

    \I__8245\ : Span4Mux_h
    port map (
            O => \N__38054\,
            I => \N__38048\
        );

    \I__8244\ : Odrv12
    port map (
            O => \N__38051\,
            I => measured_delay_tr_16
        );

    \I__8243\ : Odrv4
    port map (
            O => \N__38048\,
            I => measured_delay_tr_16
        );

    \I__8242\ : InMux
    port map (
            O => \N__38043\,
            I => \N__38038\
        );

    \I__8241\ : CascadeMux
    port map (
            O => \N__38042\,
            I => \N__38034\
        );

    \I__8240\ : CascadeMux
    port map (
            O => \N__38041\,
            I => \N__38031\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__38038\,
            I => \N__38028\
        );

    \I__8238\ : InMux
    port map (
            O => \N__38037\,
            I => \N__38025\
        );

    \I__8237\ : InMux
    port map (
            O => \N__38034\,
            I => \N__38020\
        );

    \I__8236\ : InMux
    port map (
            O => \N__38031\,
            I => \N__38020\
        );

    \I__8235\ : Span4Mux_v
    port map (
            O => \N__38028\,
            I => \N__38017\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__38025\,
            I => \N__38014\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__38020\,
            I => \N__38011\
        );

    \I__8232\ : Span4Mux_h
    port map (
            O => \N__38017\,
            I => \N__38008\
        );

    \I__8231\ : Span4Mux_h
    port map (
            O => \N__38014\,
            I => \N__38005\
        );

    \I__8230\ : Span4Mux_h
    port map (
            O => \N__38011\,
            I => \N__38002\
        );

    \I__8229\ : Odrv4
    port map (
            O => \N__38008\,
            I => measured_delay_tr_19
        );

    \I__8228\ : Odrv4
    port map (
            O => \N__38005\,
            I => measured_delay_tr_19
        );

    \I__8227\ : Odrv4
    port map (
            O => \N__38002\,
            I => measured_delay_tr_19
        );

    \I__8226\ : CascadeMux
    port map (
            O => \N__37995\,
            I => \N__37990\
        );

    \I__8225\ : InMux
    port map (
            O => \N__37994\,
            I => \N__37985\
        );

    \I__8224\ : InMux
    port map (
            O => \N__37993\,
            I => \N__37985\
        );

    \I__8223\ : InMux
    port map (
            O => \N__37990\,
            I => \N__37982\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__37985\,
            I => \N__37977\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__37982\,
            I => \N__37977\
        );

    \I__8220\ : Span4Mux_h
    port map (
            O => \N__37977\,
            I => \N__37973\
        );

    \I__8219\ : InMux
    port map (
            O => \N__37976\,
            I => \N__37970\
        );

    \I__8218\ : Odrv4
    port map (
            O => \N__37973\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__37970\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16\
        );

    \I__8216\ : CascadeMux
    port map (
            O => \N__37965\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16_cascade_\
        );

    \I__8215\ : InMux
    port map (
            O => \N__37962\,
            I => \N__37959\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__37959\,
            I => \N__37956\
        );

    \I__8213\ : Odrv12
    port map (
            O => \N__37956\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_2\
        );

    \I__8212\ : InMux
    port map (
            O => \N__37953\,
            I => \N__37950\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__37950\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_6\
        );

    \I__8210\ : InMux
    port map (
            O => \N__37947\,
            I => \N__37942\
        );

    \I__8209\ : InMux
    port map (
            O => \N__37946\,
            I => \N__37939\
        );

    \I__8208\ : InMux
    port map (
            O => \N__37945\,
            I => \N__37936\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__37942\,
            I => \N__37933\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__37939\,
            I => \N__37929\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__37936\,
            I => \N__37926\
        );

    \I__8204\ : Span4Mux_v
    port map (
            O => \N__37933\,
            I => \N__37923\
        );

    \I__8203\ : InMux
    port map (
            O => \N__37932\,
            I => \N__37920\
        );

    \I__8202\ : Span4Mux_h
    port map (
            O => \N__37929\,
            I => \N__37917\
        );

    \I__8201\ : Odrv4
    port map (
            O => \N__37926\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__37923\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__37920\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8198\ : Odrv4
    port map (
            O => \N__37917\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8197\ : InMux
    port map (
            O => \N__37908\,
            I => \N__37905\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__37905\,
            I => \N__37901\
        );

    \I__8195\ : InMux
    port map (
            O => \N__37904\,
            I => \N__37898\
        );

    \I__8194\ : Span4Mux_v
    port map (
            O => \N__37901\,
            I => \N__37895\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__37898\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__8192\ : Odrv4
    port map (
            O => \N__37895\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__8191\ : CascadeMux
    port map (
            O => \N__37890\,
            I => \N__37886\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__37889\,
            I => \N__37883\
        );

    \I__8189\ : InMux
    port map (
            O => \N__37886\,
            I => \N__37877\
        );

    \I__8188\ : InMux
    port map (
            O => \N__37883\,
            I => \N__37877\
        );

    \I__8187\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37874\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__37877\,
            I => \N__37871\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__37874\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__37871\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__8183\ : InMux
    port map (
            O => \N__37866\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__8182\ : InMux
    port map (
            O => \N__37863\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__8181\ : CEMux
    port map (
            O => \N__37860\,
            I => \N__37845\
        );

    \I__8180\ : CEMux
    port map (
            O => \N__37859\,
            I => \N__37845\
        );

    \I__8179\ : CEMux
    port map (
            O => \N__37858\,
            I => \N__37845\
        );

    \I__8178\ : CEMux
    port map (
            O => \N__37857\,
            I => \N__37845\
        );

    \I__8177\ : CEMux
    port map (
            O => \N__37856\,
            I => \N__37845\
        );

    \I__8176\ : GlobalMux
    port map (
            O => \N__37845\,
            I => \N__37842\
        );

    \I__8175\ : gio2CtrlBuf
    port map (
            O => \N__37842\,
            I => \delay_measurement_inst.delay_hc_timer.N_461_i_g\
        );

    \I__8174\ : InMux
    port map (
            O => \N__37839\,
            I => \N__37835\
        );

    \I__8173\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37832\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__37835\,
            I => \N__37829\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__37832\,
            I => \N__37826\
        );

    \I__8170\ : Span12Mux_v
    port map (
            O => \N__37829\,
            I => \N__37823\
        );

    \I__8169\ : Odrv4
    port map (
            O => \N__37826\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__8168\ : Odrv12
    port map (
            O => \N__37823\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__8167\ : CEMux
    port map (
            O => \N__37818\,
            I => \N__37815\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__37815\,
            I => \N__37812\
        );

    \I__8165\ : Span4Mux_v
    port map (
            O => \N__37812\,
            I => \N__37806\
        );

    \I__8164\ : CEMux
    port map (
            O => \N__37811\,
            I => \N__37803\
        );

    \I__8163\ : CEMux
    port map (
            O => \N__37810\,
            I => \N__37800\
        );

    \I__8162\ : CEMux
    port map (
            O => \N__37809\,
            I => \N__37797\
        );

    \I__8161\ : Span4Mux_h
    port map (
            O => \N__37806\,
            I => \N__37792\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__37803\,
            I => \N__37792\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__37800\,
            I => \N__37787\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__37797\,
            I => \N__37787\
        );

    \I__8157\ : Span4Mux_h
    port map (
            O => \N__37792\,
            I => \N__37784\
        );

    \I__8156\ : Odrv4
    port map (
            O => \N__37787\,
            I => \delay_measurement_inst.delay_hc_timer.N_462_i\
        );

    \I__8155\ : Odrv4
    port map (
            O => \N__37784\,
            I => \delay_measurement_inst.delay_hc_timer.N_462_i\
        );

    \I__8154\ : InMux
    port map (
            O => \N__37779\,
            I => \N__37755\
        );

    \I__8153\ : InMux
    port map (
            O => \N__37778\,
            I => \N__37755\
        );

    \I__8152\ : InMux
    port map (
            O => \N__37777\,
            I => \N__37755\
        );

    \I__8151\ : InMux
    port map (
            O => \N__37776\,
            I => \N__37755\
        );

    \I__8150\ : InMux
    port map (
            O => \N__37775\,
            I => \N__37746\
        );

    \I__8149\ : InMux
    port map (
            O => \N__37774\,
            I => \N__37746\
        );

    \I__8148\ : InMux
    port map (
            O => \N__37773\,
            I => \N__37746\
        );

    \I__8147\ : InMux
    port map (
            O => \N__37772\,
            I => \N__37746\
        );

    \I__8146\ : InMux
    port map (
            O => \N__37771\,
            I => \N__37737\
        );

    \I__8145\ : InMux
    port map (
            O => \N__37770\,
            I => \N__37737\
        );

    \I__8144\ : InMux
    port map (
            O => \N__37769\,
            I => \N__37737\
        );

    \I__8143\ : InMux
    port map (
            O => \N__37768\,
            I => \N__37737\
        );

    \I__8142\ : InMux
    port map (
            O => \N__37767\,
            I => \N__37714\
        );

    \I__8141\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37714\
        );

    \I__8140\ : InMux
    port map (
            O => \N__37765\,
            I => \N__37714\
        );

    \I__8139\ : InMux
    port map (
            O => \N__37764\,
            I => \N__37714\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__37755\,
            I => \N__37709\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__37746\,
            I => \N__37709\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__37737\,
            I => \N__37706\
        );

    \I__8135\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37697\
        );

    \I__8134\ : InMux
    port map (
            O => \N__37735\,
            I => \N__37697\
        );

    \I__8133\ : InMux
    port map (
            O => \N__37734\,
            I => \N__37697\
        );

    \I__8132\ : InMux
    port map (
            O => \N__37733\,
            I => \N__37697\
        );

    \I__8131\ : InMux
    port map (
            O => \N__37732\,
            I => \N__37692\
        );

    \I__8130\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37692\
        );

    \I__8129\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37683\
        );

    \I__8128\ : InMux
    port map (
            O => \N__37729\,
            I => \N__37683\
        );

    \I__8127\ : InMux
    port map (
            O => \N__37728\,
            I => \N__37683\
        );

    \I__8126\ : InMux
    port map (
            O => \N__37727\,
            I => \N__37683\
        );

    \I__8125\ : InMux
    port map (
            O => \N__37726\,
            I => \N__37674\
        );

    \I__8124\ : InMux
    port map (
            O => \N__37725\,
            I => \N__37674\
        );

    \I__8123\ : InMux
    port map (
            O => \N__37724\,
            I => \N__37674\
        );

    \I__8122\ : InMux
    port map (
            O => \N__37723\,
            I => \N__37674\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__37714\,
            I => \N__37669\
        );

    \I__8120\ : Span4Mux_v
    port map (
            O => \N__37709\,
            I => \N__37669\
        );

    \I__8119\ : Span4Mux_h
    port map (
            O => \N__37706\,
            I => \N__37666\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__37697\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__37692\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__37683\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__37674\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8114\ : Odrv4
    port map (
            O => \N__37669\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8113\ : Odrv4
    port map (
            O => \N__37666\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8112\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37650\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__37650\,
            I => \N__37645\
        );

    \I__8110\ : InMux
    port map (
            O => \N__37649\,
            I => \N__37641\
        );

    \I__8109\ : InMux
    port map (
            O => \N__37648\,
            I => \N__37638\
        );

    \I__8108\ : Span4Mux_v
    port map (
            O => \N__37645\,
            I => \N__37635\
        );

    \I__8107\ : InMux
    port map (
            O => \N__37644\,
            I => \N__37632\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__37641\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__37638\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8104\ : Odrv4
    port map (
            O => \N__37635\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__37632\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8102\ : InMux
    port map (
            O => \N__37623\,
            I => \N__37620\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__37620\,
            I => \N__37617\
        );

    \I__8100\ : Span12Mux_v
    port map (
            O => \N__37617\,
            I => \N__37614\
        );

    \I__8099\ : Odrv12
    port map (
            O => \N__37614\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__8098\ : InMux
    port map (
            O => \N__37611\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__8097\ : CascadeMux
    port map (
            O => \N__37608\,
            I => \N__37604\
        );

    \I__8096\ : CascadeMux
    port map (
            O => \N__37607\,
            I => \N__37601\
        );

    \I__8095\ : InMux
    port map (
            O => \N__37604\,
            I => \N__37596\
        );

    \I__8094\ : InMux
    port map (
            O => \N__37601\,
            I => \N__37596\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__37596\,
            I => \N__37592\
        );

    \I__8092\ : InMux
    port map (
            O => \N__37595\,
            I => \N__37589\
        );

    \I__8091\ : Span4Mux_h
    port map (
            O => \N__37592\,
            I => \N__37586\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__37589\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__8089\ : Odrv4
    port map (
            O => \N__37586\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__8088\ : InMux
    port map (
            O => \N__37581\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__8087\ : InMux
    port map (
            O => \N__37578\,
            I => \N__37572\
        );

    \I__8086\ : InMux
    port map (
            O => \N__37577\,
            I => \N__37572\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__37572\,
            I => \N__37568\
        );

    \I__8084\ : InMux
    port map (
            O => \N__37571\,
            I => \N__37565\
        );

    \I__8083\ : Span4Mux_v
    port map (
            O => \N__37568\,
            I => \N__37562\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__37565\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__8081\ : Odrv4
    port map (
            O => \N__37562\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__8080\ : InMux
    port map (
            O => \N__37557\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__8079\ : InMux
    port map (
            O => \N__37554\,
            I => \N__37548\
        );

    \I__8078\ : InMux
    port map (
            O => \N__37553\,
            I => \N__37548\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__37548\,
            I => \N__37544\
        );

    \I__8076\ : InMux
    port map (
            O => \N__37547\,
            I => \N__37541\
        );

    \I__8075\ : Span4Mux_v
    port map (
            O => \N__37544\,
            I => \N__37538\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__37541\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__8073\ : Odrv4
    port map (
            O => \N__37538\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__8072\ : InMux
    port map (
            O => \N__37533\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__8071\ : CascadeMux
    port map (
            O => \N__37530\,
            I => \N__37526\
        );

    \I__8070\ : CascadeMux
    port map (
            O => \N__37529\,
            I => \N__37523\
        );

    \I__8069\ : InMux
    port map (
            O => \N__37526\,
            I => \N__37518\
        );

    \I__8068\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37518\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__37518\,
            I => \N__37514\
        );

    \I__8066\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37511\
        );

    \I__8065\ : Span4Mux_h
    port map (
            O => \N__37514\,
            I => \N__37508\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__37511\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__8063\ : Odrv4
    port map (
            O => \N__37508\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__8062\ : InMux
    port map (
            O => \N__37503\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__8061\ : CascadeMux
    port map (
            O => \N__37500\,
            I => \N__37496\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__37499\,
            I => \N__37493\
        );

    \I__8059\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37488\
        );

    \I__8058\ : InMux
    port map (
            O => \N__37493\,
            I => \N__37488\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__37488\,
            I => \N__37484\
        );

    \I__8056\ : InMux
    port map (
            O => \N__37487\,
            I => \N__37481\
        );

    \I__8055\ : Span4Mux_h
    port map (
            O => \N__37484\,
            I => \N__37478\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__37481\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__8053\ : Odrv4
    port map (
            O => \N__37478\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__8052\ : InMux
    port map (
            O => \N__37473\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__8051\ : InMux
    port map (
            O => \N__37470\,
            I => \N__37466\
        );

    \I__8050\ : InMux
    port map (
            O => \N__37469\,
            I => \N__37463\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__37466\,
            I => \N__37459\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__37463\,
            I => \N__37456\
        );

    \I__8047\ : InMux
    port map (
            O => \N__37462\,
            I => \N__37453\
        );

    \I__8046\ : Span4Mux_h
    port map (
            O => \N__37459\,
            I => \N__37450\
        );

    \I__8045\ : Odrv4
    port map (
            O => \N__37456\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__37453\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8043\ : Odrv4
    port map (
            O => \N__37450\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8042\ : InMux
    port map (
            O => \N__37443\,
            I => \bfn_15_25_0_\
        );

    \I__8041\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37436\
        );

    \I__8040\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37433\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__37436\,
            I => \N__37429\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__37433\,
            I => \N__37426\
        );

    \I__8037\ : InMux
    port map (
            O => \N__37432\,
            I => \N__37423\
        );

    \I__8036\ : Span4Mux_h
    port map (
            O => \N__37429\,
            I => \N__37420\
        );

    \I__8035\ : Odrv4
    port map (
            O => \N__37426\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__37423\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8033\ : Odrv4
    port map (
            O => \N__37420\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8032\ : InMux
    port map (
            O => \N__37413\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__8031\ : InMux
    port map (
            O => \N__37410\,
            I => \N__37407\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__37407\,
            I => \N__37403\
        );

    \I__8029\ : InMux
    port map (
            O => \N__37406\,
            I => \N__37400\
        );

    \I__8028\ : Span4Mux_v
    port map (
            O => \N__37403\,
            I => \N__37397\
        );

    \I__8027\ : LocalMux
    port map (
            O => \N__37400\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__8026\ : Odrv4
    port map (
            O => \N__37397\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__8025\ : CascadeMux
    port map (
            O => \N__37392\,
            I => \N__37388\
        );

    \I__8024\ : CascadeMux
    port map (
            O => \N__37391\,
            I => \N__37385\
        );

    \I__8023\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37379\
        );

    \I__8022\ : InMux
    port map (
            O => \N__37385\,
            I => \N__37379\
        );

    \I__8021\ : InMux
    port map (
            O => \N__37384\,
            I => \N__37376\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__37379\,
            I => \N__37373\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__37376\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__8018\ : Odrv4
    port map (
            O => \N__37373\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__8017\ : InMux
    port map (
            O => \N__37368\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__8016\ : CascadeMux
    port map (
            O => \N__37365\,
            I => \N__37361\
        );

    \I__8015\ : CascadeMux
    port map (
            O => \N__37364\,
            I => \N__37358\
        );

    \I__8014\ : InMux
    port map (
            O => \N__37361\,
            I => \N__37352\
        );

    \I__8013\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37352\
        );

    \I__8012\ : InMux
    port map (
            O => \N__37357\,
            I => \N__37349\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__37352\,
            I => \N__37346\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__37349\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__8009\ : Odrv4
    port map (
            O => \N__37346\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__8008\ : InMux
    port map (
            O => \N__37341\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__8007\ : CascadeMux
    port map (
            O => \N__37338\,
            I => \N__37334\
        );

    \I__8006\ : CascadeMux
    port map (
            O => \N__37337\,
            I => \N__37331\
        );

    \I__8005\ : InMux
    port map (
            O => \N__37334\,
            I => \N__37326\
        );

    \I__8004\ : InMux
    port map (
            O => \N__37331\,
            I => \N__37326\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__37326\,
            I => \N__37322\
        );

    \I__8002\ : InMux
    port map (
            O => \N__37325\,
            I => \N__37319\
        );

    \I__8001\ : Span4Mux_h
    port map (
            O => \N__37322\,
            I => \N__37316\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__37319\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__7999\ : Odrv4
    port map (
            O => \N__37316\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__7998\ : InMux
    port map (
            O => \N__37311\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__7997\ : InMux
    port map (
            O => \N__37308\,
            I => \N__37301\
        );

    \I__7996\ : InMux
    port map (
            O => \N__37307\,
            I => \N__37301\
        );

    \I__7995\ : InMux
    port map (
            O => \N__37306\,
            I => \N__37298\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__37301\,
            I => \N__37295\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__37298\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__7992\ : Odrv4
    port map (
            O => \N__37295\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__7991\ : InMux
    port map (
            O => \N__37290\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__7990\ : InMux
    port map (
            O => \N__37287\,
            I => \N__37281\
        );

    \I__7989\ : InMux
    port map (
            O => \N__37286\,
            I => \N__37281\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__37281\,
            I => \N__37277\
        );

    \I__7987\ : InMux
    port map (
            O => \N__37280\,
            I => \N__37274\
        );

    \I__7986\ : Span4Mux_v
    port map (
            O => \N__37277\,
            I => \N__37271\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__37274\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__7984\ : Odrv4
    port map (
            O => \N__37271\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__7983\ : InMux
    port map (
            O => \N__37266\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__7982\ : CascadeMux
    port map (
            O => \N__37263\,
            I => \N__37259\
        );

    \I__7981\ : CascadeMux
    port map (
            O => \N__37262\,
            I => \N__37256\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37259\,
            I => \N__37251\
        );

    \I__7979\ : InMux
    port map (
            O => \N__37256\,
            I => \N__37251\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__37251\,
            I => \N__37247\
        );

    \I__7977\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37244\
        );

    \I__7976\ : Span4Mux_h
    port map (
            O => \N__37247\,
            I => \N__37241\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__37244\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__7974\ : Odrv4
    port map (
            O => \N__37241\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__7973\ : InMux
    port map (
            O => \N__37236\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__7972\ : CascadeMux
    port map (
            O => \N__37233\,
            I => \N__37229\
        );

    \I__7971\ : CascadeMux
    port map (
            O => \N__37232\,
            I => \N__37226\
        );

    \I__7970\ : InMux
    port map (
            O => \N__37229\,
            I => \N__37221\
        );

    \I__7969\ : InMux
    port map (
            O => \N__37226\,
            I => \N__37221\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__37221\,
            I => \N__37217\
        );

    \I__7967\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37214\
        );

    \I__7966\ : Span4Mux_h
    port map (
            O => \N__37217\,
            I => \N__37211\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__37214\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__7964\ : Odrv4
    port map (
            O => \N__37211\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__7963\ : InMux
    port map (
            O => \N__37206\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__7962\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37199\
        );

    \I__7961\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37196\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__37199\,
            I => \N__37192\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__37196\,
            I => \N__37189\
        );

    \I__7958\ : InMux
    port map (
            O => \N__37195\,
            I => \N__37186\
        );

    \I__7957\ : Span4Mux_h
    port map (
            O => \N__37192\,
            I => \N__37183\
        );

    \I__7956\ : Odrv4
    port map (
            O => \N__37189\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__37186\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__7954\ : Odrv4
    port map (
            O => \N__37183\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__7953\ : InMux
    port map (
            O => \N__37176\,
            I => \bfn_15_24_0_\
        );

    \I__7952\ : InMux
    port map (
            O => \N__37173\,
            I => \N__37169\
        );

    \I__7951\ : InMux
    port map (
            O => \N__37172\,
            I => \N__37166\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__37169\,
            I => \N__37162\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__37166\,
            I => \N__37159\
        );

    \I__7948\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37156\
        );

    \I__7947\ : Span4Mux_h
    port map (
            O => \N__37162\,
            I => \N__37153\
        );

    \I__7946\ : Odrv4
    port map (
            O => \N__37159\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__37156\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__7944\ : Odrv4
    port map (
            O => \N__37153\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__7943\ : InMux
    port map (
            O => \N__37146\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__7942\ : CascadeMux
    port map (
            O => \N__37143\,
            I => \N__37139\
        );

    \I__7941\ : CascadeMux
    port map (
            O => \N__37142\,
            I => \N__37136\
        );

    \I__7940\ : InMux
    port map (
            O => \N__37139\,
            I => \N__37130\
        );

    \I__7939\ : InMux
    port map (
            O => \N__37136\,
            I => \N__37130\
        );

    \I__7938\ : InMux
    port map (
            O => \N__37135\,
            I => \N__37127\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__37130\,
            I => \N__37124\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__37127\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__7935\ : Odrv4
    port map (
            O => \N__37124\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__7934\ : CascadeMux
    port map (
            O => \N__37119\,
            I => \N__37115\
        );

    \I__7933\ : CascadeMux
    port map (
            O => \N__37118\,
            I => \N__37112\
        );

    \I__7932\ : InMux
    port map (
            O => \N__37115\,
            I => \N__37106\
        );

    \I__7931\ : InMux
    port map (
            O => \N__37112\,
            I => \N__37106\
        );

    \I__7930\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37103\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__37106\,
            I => \N__37100\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__37103\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__7927\ : Odrv4
    port map (
            O => \N__37100\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__7926\ : InMux
    port map (
            O => \N__37095\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__7925\ : CascadeMux
    port map (
            O => \N__37092\,
            I => \N__37088\
        );

    \I__7924\ : CascadeMux
    port map (
            O => \N__37091\,
            I => \N__37085\
        );

    \I__7923\ : InMux
    port map (
            O => \N__37088\,
            I => \N__37080\
        );

    \I__7922\ : InMux
    port map (
            O => \N__37085\,
            I => \N__37080\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__37080\,
            I => \N__37076\
        );

    \I__7920\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37073\
        );

    \I__7919\ : Span4Mux_h
    port map (
            O => \N__37076\,
            I => \N__37070\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__37073\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__7917\ : Odrv4
    port map (
            O => \N__37070\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__7916\ : InMux
    port map (
            O => \N__37065\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__7915\ : InMux
    port map (
            O => \N__37062\,
            I => \N__37056\
        );

    \I__7914\ : InMux
    port map (
            O => \N__37061\,
            I => \N__37056\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__37056\,
            I => \N__37052\
        );

    \I__7912\ : InMux
    port map (
            O => \N__37055\,
            I => \N__37049\
        );

    \I__7911\ : Span4Mux_v
    port map (
            O => \N__37052\,
            I => \N__37046\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__37049\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__37046\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__7908\ : InMux
    port map (
            O => \N__37041\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__7907\ : InMux
    port map (
            O => \N__37038\,
            I => \N__37032\
        );

    \I__7906\ : InMux
    port map (
            O => \N__37037\,
            I => \N__37032\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__37032\,
            I => \N__37028\
        );

    \I__7904\ : InMux
    port map (
            O => \N__37031\,
            I => \N__37025\
        );

    \I__7903\ : Span4Mux_v
    port map (
            O => \N__37028\,
            I => \N__37022\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__37025\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__7901\ : Odrv4
    port map (
            O => \N__37022\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__7900\ : InMux
    port map (
            O => \N__37017\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__7899\ : CascadeMux
    port map (
            O => \N__37014\,
            I => \N__37010\
        );

    \I__7898\ : CascadeMux
    port map (
            O => \N__37013\,
            I => \N__37007\
        );

    \I__7897\ : InMux
    port map (
            O => \N__37010\,
            I => \N__37002\
        );

    \I__7896\ : InMux
    port map (
            O => \N__37007\,
            I => \N__37002\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__37002\,
            I => \N__36998\
        );

    \I__7894\ : InMux
    port map (
            O => \N__37001\,
            I => \N__36995\
        );

    \I__7893\ : Span4Mux_h
    port map (
            O => \N__36998\,
            I => \N__36992\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__36995\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__7891\ : Odrv4
    port map (
            O => \N__36992\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__7890\ : InMux
    port map (
            O => \N__36987\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__7889\ : CascadeMux
    port map (
            O => \N__36984\,
            I => \N__36980\
        );

    \I__7888\ : CascadeMux
    port map (
            O => \N__36983\,
            I => \N__36977\
        );

    \I__7887\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36972\
        );

    \I__7886\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36972\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__36972\,
            I => \N__36968\
        );

    \I__7884\ : InMux
    port map (
            O => \N__36971\,
            I => \N__36965\
        );

    \I__7883\ : Span4Mux_h
    port map (
            O => \N__36968\,
            I => \N__36962\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__36965\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__7881\ : Odrv4
    port map (
            O => \N__36962\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__7880\ : InMux
    port map (
            O => \N__36957\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__7879\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36950\
        );

    \I__7878\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36947\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__36950\,
            I => \N__36944\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__36947\,
            I => \N__36940\
        );

    \I__7875\ : Span4Mux_h
    port map (
            O => \N__36944\,
            I => \N__36937\
        );

    \I__7874\ : InMux
    port map (
            O => \N__36943\,
            I => \N__36934\
        );

    \I__7873\ : Span4Mux_h
    port map (
            O => \N__36940\,
            I => \N__36931\
        );

    \I__7872\ : Odrv4
    port map (
            O => \N__36937\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__36934\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__7870\ : Odrv4
    port map (
            O => \N__36931\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__7869\ : InMux
    port map (
            O => \N__36924\,
            I => \bfn_15_23_0_\
        );

    \I__7868\ : InMux
    port map (
            O => \N__36921\,
            I => \N__36917\
        );

    \I__7867\ : InMux
    port map (
            O => \N__36920\,
            I => \N__36914\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__36917\,
            I => \N__36910\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__36914\,
            I => \N__36907\
        );

    \I__7864\ : InMux
    port map (
            O => \N__36913\,
            I => \N__36904\
        );

    \I__7863\ : Span4Mux_h
    port map (
            O => \N__36910\,
            I => \N__36901\
        );

    \I__7862\ : Odrv4
    port map (
            O => \N__36907\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__36904\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__36901\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__7859\ : InMux
    port map (
            O => \N__36894\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__7858\ : InMux
    port map (
            O => \N__36891\,
            I => \N__36888\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__36888\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\
        );

    \I__7856\ : InMux
    port map (
            O => \N__36885\,
            I => \N__36881\
        );

    \I__7855\ : InMux
    port map (
            O => \N__36884\,
            I => \N__36878\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__36881\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__36878\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__7852\ : InMux
    port map (
            O => \N__36873\,
            I => \N__36870\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__36870\,
            I => \N__36867\
        );

    \I__7850\ : Odrv4
    port map (
            O => \N__36867\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\
        );

    \I__7849\ : InMux
    port map (
            O => \N__36864\,
            I => \N__36861\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__36861\,
            I => \N__36857\
        );

    \I__7847\ : InMux
    port map (
            O => \N__36860\,
            I => \N__36854\
        );

    \I__7846\ : Odrv4
    port map (
            O => \N__36857\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__36854\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7844\ : InMux
    port map (
            O => \N__36849\,
            I => \N__36846\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__36846\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\
        );

    \I__7842\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36839\
        );

    \I__7841\ : InMux
    port map (
            O => \N__36842\,
            I => \N__36836\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__36839\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__36836\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7838\ : CascadeMux
    port map (
            O => \N__36831\,
            I => \N__36828\
        );

    \I__7837\ : InMux
    port map (
            O => \N__36828\,
            I => \N__36825\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__36825\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__7835\ : CascadeMux
    port map (
            O => \N__36822\,
            I => \N__36819\
        );

    \I__7834\ : InMux
    port map (
            O => \N__36819\,
            I => \N__36816\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__36816\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__7832\ : CascadeMux
    port map (
            O => \N__36813\,
            I => \N__36810\
        );

    \I__7831\ : InMux
    port map (
            O => \N__36810\,
            I => \N__36807\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__36807\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__7829\ : CascadeMux
    port map (
            O => \N__36804\,
            I => \N__36801\
        );

    \I__7828\ : InMux
    port map (
            O => \N__36801\,
            I => \N__36798\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__36798\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__7826\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36791\
        );

    \I__7825\ : InMux
    port map (
            O => \N__36794\,
            I => \N__36787\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__36791\,
            I => \N__36784\
        );

    \I__7823\ : InMux
    port map (
            O => \N__36790\,
            I => \N__36781\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__36787\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__7821\ : Odrv4
    port map (
            O => \N__36784\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__36781\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__7819\ : InMux
    port map (
            O => \N__36774\,
            I => \N__36770\
        );

    \I__7818\ : InMux
    port map (
            O => \N__36773\,
            I => \N__36766\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__36770\,
            I => \N__36763\
        );

    \I__7816\ : InMux
    port map (
            O => \N__36769\,
            I => \N__36760\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__36766\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__7814\ : Odrv4
    port map (
            O => \N__36763\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__36760\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__7812\ : InMux
    port map (
            O => \N__36753\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__7811\ : InMux
    port map (
            O => \N__36750\,
            I => \N__36746\
        );

    \I__7810\ : InMux
    port map (
            O => \N__36749\,
            I => \N__36743\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__36746\,
            I => \N__36740\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__36743\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7807\ : Odrv4
    port map (
            O => \N__36740\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7806\ : InMux
    port map (
            O => \N__36735\,
            I => \N__36732\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__36732\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\
        );

    \I__7804\ : InMux
    port map (
            O => \N__36729\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__7803\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36722\
        );

    \I__7802\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36719\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__36722\,
            I => \N__36716\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__36719\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__7799\ : Odrv4
    port map (
            O => \N__36716\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__7798\ : InMux
    port map (
            O => \N__36711\,
            I => \N__36708\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__36708\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\
        );

    \I__7796\ : InMux
    port map (
            O => \N__36705\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__7795\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36698\
        );

    \I__7794\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36695\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__36698\,
            I => \N__36692\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__36695\,
            I => \N__36687\
        );

    \I__7791\ : Span4Mux_v
    port map (
            O => \N__36692\,
            I => \N__36687\
        );

    \I__7790\ : Odrv4
    port map (
            O => \N__36687\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__7789\ : InMux
    port map (
            O => \N__36684\,
            I => \N__36681\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__36681\,
            I => \N__36678\
        );

    \I__7787\ : Odrv12
    port map (
            O => \N__36678\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\
        );

    \I__7786\ : InMux
    port map (
            O => \N__36675\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__7785\ : InMux
    port map (
            O => \N__36672\,
            I => \bfn_15_19_0_\
        );

    \I__7784\ : InMux
    port map (
            O => \N__36669\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__7783\ : InMux
    port map (
            O => \N__36666\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__7782\ : InMux
    port map (
            O => \N__36663\,
            I => \N__36660\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__36660\,
            I => \N__36657\
        );

    \I__7780\ : Odrv4
    port map (
            O => \N__36657\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__7779\ : InMux
    port map (
            O => \N__36654\,
            I => \N__36651\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__36651\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\
        );

    \I__7777\ : InMux
    port map (
            O => \N__36648\,
            I => \N__36644\
        );

    \I__7776\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36641\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__36644\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__36641\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7773\ : InMux
    port map (
            O => \N__36636\,
            I => \N__36633\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__36633\,
            I => \N__36630\
        );

    \I__7771\ : Span4Mux_h
    port map (
            O => \N__36630\,
            I => \N__36626\
        );

    \I__7770\ : InMux
    port map (
            O => \N__36629\,
            I => \N__36623\
        );

    \I__7769\ : Odrv4
    port map (
            O => \N__36626\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__36623\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7767\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36615\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__36615\,
            I => \N__36612\
        );

    \I__7765\ : Span4Mux_h
    port map (
            O => \N__36612\,
            I => \N__36609\
        );

    \I__7764\ : Odrv4
    port map (
            O => \N__36609\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\
        );

    \I__7763\ : InMux
    port map (
            O => \N__36606\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__7762\ : InMux
    port map (
            O => \N__36603\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__7761\ : InMux
    port map (
            O => \N__36600\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__7760\ : InMux
    port map (
            O => \N__36597\,
            I => \bfn_15_18_0_\
        );

    \I__7759\ : InMux
    port map (
            O => \N__36594\,
            I => \N__36590\
        );

    \I__7758\ : InMux
    port map (
            O => \N__36593\,
            I => \N__36587\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__36590\,
            I => \N__36584\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__36587\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7755\ : Odrv4
    port map (
            O => \N__36584\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7754\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36576\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__36576\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\
        );

    \I__7752\ : InMux
    port map (
            O => \N__36573\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__7751\ : InMux
    port map (
            O => \N__36570\,
            I => \N__36566\
        );

    \I__7750\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36563\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__36566\,
            I => \N__36560\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__36563\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7747\ : Odrv4
    port map (
            O => \N__36560\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7746\ : InMux
    port map (
            O => \N__36555\,
            I => \N__36552\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__36552\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\
        );

    \I__7744\ : InMux
    port map (
            O => \N__36549\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__7743\ : InMux
    port map (
            O => \N__36546\,
            I => \N__36542\
        );

    \I__7742\ : InMux
    port map (
            O => \N__36545\,
            I => \N__36539\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__36542\,
            I => \N__36536\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__36539\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7739\ : Odrv4
    port map (
            O => \N__36536\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7738\ : InMux
    port map (
            O => \N__36531\,
            I => \N__36528\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__36528\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\
        );

    \I__7736\ : InMux
    port map (
            O => \N__36525\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__7735\ : InMux
    port map (
            O => \N__36522\,
            I => \N__36519\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__36519\,
            I => \N__36516\
        );

    \I__7733\ : Span4Mux_v
    port map (
            O => \N__36516\,
            I => \N__36512\
        );

    \I__7732\ : InMux
    port map (
            O => \N__36515\,
            I => \N__36509\
        );

    \I__7731\ : Odrv4
    port map (
            O => \N__36512\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__36509\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7729\ : InMux
    port map (
            O => \N__36504\,
            I => \N__36501\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__36501\,
            I => \N__36498\
        );

    \I__7727\ : Span4Mux_v
    port map (
            O => \N__36498\,
            I => \N__36495\
        );

    \I__7726\ : Odrv4
    port map (
            O => \N__36495\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\
        );

    \I__7725\ : InMux
    port map (
            O => \N__36492\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__7724\ : CascadeMux
    port map (
            O => \N__36489\,
            I => \N__36485\
        );

    \I__7723\ : CascadeMux
    port map (
            O => \N__36488\,
            I => \N__36482\
        );

    \I__7722\ : InMux
    port map (
            O => \N__36485\,
            I => \N__36479\
        );

    \I__7721\ : InMux
    port map (
            O => \N__36482\,
            I => \N__36476\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36472\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__36476\,
            I => \N__36469\
        );

    \I__7718\ : CascadeMux
    port map (
            O => \N__36475\,
            I => \N__36466\
        );

    \I__7717\ : Span4Mux_h
    port map (
            O => \N__36472\,
            I => \N__36463\
        );

    \I__7716\ : Span4Mux_h
    port map (
            O => \N__36469\,
            I => \N__36460\
        );

    \I__7715\ : InMux
    port map (
            O => \N__36466\,
            I => \N__36457\
        );

    \I__7714\ : Span4Mux_v
    port map (
            O => \N__36463\,
            I => \N__36454\
        );

    \I__7713\ : Span4Mux_v
    port map (
            O => \N__36460\,
            I => \N__36451\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__36457\,
            I => \N__36448\
        );

    \I__7711\ : Odrv4
    port map (
            O => \N__36454\,
            I => measured_delay_tr_1
        );

    \I__7710\ : Odrv4
    port map (
            O => \N__36451\,
            I => measured_delay_tr_1
        );

    \I__7709\ : Odrv4
    port map (
            O => \N__36448\,
            I => measured_delay_tr_1
        );

    \I__7708\ : InMux
    port map (
            O => \N__36441\,
            I => \N__36435\
        );

    \I__7707\ : InMux
    port map (
            O => \N__36440\,
            I => \N__36435\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__36435\,
            I => \N__36427\
        );

    \I__7705\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36416\
        );

    \I__7704\ : InMux
    port map (
            O => \N__36433\,
            I => \N__36416\
        );

    \I__7703\ : InMux
    port map (
            O => \N__36432\,
            I => \N__36416\
        );

    \I__7702\ : InMux
    port map (
            O => \N__36431\,
            I => \N__36416\
        );

    \I__7701\ : InMux
    port map (
            O => \N__36430\,
            I => \N__36416\
        );

    \I__7700\ : Span4Mux_v
    port map (
            O => \N__36427\,
            I => \N__36410\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__36416\,
            I => \N__36410\
        );

    \I__7698\ : InMux
    port map (
            O => \N__36415\,
            I => \N__36407\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__36410\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__36407\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i\
        );

    \I__7695\ : CascadeMux
    port map (
            O => \N__36402\,
            I => \N__36399\
        );

    \I__7694\ : InMux
    port map (
            O => \N__36399\,
            I => \N__36392\
        );

    \I__7693\ : InMux
    port map (
            O => \N__36398\,
            I => \N__36392\
        );

    \I__7692\ : CascadeMux
    port map (
            O => \N__36397\,
            I => \N__36389\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__36392\,
            I => \N__36384\
        );

    \I__7690\ : InMux
    port map (
            O => \N__36389\,
            I => \N__36377\
        );

    \I__7689\ : InMux
    port map (
            O => \N__36388\,
            I => \N__36377\
        );

    \I__7688\ : InMux
    port map (
            O => \N__36387\,
            I => \N__36377\
        );

    \I__7687\ : Odrv12
    port map (
            O => \N__36384\,
            I => \delay_measurement_inst.delay_tr_reg_5_tz_1\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__36377\,
            I => \delay_measurement_inst.delay_tr_reg_5_tz_1\
        );

    \I__7685\ : InMux
    port map (
            O => \N__36372\,
            I => \N__36369\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__36369\,
            I => \N__36364\
        );

    \I__7683\ : InMux
    port map (
            O => \N__36368\,
            I => \N__36361\
        );

    \I__7682\ : InMux
    port map (
            O => \N__36367\,
            I => \N__36358\
        );

    \I__7681\ : Span4Mux_v
    port map (
            O => \N__36364\,
            I => \N__36353\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__36361\,
            I => \N__36353\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__36358\,
            I => \N__36350\
        );

    \I__7678\ : Span4Mux_v
    port map (
            O => \N__36353\,
            I => \N__36344\
        );

    \I__7677\ : Span4Mux_v
    port map (
            O => \N__36350\,
            I => \N__36344\
        );

    \I__7676\ : InMux
    port map (
            O => \N__36349\,
            I => \N__36341\
        );

    \I__7675\ : Span4Mux_h
    port map (
            O => \N__36344\,
            I => \N__36338\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__36341\,
            I => measured_delay_tr_2
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__36338\,
            I => measured_delay_tr_2
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__36333\,
            I => \N__36329\
        );

    \I__7671\ : InMux
    port map (
            O => \N__36332\,
            I => \N__36325\
        );

    \I__7670\ : InMux
    port map (
            O => \N__36329\,
            I => \N__36322\
        );

    \I__7669\ : InMux
    port map (
            O => \N__36328\,
            I => \N__36319\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__36325\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__36322\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__36319\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7665\ : InMux
    port map (
            O => \N__36312\,
            I => \N__36309\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__36309\,
            I => \N__36306\
        );

    \I__7663\ : Span4Mux_v
    port map (
            O => \N__36306\,
            I => \N__36302\
        );

    \I__7662\ : InMux
    port map (
            O => \N__36305\,
            I => \N__36299\
        );

    \I__7661\ : Odrv4
    port map (
            O => \N__36302\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__36299\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7659\ : InMux
    port map (
            O => \N__36294\,
            I => \N__36291\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__36291\,
            I => \N__36288\
        );

    \I__7657\ : Span4Mux_v
    port map (
            O => \N__36288\,
            I => \N__36285\
        );

    \I__7656\ : Odrv4
    port map (
            O => \N__36285\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\
        );

    \I__7655\ : InMux
    port map (
            O => \N__36282\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__7654\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36276\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__36276\,
            I => \N__36273\
        );

    \I__7652\ : Span4Mux_h
    port map (
            O => \N__36273\,
            I => \N__36269\
        );

    \I__7651\ : InMux
    port map (
            O => \N__36272\,
            I => \N__36266\
        );

    \I__7650\ : Odrv4
    port map (
            O => \N__36269\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__36266\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7648\ : CascadeMux
    port map (
            O => \N__36261\,
            I => \N__36258\
        );

    \I__7647\ : InMux
    port map (
            O => \N__36258\,
            I => \N__36255\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__36255\,
            I => \N__36252\
        );

    \I__7645\ : Span4Mux_h
    port map (
            O => \N__36252\,
            I => \N__36249\
        );

    \I__7644\ : Odrv4
    port map (
            O => \N__36249\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\
        );

    \I__7643\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36243\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__36243\,
            I => \N__36240\
        );

    \I__7641\ : Span12Mux_h
    port map (
            O => \N__36240\,
            I => \N__36237\
        );

    \I__7640\ : Odrv12
    port map (
            O => \N__36237\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\
        );

    \I__7639\ : InMux
    port map (
            O => \N__36234\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__7638\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36228\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__36228\,
            I => \N__36225\
        );

    \I__7636\ : Span4Mux_h
    port map (
            O => \N__36225\,
            I => \N__36221\
        );

    \I__7635\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36218\
        );

    \I__7634\ : Odrv4
    port map (
            O => \N__36221\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__36218\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7632\ : InMux
    port map (
            O => \N__36213\,
            I => \N__36210\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__36210\,
            I => \N__36207\
        );

    \I__7630\ : Span4Mux_v
    port map (
            O => \N__36207\,
            I => \N__36204\
        );

    \I__7629\ : Odrv4
    port map (
            O => \N__36204\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\
        );

    \I__7628\ : InMux
    port map (
            O => \N__36201\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__7627\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36195\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__36195\,
            I => \N__36192\
        );

    \I__7625\ : Span4Mux_h
    port map (
            O => \N__36192\,
            I => \N__36188\
        );

    \I__7624\ : InMux
    port map (
            O => \N__36191\,
            I => \N__36185\
        );

    \I__7623\ : Odrv4
    port map (
            O => \N__36188\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__36185\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7621\ : InMux
    port map (
            O => \N__36180\,
            I => \N__36177\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__36177\,
            I => \N__36174\
        );

    \I__7619\ : Span4Mux_h
    port map (
            O => \N__36174\,
            I => \N__36171\
        );

    \I__7618\ : Odrv4
    port map (
            O => \N__36171\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\
        );

    \I__7617\ : InMux
    port map (
            O => \N__36168\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__7616\ : InMux
    port map (
            O => \N__36165\,
            I => \N__36162\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__36162\,
            I => \N__36159\
        );

    \I__7614\ : Span4Mux_h
    port map (
            O => \N__36159\,
            I => \N__36156\
        );

    \I__7613\ : Odrv4
    port map (
            O => \N__36156\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__7612\ : CascadeMux
    port map (
            O => \N__36153\,
            I => \phase_controller_inst1.start_timer_hc_RNOZ0Z_0_cascade_\
        );

    \I__7611\ : InMux
    port map (
            O => \N__36150\,
            I => \N__36145\
        );

    \I__7610\ : InMux
    port map (
            O => \N__36149\,
            I => \N__36142\
        );

    \I__7609\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36139\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__36145\,
            I => \N__36136\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__36142\,
            I => \N__36131\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__36139\,
            I => \N__36131\
        );

    \I__7605\ : Span4Mux_h
    port map (
            O => \N__36136\,
            I => \N__36126\
        );

    \I__7604\ : Span4Mux_v
    port map (
            O => \N__36131\,
            I => \N__36126\
        );

    \I__7603\ : Span4Mux_v
    port map (
            O => \N__36126\,
            I => \N__36123\
        );

    \I__7602\ : Span4Mux_v
    port map (
            O => \N__36123\,
            I => \N__36120\
        );

    \I__7601\ : Odrv4
    port map (
            O => \N__36120\,
            I => \il_max_comp1_D2\
        );

    \I__7600\ : InMux
    port map (
            O => \N__36117\,
            I => \N__36112\
        );

    \I__7599\ : InMux
    port map (
            O => \N__36116\,
            I => \N__36107\
        );

    \I__7598\ : CascadeMux
    port map (
            O => \N__36115\,
            I => \N__36104\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__36112\,
            I => \N__36101\
        );

    \I__7596\ : InMux
    port map (
            O => \N__36111\,
            I => \N__36096\
        );

    \I__7595\ : InMux
    port map (
            O => \N__36110\,
            I => \N__36096\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__36107\,
            I => \N__36092\
        );

    \I__7593\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36089\
        );

    \I__7592\ : Span4Mux_h
    port map (
            O => \N__36101\,
            I => \N__36086\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__36096\,
            I => \N__36083\
        );

    \I__7590\ : InMux
    port map (
            O => \N__36095\,
            I => \N__36080\
        );

    \I__7589\ : Odrv4
    port map (
            O => \N__36092\,
            I => state_3
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__36089\,
            I => state_3
        );

    \I__7587\ : Odrv4
    port map (
            O => \N__36086\,
            I => state_3
        );

    \I__7586\ : Odrv4
    port map (
            O => \N__36083\,
            I => state_3
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__36080\,
            I => state_3
        );

    \I__7584\ : InMux
    port map (
            O => \N__36069\,
            I => \N__36066\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__36066\,
            I => \N__36061\
        );

    \I__7582\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36058\
        );

    \I__7581\ : InMux
    port map (
            O => \N__36064\,
            I => \N__36055\
        );

    \I__7580\ : Odrv4
    port map (
            O => \N__36061\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__36058\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__36055\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__7577\ : CascadeMux
    port map (
            O => \N__36048\,
            I => \N__36045\
        );

    \I__7576\ : InMux
    port map (
            O => \N__36045\,
            I => \N__36041\
        );

    \I__7575\ : CascadeMux
    port map (
            O => \N__36044\,
            I => \N__36037\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__36041\,
            I => \N__36033\
        );

    \I__7573\ : InMux
    port map (
            O => \N__36040\,
            I => \N__36026\
        );

    \I__7572\ : InMux
    port map (
            O => \N__36037\,
            I => \N__36026\
        );

    \I__7571\ : InMux
    port map (
            O => \N__36036\,
            I => \N__36026\
        );

    \I__7570\ : Odrv12
    port map (
            O => \N__36033\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__36026\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__7568\ : IoInMux
    port map (
            O => \N__36021\,
            I => \N__36018\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__36018\,
            I => \N__36015\
        );

    \I__7566\ : IoSpan4Mux
    port map (
            O => \N__36015\,
            I => \N__36012\
        );

    \I__7565\ : Span4Mux_s2_v
    port map (
            O => \N__36012\,
            I => \N__36009\
        );

    \I__7564\ : Sp12to4
    port map (
            O => \N__36009\,
            I => \N__36006\
        );

    \I__7563\ : Span12Mux_v
    port map (
            O => \N__36006\,
            I => \N__36003\
        );

    \I__7562\ : Odrv12
    port map (
            O => \N__36003\,
            I => s2_phy_c
        );

    \I__7561\ : CascadeMux
    port map (
            O => \N__36000\,
            I => \delay_measurement_inst.N_384_cascade_\
        );

    \I__7560\ : InMux
    port map (
            O => \N__35997\,
            I => \N__35993\
        );

    \I__7559\ : CascadeMux
    port map (
            O => \N__35996\,
            I => \N__35990\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__35993\,
            I => \N__35986\
        );

    \I__7557\ : InMux
    port map (
            O => \N__35990\,
            I => \N__35983\
        );

    \I__7556\ : InMux
    port map (
            O => \N__35989\,
            I => \N__35979\
        );

    \I__7555\ : Span4Mux_v
    port map (
            O => \N__35986\,
            I => \N__35974\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__35983\,
            I => \N__35974\
        );

    \I__7553\ : CascadeMux
    port map (
            O => \N__35982\,
            I => \N__35971\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__35979\,
            I => \N__35968\
        );

    \I__7551\ : Span4Mux_v
    port map (
            O => \N__35974\,
            I => \N__35965\
        );

    \I__7550\ : InMux
    port map (
            O => \N__35971\,
            I => \N__35962\
        );

    \I__7549\ : Span12Mux_v
    port map (
            O => \N__35968\,
            I => \N__35959\
        );

    \I__7548\ : Span4Mux_v
    port map (
            O => \N__35965\,
            I => \N__35956\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__35962\,
            I => measured_delay_tr_4
        );

    \I__7546\ : Odrv12
    port map (
            O => \N__35959\,
            I => measured_delay_tr_4
        );

    \I__7545\ : Odrv4
    port map (
            O => \N__35956\,
            I => measured_delay_tr_4
        );

    \I__7544\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35945\
        );

    \I__7543\ : InMux
    port map (
            O => \N__35948\,
            I => \N__35942\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__35945\,
            I => \N__35938\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__35942\,
            I => \N__35935\
        );

    \I__7540\ : InMux
    port map (
            O => \N__35941\,
            I => \N__35932\
        );

    \I__7539\ : Span4Mux_h
    port map (
            O => \N__35938\,
            I => \N__35927\
        );

    \I__7538\ : Span4Mux_v
    port map (
            O => \N__35935\,
            I => \N__35927\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__35932\,
            I => \N__35923\
        );

    \I__7536\ : Span4Mux_h
    port map (
            O => \N__35927\,
            I => \N__35920\
        );

    \I__7535\ : InMux
    port map (
            O => \N__35926\,
            I => \N__35917\
        );

    \I__7534\ : Span4Mux_h
    port map (
            O => \N__35923\,
            I => \N__35914\
        );

    \I__7533\ : Odrv4
    port map (
            O => \N__35920\,
            I => measured_delay_tr_5
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__35917\,
            I => measured_delay_tr_5
        );

    \I__7531\ : Odrv4
    port map (
            O => \N__35914\,
            I => measured_delay_tr_5
        );

    \I__7530\ : InMux
    port map (
            O => \N__35907\,
            I => \N__35903\
        );

    \I__7529\ : InMux
    port map (
            O => \N__35906\,
            I => \N__35900\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__35903\,
            I => \N__35895\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__35900\,
            I => \N__35892\
        );

    \I__7526\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35889\
        );

    \I__7525\ : CascadeMux
    port map (
            O => \N__35898\,
            I => \N__35886\
        );

    \I__7524\ : Span4Mux_h
    port map (
            O => \N__35895\,
            I => \N__35883\
        );

    \I__7523\ : Span4Mux_h
    port map (
            O => \N__35892\,
            I => \N__35878\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__35889\,
            I => \N__35878\
        );

    \I__7521\ : InMux
    port map (
            O => \N__35886\,
            I => \N__35875\
        );

    \I__7520\ : Span4Mux_h
    port map (
            O => \N__35883\,
            I => \N__35872\
        );

    \I__7519\ : Span4Mux_v
    port map (
            O => \N__35878\,
            I => \N__35869\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__35875\,
            I => measured_delay_tr_7
        );

    \I__7517\ : Odrv4
    port map (
            O => \N__35872\,
            I => measured_delay_tr_7
        );

    \I__7516\ : Odrv4
    port map (
            O => \N__35869\,
            I => measured_delay_tr_7
        );

    \I__7515\ : CascadeMux
    port map (
            O => \N__35862\,
            I => \N__35859\
        );

    \I__7514\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35853\
        );

    \I__7513\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35853\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__35853\,
            I => \N__35849\
        );

    \I__7511\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35846\
        );

    \I__7510\ : Odrv4
    port map (
            O => \N__35849\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__35846\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31\
        );

    \I__7508\ : InMux
    port map (
            O => \N__35841\,
            I => \N__35837\
        );

    \I__7507\ : InMux
    port map (
            O => \N__35840\,
            I => \N__35834\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__35837\,
            I => \N__35830\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__35834\,
            I => \N__35827\
        );

    \I__7504\ : InMux
    port map (
            O => \N__35833\,
            I => \N__35824\
        );

    \I__7503\ : Span4Mux_h
    port map (
            O => \N__35830\,
            I => \N__35820\
        );

    \I__7502\ : Span4Mux_h
    port map (
            O => \N__35827\,
            I => \N__35815\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__35824\,
            I => \N__35815\
        );

    \I__7500\ : InMux
    port map (
            O => \N__35823\,
            I => \N__35812\
        );

    \I__7499\ : Span4Mux_h
    port map (
            O => \N__35820\,
            I => \N__35809\
        );

    \I__7498\ : Span4Mux_v
    port map (
            O => \N__35815\,
            I => \N__35806\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__35812\,
            I => measured_delay_tr_8
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__35809\,
            I => measured_delay_tr_8
        );

    \I__7495\ : Odrv4
    port map (
            O => \N__35806\,
            I => measured_delay_tr_8
        );

    \I__7494\ : CascadeMux
    port map (
            O => \N__35799\,
            I => \N__35796\
        );

    \I__7493\ : InMux
    port map (
            O => \N__35796\,
            I => \N__35792\
        );

    \I__7492\ : CascadeMux
    port map (
            O => \N__35795\,
            I => \N__35789\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__35792\,
            I => \N__35784\
        );

    \I__7490\ : InMux
    port map (
            O => \N__35789\,
            I => \N__35781\
        );

    \I__7489\ : InMux
    port map (
            O => \N__35788\,
            I => \N__35778\
        );

    \I__7488\ : CascadeMux
    port map (
            O => \N__35787\,
            I => \N__35775\
        );

    \I__7487\ : Span4Mux_h
    port map (
            O => \N__35784\,
            I => \N__35772\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__35781\,
            I => \N__35767\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__35778\,
            I => \N__35767\
        );

    \I__7484\ : InMux
    port map (
            O => \N__35775\,
            I => \N__35764\
        );

    \I__7483\ : Span4Mux_v
    port map (
            O => \N__35772\,
            I => \N__35761\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__35767\,
            I => \N__35758\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__35764\,
            I => measured_delay_tr_3
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__35761\,
            I => measured_delay_tr_3
        );

    \I__7479\ : Odrv4
    port map (
            O => \N__35758\,
            I => measured_delay_tr_3
        );

    \I__7478\ : InMux
    port map (
            O => \N__35751\,
            I => \N__35748\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__35748\,
            I => \N__35745\
        );

    \I__7476\ : Odrv4
    port map (
            O => \N__35745\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\
        );

    \I__7475\ : InMux
    port map (
            O => \N__35742\,
            I => \N__35739\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__35739\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5\
        );

    \I__7473\ : CascadeMux
    port map (
            O => \N__35736\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31_cascade_\
        );

    \I__7472\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35730\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__35730\,
            I => \N__35725\
        );

    \I__7470\ : InMux
    port map (
            O => \N__35729\,
            I => \N__35722\
        );

    \I__7469\ : InMux
    port map (
            O => \N__35728\,
            I => \N__35719\
        );

    \I__7468\ : Span4Mux_h
    port map (
            O => \N__35725\,
            I => \N__35716\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__35722\,
            I => \N__35711\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__35719\,
            I => \N__35711\
        );

    \I__7465\ : Odrv4
    port map (
            O => \N__35716\,
            I => measured_delay_tr_6
        );

    \I__7464\ : Odrv12
    port map (
            O => \N__35711\,
            I => measured_delay_tr_6
        );

    \I__7463\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35703\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__35703\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0\
        );

    \I__7461\ : CascadeMux
    port map (
            O => \N__35700\,
            I => \delay_measurement_inst.N_381_cascade_\
        );

    \I__7460\ : InMux
    port map (
            O => \N__35697\,
            I => \N__35694\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__35694\,
            I => \delay_measurement_inst.delay_tr_timer.N_376\
        );

    \I__7458\ : CascadeMux
    port map (
            O => \N__35691\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_\
        );

    \I__7457\ : CascadeMux
    port map (
            O => \N__35688\,
            I => \delay_measurement_inst.N_498_cascade_\
        );

    \I__7456\ : InMux
    port map (
            O => \N__35685\,
            I => \N__35681\
        );

    \I__7455\ : InMux
    port map (
            O => \N__35684\,
            I => \N__35678\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__35681\,
            I => \delay_measurement_inst.N_381\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__35678\,
            I => \delay_measurement_inst.N_381\
        );

    \I__7452\ : InMux
    port map (
            O => \N__35673\,
            I => \N__35668\
        );

    \I__7451\ : InMux
    port map (
            O => \N__35672\,
            I => \N__35663\
        );

    \I__7450\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35663\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__35668\,
            I => \N__35660\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__35663\,
            I => \delay_measurement_inst.N_384\
        );

    \I__7447\ : Odrv4
    port map (
            O => \N__35660\,
            I => \delay_measurement_inst.N_384\
        );

    \I__7446\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35651\
        );

    \I__7445\ : InMux
    port map (
            O => \N__35654\,
            I => \N__35648\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__35651\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__35648\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7442\ : CascadeMux
    port map (
            O => \N__35643\,
            I => \N__35640\
        );

    \I__7441\ : InMux
    port map (
            O => \N__35640\,
            I => \N__35637\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__35637\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\
        );

    \I__7439\ : InMux
    port map (
            O => \N__35634\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__7438\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35627\
        );

    \I__7437\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35624\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__35627\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__35624\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7434\ : InMux
    port map (
            O => \N__35619\,
            I => \N__35616\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__35616\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\
        );

    \I__7432\ : InMux
    port map (
            O => \N__35613\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__7431\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35606\
        );

    \I__7430\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35603\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__35606\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__35603\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7427\ : CascadeMux
    port map (
            O => \N__35598\,
            I => \N__35595\
        );

    \I__7426\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35592\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__35592\,
            I => \N__35589\
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__35589\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\
        );

    \I__7423\ : InMux
    port map (
            O => \N__35586\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__7422\ : InMux
    port map (
            O => \N__35583\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__7421\ : InMux
    port map (
            O => \N__35580\,
            I => \N__35576\
        );

    \I__7420\ : InMux
    port map (
            O => \N__35579\,
            I => \N__35573\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__35576\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__35573\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7417\ : CascadeMux
    port map (
            O => \N__35568\,
            I => \N__35565\
        );

    \I__7416\ : InMux
    port map (
            O => \N__35565\,
            I => \N__35562\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__35562\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\
        );

    \I__7414\ : InMux
    port map (
            O => \N__35559\,
            I => \bfn_15_10_0_\
        );

    \I__7413\ : InMux
    port map (
            O => \N__35556\,
            I => \N__35552\
        );

    \I__7412\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35549\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__35552\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__35549\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__7409\ : InMux
    port map (
            O => \N__35544\,
            I => \N__35541\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__35541\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\
        );

    \I__7407\ : InMux
    port map (
            O => \N__35538\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__7406\ : InMux
    port map (
            O => \N__35535\,
            I => \N__35531\
        );

    \I__7405\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35528\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__35531\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__35528\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__7402\ : InMux
    port map (
            O => \N__35523\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__7401\ : CascadeMux
    port map (
            O => \N__35520\,
            I => \N__35517\
        );

    \I__7400\ : InMux
    port map (
            O => \N__35517\,
            I => \N__35514\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__35514\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\
        );

    \I__7398\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35507\
        );

    \I__7397\ : InMux
    port map (
            O => \N__35510\,
            I => \N__35504\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__35507\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__35504\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7394\ : CascadeMux
    port map (
            O => \N__35499\,
            I => \N__35496\
        );

    \I__7393\ : InMux
    port map (
            O => \N__35496\,
            I => \N__35493\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__35493\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\
        );

    \I__7391\ : InMux
    port map (
            O => \N__35490\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__7390\ : InMux
    port map (
            O => \N__35487\,
            I => \N__35483\
        );

    \I__7389\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35480\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__35483\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__35480\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7386\ : InMux
    port map (
            O => \N__35475\,
            I => \N__35472\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__35472\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\
        );

    \I__7384\ : InMux
    port map (
            O => \N__35469\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__7383\ : InMux
    port map (
            O => \N__35466\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__7382\ : InMux
    port map (
            O => \N__35463\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__7381\ : InMux
    port map (
            O => \N__35460\,
            I => \bfn_15_9_0_\
        );

    \I__7380\ : InMux
    port map (
            O => \N__35457\,
            I => \N__35453\
        );

    \I__7379\ : InMux
    port map (
            O => \N__35456\,
            I => \N__35450\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__35453\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__35450\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7376\ : InMux
    port map (
            O => \N__35445\,
            I => \N__35442\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__35442\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\
        );

    \I__7374\ : InMux
    port map (
            O => \N__35439\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__7373\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35432\
        );

    \I__7372\ : InMux
    port map (
            O => \N__35435\,
            I => \N__35429\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__35432\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__35429\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7369\ : InMux
    port map (
            O => \N__35424\,
            I => \N__35421\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__35421\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\
        );

    \I__7367\ : InMux
    port map (
            O => \N__35418\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__7366\ : InMux
    port map (
            O => \N__35415\,
            I => \N__35411\
        );

    \I__7365\ : InMux
    port map (
            O => \N__35414\,
            I => \N__35408\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__35411\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__35408\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7362\ : InMux
    port map (
            O => \N__35403\,
            I => \N__35400\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__35400\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\
        );

    \I__7360\ : InMux
    port map (
            O => \N__35397\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__7359\ : InMux
    port map (
            O => \N__35394\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__7358\ : InMux
    port map (
            O => \N__35391\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__7357\ : InMux
    port map (
            O => \N__35388\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__7356\ : InMux
    port map (
            O => \N__35385\,
            I => \N__35382\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__35382\,
            I => \il_min_comp1_D1\
        );

    \I__7354\ : CEMux
    port map (
            O => \N__35379\,
            I => \N__35375\
        );

    \I__7353\ : CEMux
    port map (
            O => \N__35378\,
            I => \N__35371\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__35375\,
            I => \N__35366\
        );

    \I__7351\ : CEMux
    port map (
            O => \N__35374\,
            I => \N__35363\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__35371\,
            I => \N__35360\
        );

    \I__7349\ : CEMux
    port map (
            O => \N__35370\,
            I => \N__35357\
        );

    \I__7348\ : CEMux
    port map (
            O => \N__35369\,
            I => \N__35354\
        );

    \I__7347\ : Span4Mux_h
    port map (
            O => \N__35366\,
            I => \N__35351\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__35363\,
            I => \N__35348\
        );

    \I__7345\ : Span4Mux_h
    port map (
            O => \N__35360\,
            I => \N__35341\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__35357\,
            I => \N__35341\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__35354\,
            I => \N__35341\
        );

    \I__7342\ : Span4Mux_h
    port map (
            O => \N__35351\,
            I => \N__35338\
        );

    \I__7341\ : Span4Mux_h
    port map (
            O => \N__35348\,
            I => \N__35335\
        );

    \I__7340\ : Span4Mux_v
    port map (
            O => \N__35341\,
            I => \N__35332\
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__35338\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__7338\ : Odrv4
    port map (
            O => \N__35335\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__7337\ : Odrv4
    port map (
            O => \N__35332\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__7336\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35322\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__35322\,
            I => \N__35319\
        );

    \I__7334\ : Odrv4
    port map (
            O => \N__35319\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__7333\ : CascadeMux
    port map (
            O => \N__35316\,
            I => \N__35312\
        );

    \I__7332\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35308\
        );

    \I__7331\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35305\
        );

    \I__7330\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35302\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__35308\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__35305\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__35302\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7326\ : InMux
    port map (
            O => \N__35295\,
            I => \N__35291\
        );

    \I__7325\ : InMux
    port map (
            O => \N__35294\,
            I => \N__35288\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__35291\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__35288\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7322\ : InMux
    port map (
            O => \N__35283\,
            I => \N__35280\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__35280\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\
        );

    \I__7320\ : InMux
    port map (
            O => \N__35277\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__7319\ : InMux
    port map (
            O => \N__35274\,
            I => \N__35271\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__35271\,
            I => \N__35268\
        );

    \I__7317\ : Odrv4
    port map (
            O => \N__35268\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\
        );

    \I__7316\ : CascadeMux
    port map (
            O => \N__35265\,
            I => \N__35262\
        );

    \I__7315\ : InMux
    port map (
            O => \N__35262\,
            I => \N__35258\
        );

    \I__7314\ : InMux
    port map (
            O => \N__35261\,
            I => \N__35255\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__35258\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__35255\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7311\ : CascadeMux
    port map (
            O => \N__35250\,
            I => \N__35247\
        );

    \I__7310\ : InMux
    port map (
            O => \N__35247\,
            I => \N__35244\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__35244\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\
        );

    \I__7308\ : InMux
    port map (
            O => \N__35241\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__7307\ : InMux
    port map (
            O => \N__35238\,
            I => \N__35234\
        );

    \I__7306\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35231\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__35234\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__35231\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7303\ : InMux
    port map (
            O => \N__35226\,
            I => \N__35223\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__35223\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\
        );

    \I__7301\ : InMux
    port map (
            O => \N__35220\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__7300\ : InMux
    port map (
            O => \N__35217\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__7299\ : InMux
    port map (
            O => \N__35214\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__7298\ : InMux
    port map (
            O => \N__35211\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__7297\ : InMux
    port map (
            O => \N__35208\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__7296\ : InMux
    port map (
            O => \N__35205\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__7295\ : InMux
    port map (
            O => \N__35202\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__7294\ : InMux
    port map (
            O => \N__35199\,
            I => \bfn_14_28_0_\
        );

    \I__7293\ : InMux
    port map (
            O => \N__35196\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__7292\ : InMux
    port map (
            O => \N__35193\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__7291\ : InMux
    port map (
            O => \N__35190\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__7290\ : InMux
    port map (
            O => \N__35187\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__7289\ : InMux
    port map (
            O => \N__35184\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__7288\ : InMux
    port map (
            O => \N__35181\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__7287\ : InMux
    port map (
            O => \N__35178\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__7286\ : InMux
    port map (
            O => \N__35175\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__7285\ : InMux
    port map (
            O => \N__35172\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__7284\ : InMux
    port map (
            O => \N__35169\,
            I => \bfn_14_27_0_\
        );

    \I__7283\ : InMux
    port map (
            O => \N__35166\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__7282\ : InMux
    port map (
            O => \N__35163\,
            I => \bfn_14_25_0_\
        );

    \I__7281\ : InMux
    port map (
            O => \N__35160\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__7280\ : InMux
    port map (
            O => \N__35157\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__7279\ : InMux
    port map (
            O => \N__35154\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__7278\ : InMux
    port map (
            O => \N__35151\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__7277\ : InMux
    port map (
            O => \N__35148\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__7276\ : InMux
    port map (
            O => \N__35145\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__7275\ : InMux
    port map (
            O => \N__35142\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__7274\ : InMux
    port map (
            O => \N__35139\,
            I => \bfn_14_26_0_\
        );

    \I__7273\ : InMux
    port map (
            O => \N__35136\,
            I => \N__35133\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__35133\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__7271\ : InMux
    port map (
            O => \N__35130\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__7270\ : CascadeMux
    port map (
            O => \N__35127\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\
        );

    \I__7269\ : CascadeMux
    port map (
            O => \N__35124\,
            I => \N__35121\
        );

    \I__7268\ : InMux
    port map (
            O => \N__35121\,
            I => \N__35118\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__35118\,
            I => \N__35115\
        );

    \I__7266\ : Odrv4
    port map (
            O => \N__35115\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__7265\ : InMux
    port map (
            O => \N__35112\,
            I => \N__35109\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__35109\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__7263\ : CascadeMux
    port map (
            O => \N__35106\,
            I => \N__35103\
        );

    \I__7262\ : InMux
    port map (
            O => \N__35103\,
            I => \N__35100\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__35100\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__7260\ : InMux
    port map (
            O => \N__35097\,
            I => \N__35094\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__35094\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__7258\ : CascadeMux
    port map (
            O => \N__35091\,
            I => \N__35088\
        );

    \I__7257\ : InMux
    port map (
            O => \N__35088\,
            I => \N__35085\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__35085\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__7255\ : InMux
    port map (
            O => \N__35082\,
            I => \N__35079\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__35079\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__7253\ : InMux
    port map (
            O => \N__35076\,
            I => \N__35073\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__35073\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__7251\ : InMux
    port map (
            O => \N__35070\,
            I => \N__35067\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__35067\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__7249\ : InMux
    port map (
            O => \N__35064\,
            I => \N__35061\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__35061\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__7247\ : InMux
    port map (
            O => \N__35058\,
            I => \N__35055\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__35055\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__7245\ : InMux
    port map (
            O => \N__35052\,
            I => \N__35049\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__35049\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__7243\ : InMux
    port map (
            O => \N__35046\,
            I => \N__35043\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__35043\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__7241\ : CascadeMux
    port map (
            O => \N__35040\,
            I => \N__35037\
        );

    \I__7240\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35034\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__35034\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__7238\ : InMux
    port map (
            O => \N__35031\,
            I => \N__35028\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__35028\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__7236\ : InMux
    port map (
            O => \N__35025\,
            I => \N__35022\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__35022\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__7234\ : InMux
    port map (
            O => \N__35019\,
            I => \N__35016\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__35016\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__7232\ : InMux
    port map (
            O => \N__35013\,
            I => \N__35010\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__35010\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__7230\ : InMux
    port map (
            O => \N__35007\,
            I => \N__35004\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__35004\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__7228\ : CascadeMux
    port map (
            O => \N__35001\,
            I => \N__34998\
        );

    \I__7227\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34995\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__34995\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__7225\ : CascadeMux
    port map (
            O => \N__34992\,
            I => \N__34989\
        );

    \I__7224\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34986\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__34986\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__7222\ : InMux
    port map (
            O => \N__34983\,
            I => \N__34980\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__34980\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__7220\ : CascadeMux
    port map (
            O => \N__34977\,
            I => \N__34974\
        );

    \I__7219\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34971\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__34971\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__7217\ : InMux
    port map (
            O => \N__34968\,
            I => \N__34965\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__34965\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__7215\ : CascadeMux
    port map (
            O => \N__34962\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__7214\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34956\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__34956\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\
        );

    \I__7212\ : CascadeMux
    port map (
            O => \N__34953\,
            I => \N__34950\
        );

    \I__7211\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34947\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__34947\,
            I => \N__34944\
        );

    \I__7209\ : Odrv4
    port map (
            O => \N__34944\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__7208\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34938\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__34938\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__7206\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34932\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__34932\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__7204\ : InMux
    port map (
            O => \N__34929\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__7203\ : CascadeMux
    port map (
            O => \N__34926\,
            I => \N__34923\
        );

    \I__7202\ : InMux
    port map (
            O => \N__34923\,
            I => \N__34919\
        );

    \I__7201\ : InMux
    port map (
            O => \N__34922\,
            I => \N__34916\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__34919\,
            I => \N__34910\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__34916\,
            I => \N__34910\
        );

    \I__7198\ : InMux
    port map (
            O => \N__34915\,
            I => \N__34907\
        );

    \I__7197\ : Span4Mux_v
    port map (
            O => \N__34910\,
            I => \N__34904\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__34907\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__7195\ : Odrv4
    port map (
            O => \N__34904\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__7194\ : InMux
    port map (
            O => \N__34899\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__7193\ : InMux
    port map (
            O => \N__34896\,
            I => \N__34889\
        );

    \I__7192\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34889\
        );

    \I__7191\ : InMux
    port map (
            O => \N__34894\,
            I => \N__34886\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__34889\,
            I => \N__34883\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__34886\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__7188\ : Odrv4
    port map (
            O => \N__34883\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__7187\ : InMux
    port map (
            O => \N__34878\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__7186\ : InMux
    port map (
            O => \N__34875\,
            I => \N__34871\
        );

    \I__7185\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34868\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__34871\,
            I => \N__34865\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__34868\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__7182\ : Odrv4
    port map (
            O => \N__34865\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__7181\ : InMux
    port map (
            O => \N__34860\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__7180\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34821\
        );

    \I__7179\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34821\
        );

    \I__7178\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34821\
        );

    \I__7177\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34821\
        );

    \I__7176\ : InMux
    port map (
            O => \N__34853\,
            I => \N__34812\
        );

    \I__7175\ : InMux
    port map (
            O => \N__34852\,
            I => \N__34812\
        );

    \I__7174\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34812\
        );

    \I__7173\ : InMux
    port map (
            O => \N__34850\,
            I => \N__34812\
        );

    \I__7172\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34803\
        );

    \I__7171\ : InMux
    port map (
            O => \N__34848\,
            I => \N__34803\
        );

    \I__7170\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34803\
        );

    \I__7169\ : InMux
    port map (
            O => \N__34846\,
            I => \N__34803\
        );

    \I__7168\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34794\
        );

    \I__7167\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34794\
        );

    \I__7166\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34794\
        );

    \I__7165\ : InMux
    port map (
            O => \N__34842\,
            I => \N__34794\
        );

    \I__7164\ : InMux
    port map (
            O => \N__34841\,
            I => \N__34785\
        );

    \I__7163\ : InMux
    port map (
            O => \N__34840\,
            I => \N__34785\
        );

    \I__7162\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34785\
        );

    \I__7161\ : InMux
    port map (
            O => \N__34838\,
            I => \N__34785\
        );

    \I__7160\ : InMux
    port map (
            O => \N__34837\,
            I => \N__34776\
        );

    \I__7159\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34776\
        );

    \I__7158\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34776\
        );

    \I__7157\ : InMux
    port map (
            O => \N__34834\,
            I => \N__34776\
        );

    \I__7156\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34765\
        );

    \I__7155\ : InMux
    port map (
            O => \N__34832\,
            I => \N__34765\
        );

    \I__7154\ : InMux
    port map (
            O => \N__34831\,
            I => \N__34765\
        );

    \I__7153\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34765\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__34821\,
            I => \N__34760\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__34812\,
            I => \N__34760\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__34803\,
            I => \N__34751\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__34794\,
            I => \N__34751\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__34785\,
            I => \N__34751\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__34776\,
            I => \N__34751\
        );

    \I__7146\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34746\
        );

    \I__7145\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34746\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__34765\,
            I => \N__34739\
        );

    \I__7143\ : Span4Mux_v
    port map (
            O => \N__34760\,
            I => \N__34739\
        );

    \I__7142\ : Span4Mux_v
    port map (
            O => \N__34751\,
            I => \N__34739\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__34746\,
            I => \N__34736\
        );

    \I__7140\ : Span4Mux_v
    port map (
            O => \N__34739\,
            I => \N__34733\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__34736\,
            I => \N__34730\
        );

    \I__7138\ : Span4Mux_h
    port map (
            O => \N__34733\,
            I => \N__34727\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__34730\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__7136\ : Odrv4
    port map (
            O => \N__34727\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__7135\ : InMux
    port map (
            O => \N__34722\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__7134\ : CascadeMux
    port map (
            O => \N__34719\,
            I => \N__34716\
        );

    \I__7133\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34712\
        );

    \I__7132\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34709\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34706\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__34709\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__7129\ : Odrv4
    port map (
            O => \N__34706\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__7128\ : CEMux
    port map (
            O => \N__34701\,
            I => \N__34697\
        );

    \I__7127\ : CEMux
    port map (
            O => \N__34700\,
            I => \N__34692\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__34697\,
            I => \N__34689\
        );

    \I__7125\ : CEMux
    port map (
            O => \N__34696\,
            I => \N__34686\
        );

    \I__7124\ : CEMux
    port map (
            O => \N__34695\,
            I => \N__34683\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__34692\,
            I => \N__34680\
        );

    \I__7122\ : Span4Mux_v
    port map (
            O => \N__34689\,
            I => \N__34675\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__34686\,
            I => \N__34675\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__34683\,
            I => \N__34672\
        );

    \I__7119\ : Span4Mux_v
    port map (
            O => \N__34680\,
            I => \N__34667\
        );

    \I__7118\ : Span4Mux_h
    port map (
            O => \N__34675\,
            I => \N__34667\
        );

    \I__7117\ : Span4Mux_h
    port map (
            O => \N__34672\,
            I => \N__34664\
        );

    \I__7116\ : Span4Mux_v
    port map (
            O => \N__34667\,
            I => \N__34661\
        );

    \I__7115\ : Span4Mux_h
    port map (
            O => \N__34664\,
            I => \N__34658\
        );

    \I__7114\ : Odrv4
    port map (
            O => \N__34661\,
            I => \current_shift_inst.timer_s1.N_186_i\
        );

    \I__7113\ : Odrv4
    port map (
            O => \N__34658\,
            I => \current_shift_inst.timer_s1.N_186_i\
        );

    \I__7112\ : InMux
    port map (
            O => \N__34653\,
            I => \N__34649\
        );

    \I__7111\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34646\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__34649\,
            I => \N__34643\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__34646\,
            I => \N__34640\
        );

    \I__7108\ : Span4Mux_v
    port map (
            O => \N__34643\,
            I => \N__34637\
        );

    \I__7107\ : Span4Mux_h
    port map (
            O => \N__34640\,
            I => \N__34634\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__34637\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__7105\ : Odrv4
    port map (
            O => \N__34634\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__7104\ : InMux
    port map (
            O => \N__34629\,
            I => \N__34626\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__34626\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__7102\ : CascadeMux
    port map (
            O => \N__34623\,
            I => \N__34620\
        );

    \I__7101\ : InMux
    port map (
            O => \N__34620\,
            I => \N__34615\
        );

    \I__7100\ : InMux
    port map (
            O => \N__34619\,
            I => \N__34610\
        );

    \I__7099\ : InMux
    port map (
            O => \N__34618\,
            I => \N__34610\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__34615\,
            I => \N__34607\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__34610\,
            I => \N__34604\
        );

    \I__7096\ : Span4Mux_h
    port map (
            O => \N__34607\,
            I => \N__34601\
        );

    \I__7095\ : Span4Mux_h
    port map (
            O => \N__34604\,
            I => \N__34598\
        );

    \I__7094\ : Span4Mux_h
    port map (
            O => \N__34601\,
            I => \N__34593\
        );

    \I__7093\ : Span4Mux_h
    port map (
            O => \N__34598\,
            I => \N__34593\
        );

    \I__7092\ : Odrv4
    port map (
            O => \N__34593\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__7091\ : CascadeMux
    port map (
            O => \N__34590\,
            I => \N__34553\
        );

    \I__7090\ : CascadeMux
    port map (
            O => \N__34589\,
            I => \N__34550\
        );

    \I__7089\ : CascadeMux
    port map (
            O => \N__34588\,
            I => \N__34547\
        );

    \I__7088\ : CascadeMux
    port map (
            O => \N__34587\,
            I => \N__34544\
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__34586\,
            I => \N__34541\
        );

    \I__7086\ : CascadeMux
    port map (
            O => \N__34585\,
            I => \N__34538\
        );

    \I__7085\ : CascadeMux
    port map (
            O => \N__34584\,
            I => \N__34535\
        );

    \I__7084\ : CascadeMux
    port map (
            O => \N__34583\,
            I => \N__34532\
        );

    \I__7083\ : CascadeMux
    port map (
            O => \N__34582\,
            I => \N__34529\
        );

    \I__7082\ : CascadeMux
    port map (
            O => \N__34581\,
            I => \N__34526\
        );

    \I__7081\ : CascadeMux
    port map (
            O => \N__34580\,
            I => \N__34523\
        );

    \I__7080\ : CascadeMux
    port map (
            O => \N__34579\,
            I => \N__34520\
        );

    \I__7079\ : CascadeMux
    port map (
            O => \N__34578\,
            I => \N__34517\
        );

    \I__7078\ : CascadeMux
    port map (
            O => \N__34577\,
            I => \N__34514\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__34576\,
            I => \N__34511\
        );

    \I__7076\ : InMux
    port map (
            O => \N__34575\,
            I => \N__34506\
        );

    \I__7075\ : InMux
    port map (
            O => \N__34574\,
            I => \N__34506\
        );

    \I__7074\ : CascadeMux
    port map (
            O => \N__34573\,
            I => \N__34503\
        );

    \I__7073\ : CascadeMux
    port map (
            O => \N__34572\,
            I => \N__34500\
        );

    \I__7072\ : CascadeMux
    port map (
            O => \N__34571\,
            I => \N__34497\
        );

    \I__7071\ : CascadeMux
    port map (
            O => \N__34570\,
            I => \N__34494\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__34569\,
            I => \N__34491\
        );

    \I__7069\ : CascadeMux
    port map (
            O => \N__34568\,
            I => \N__34487\
        );

    \I__7068\ : CascadeMux
    port map (
            O => \N__34567\,
            I => \N__34484\
        );

    \I__7067\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34475\
        );

    \I__7066\ : InMux
    port map (
            O => \N__34565\,
            I => \N__34472\
        );

    \I__7065\ : InMux
    port map (
            O => \N__34564\,
            I => \N__34465\
        );

    \I__7064\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34465\
        );

    \I__7063\ : InMux
    port map (
            O => \N__34562\,
            I => \N__34465\
        );

    \I__7062\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34456\
        );

    \I__7061\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34456\
        );

    \I__7060\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34456\
        );

    \I__7059\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34456\
        );

    \I__7058\ : CascadeMux
    port map (
            O => \N__34557\,
            I => \N__34453\
        );

    \I__7057\ : CascadeMux
    port map (
            O => \N__34556\,
            I => \N__34450\
        );

    \I__7056\ : InMux
    port map (
            O => \N__34553\,
            I => \N__34442\
        );

    \I__7055\ : InMux
    port map (
            O => \N__34550\,
            I => \N__34442\
        );

    \I__7054\ : InMux
    port map (
            O => \N__34547\,
            I => \N__34442\
        );

    \I__7053\ : InMux
    port map (
            O => \N__34544\,
            I => \N__34433\
        );

    \I__7052\ : InMux
    port map (
            O => \N__34541\,
            I => \N__34433\
        );

    \I__7051\ : InMux
    port map (
            O => \N__34538\,
            I => \N__34433\
        );

    \I__7050\ : InMux
    port map (
            O => \N__34535\,
            I => \N__34433\
        );

    \I__7049\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34424\
        );

    \I__7048\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34424\
        );

    \I__7047\ : InMux
    port map (
            O => \N__34526\,
            I => \N__34424\
        );

    \I__7046\ : InMux
    port map (
            O => \N__34523\,
            I => \N__34424\
        );

    \I__7045\ : InMux
    port map (
            O => \N__34520\,
            I => \N__34415\
        );

    \I__7044\ : InMux
    port map (
            O => \N__34517\,
            I => \N__34415\
        );

    \I__7043\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34415\
        );

    \I__7042\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34415\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__34506\,
            I => \N__34412\
        );

    \I__7040\ : InMux
    port map (
            O => \N__34503\,
            I => \N__34405\
        );

    \I__7039\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34405\
        );

    \I__7038\ : InMux
    port map (
            O => \N__34497\,
            I => \N__34405\
        );

    \I__7037\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34394\
        );

    \I__7036\ : InMux
    port map (
            O => \N__34491\,
            I => \N__34394\
        );

    \I__7035\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34394\
        );

    \I__7034\ : InMux
    port map (
            O => \N__34487\,
            I => \N__34394\
        );

    \I__7033\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34394\
        );

    \I__7032\ : CascadeMux
    port map (
            O => \N__34483\,
            I => \N__34391\
        );

    \I__7031\ : CascadeMux
    port map (
            O => \N__34482\,
            I => \N__34388\
        );

    \I__7030\ : CascadeMux
    port map (
            O => \N__34481\,
            I => \N__34385\
        );

    \I__7029\ : CascadeMux
    port map (
            O => \N__34480\,
            I => \N__34382\
        );

    \I__7028\ : CascadeMux
    port map (
            O => \N__34479\,
            I => \N__34379\
        );

    \I__7027\ : CascadeMux
    port map (
            O => \N__34478\,
            I => \N__34376\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__34475\,
            I => \N__34364\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__34472\,
            I => \N__34361\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__34465\,
            I => \N__34356\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__34456\,
            I => \N__34356\
        );

    \I__7022\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34353\
        );

    \I__7021\ : InMux
    port map (
            O => \N__34450\,
            I => \N__34348\
        );

    \I__7020\ : InMux
    port map (
            O => \N__34449\,
            I => \N__34348\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__34442\,
            I => \N__34343\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__34433\,
            I => \N__34343\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__34424\,
            I => \N__34338\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__34415\,
            I => \N__34338\
        );

    \I__7015\ : Span4Mux_h
    port map (
            O => \N__34412\,
            I => \N__34331\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__34405\,
            I => \N__34331\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__34394\,
            I => \N__34331\
        );

    \I__7012\ : InMux
    port map (
            O => \N__34391\,
            I => \N__34324\
        );

    \I__7011\ : InMux
    port map (
            O => \N__34388\,
            I => \N__34324\
        );

    \I__7010\ : InMux
    port map (
            O => \N__34385\,
            I => \N__34324\
        );

    \I__7009\ : InMux
    port map (
            O => \N__34382\,
            I => \N__34315\
        );

    \I__7008\ : InMux
    port map (
            O => \N__34379\,
            I => \N__34315\
        );

    \I__7007\ : InMux
    port map (
            O => \N__34376\,
            I => \N__34315\
        );

    \I__7006\ : InMux
    port map (
            O => \N__34375\,
            I => \N__34315\
        );

    \I__7005\ : InMux
    port map (
            O => \N__34374\,
            I => \N__34312\
        );

    \I__7004\ : InMux
    port map (
            O => \N__34373\,
            I => \N__34305\
        );

    \I__7003\ : InMux
    port map (
            O => \N__34372\,
            I => \N__34305\
        );

    \I__7002\ : InMux
    port map (
            O => \N__34371\,
            I => \N__34305\
        );

    \I__7001\ : InMux
    port map (
            O => \N__34370\,
            I => \N__34296\
        );

    \I__7000\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34296\
        );

    \I__6999\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34296\
        );

    \I__6998\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34296\
        );

    \I__6997\ : Span4Mux_s2_v
    port map (
            O => \N__34364\,
            I => \N__34293\
        );

    \I__6996\ : Span4Mux_v
    port map (
            O => \N__34361\,
            I => \N__34287\
        );

    \I__6995\ : Span4Mux_v
    port map (
            O => \N__34356\,
            I => \N__34280\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__34353\,
            I => \N__34280\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__34348\,
            I => \N__34280\
        );

    \I__6992\ : Span4Mux_v
    port map (
            O => \N__34343\,
            I => \N__34269\
        );

    \I__6991\ : Span4Mux_v
    port map (
            O => \N__34338\,
            I => \N__34269\
        );

    \I__6990\ : Span4Mux_h
    port map (
            O => \N__34331\,
            I => \N__34269\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__34324\,
            I => \N__34269\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__34315\,
            I => \N__34269\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__34312\,
            I => \N__34262\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__34305\,
            I => \N__34262\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__34296\,
            I => \N__34262\
        );

    \I__6984\ : Span4Mux_v
    port map (
            O => \N__34293\,
            I => \N__34259\
        );

    \I__6983\ : InMux
    port map (
            O => \N__34292\,
            I => \N__34256\
        );

    \I__6982\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34253\
        );

    \I__6981\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34250\
        );

    \I__6980\ : Span4Mux_h
    port map (
            O => \N__34287\,
            I => \N__34245\
        );

    \I__6979\ : Span4Mux_h
    port map (
            O => \N__34280\,
            I => \N__34245\
        );

    \I__6978\ : Span4Mux_v
    port map (
            O => \N__34269\,
            I => \N__34242\
        );

    \I__6977\ : Span12Mux_s11_v
    port map (
            O => \N__34262\,
            I => \N__34239\
        );

    \I__6976\ : Sp12to4
    port map (
            O => \N__34259\,
            I => \N__34236\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__34256\,
            I => \N__34229\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__34253\,
            I => \N__34229\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__34250\,
            I => \N__34229\
        );

    \I__6972\ : Sp12to4
    port map (
            O => \N__34245\,
            I => \N__34226\
        );

    \I__6971\ : Span4Mux_h
    port map (
            O => \N__34242\,
            I => \N__34223\
        );

    \I__6970\ : Span12Mux_v
    port map (
            O => \N__34239\,
            I => \N__34216\
        );

    \I__6969\ : Span12Mux_h
    port map (
            O => \N__34236\,
            I => \N__34216\
        );

    \I__6968\ : Span12Mux_s6_v
    port map (
            O => \N__34229\,
            I => \N__34216\
        );

    \I__6967\ : Odrv12
    port map (
            O => \N__34226\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6966\ : Odrv4
    port map (
            O => \N__34223\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6965\ : Odrv12
    port map (
            O => \N__34216\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6964\ : CascadeMux
    port map (
            O => \N__34209\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__6963\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34202\
        );

    \I__6962\ : InMux
    port map (
            O => \N__34205\,
            I => \N__34199\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__34202\,
            I => \N__34196\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__34199\,
            I => \N__34193\
        );

    \I__6959\ : Span4Mux_h
    port map (
            O => \N__34196\,
            I => \N__34190\
        );

    \I__6958\ : Span4Mux_v
    port map (
            O => \N__34193\,
            I => \N__34187\
        );

    \I__6957\ : Span4Mux_v
    port map (
            O => \N__34190\,
            I => \N__34184\
        );

    \I__6956\ : Odrv4
    port map (
            O => \N__34187\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__6955\ : Odrv4
    port map (
            O => \N__34184\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__6954\ : CascadeMux
    port map (
            O => \N__34179\,
            I => \N__34175\
        );

    \I__6953\ : CascadeMux
    port map (
            O => \N__34178\,
            I => \N__34172\
        );

    \I__6952\ : InMux
    port map (
            O => \N__34175\,
            I => \N__34169\
        );

    \I__6951\ : InMux
    port map (
            O => \N__34172\,
            I => \N__34166\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__34169\,
            I => \N__34161\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__34166\,
            I => \N__34161\
        );

    \I__6948\ : Span4Mux_h
    port map (
            O => \N__34161\,
            I => \N__34158\
        );

    \I__6947\ : Span4Mux_h
    port map (
            O => \N__34158\,
            I => \N__34155\
        );

    \I__6946\ : Odrv4
    port map (
            O => \N__34155\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__6945\ : CascadeMux
    port map (
            O => \N__34152\,
            I => \N__34149\
        );

    \I__6944\ : InMux
    port map (
            O => \N__34149\,
            I => \N__34146\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__34146\,
            I => \N__34141\
        );

    \I__6942\ : CascadeMux
    port map (
            O => \N__34145\,
            I => \N__34138\
        );

    \I__6941\ : InMux
    port map (
            O => \N__34144\,
            I => \N__34135\
        );

    \I__6940\ : Span4Mux_h
    port map (
            O => \N__34141\,
            I => \N__34132\
        );

    \I__6939\ : InMux
    port map (
            O => \N__34138\,
            I => \N__34129\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__34135\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__6937\ : Odrv4
    port map (
            O => \N__34132\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__34129\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__6935\ : InMux
    port map (
            O => \N__34122\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__6934\ : InMux
    port map (
            O => \N__34119\,
            I => \N__34113\
        );

    \I__6933\ : InMux
    port map (
            O => \N__34118\,
            I => \N__34113\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__34113\,
            I => \N__34109\
        );

    \I__6931\ : InMux
    port map (
            O => \N__34112\,
            I => \N__34106\
        );

    \I__6930\ : Span4Mux_v
    port map (
            O => \N__34109\,
            I => \N__34103\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__34106\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__6928\ : Odrv4
    port map (
            O => \N__34103\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__6927\ : InMux
    port map (
            O => \N__34098\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__6926\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34088\
        );

    \I__6925\ : InMux
    port map (
            O => \N__34094\,
            I => \N__34088\
        );

    \I__6924\ : InMux
    port map (
            O => \N__34093\,
            I => \N__34085\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__34088\,
            I => \N__34082\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__34085\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__6921\ : Odrv4
    port map (
            O => \N__34082\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__6920\ : InMux
    port map (
            O => \N__34077\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__6919\ : CascadeMux
    port map (
            O => \N__34074\,
            I => \N__34070\
        );

    \I__6918\ : CascadeMux
    port map (
            O => \N__34073\,
            I => \N__34067\
        );

    \I__6917\ : InMux
    port map (
            O => \N__34070\,
            I => \N__34062\
        );

    \I__6916\ : InMux
    port map (
            O => \N__34067\,
            I => \N__34062\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__34062\,
            I => \N__34058\
        );

    \I__6914\ : InMux
    port map (
            O => \N__34061\,
            I => \N__34055\
        );

    \I__6913\ : Span4Mux_h
    port map (
            O => \N__34058\,
            I => \N__34052\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__34055\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__6911\ : Odrv4
    port map (
            O => \N__34052\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__6910\ : InMux
    port map (
            O => \N__34047\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__6909\ : CascadeMux
    port map (
            O => \N__34044\,
            I => \N__34040\
        );

    \I__6908\ : CascadeMux
    port map (
            O => \N__34043\,
            I => \N__34037\
        );

    \I__6907\ : InMux
    port map (
            O => \N__34040\,
            I => \N__34031\
        );

    \I__6906\ : InMux
    port map (
            O => \N__34037\,
            I => \N__34031\
        );

    \I__6905\ : InMux
    port map (
            O => \N__34036\,
            I => \N__34028\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__34031\,
            I => \N__34025\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__34028\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__6902\ : Odrv4
    port map (
            O => \N__34025\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__6901\ : InMux
    port map (
            O => \N__34020\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__6900\ : InMux
    port map (
            O => \N__34017\,
            I => \N__34010\
        );

    \I__6899\ : InMux
    port map (
            O => \N__34016\,
            I => \N__34010\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34015\,
            I => \N__34007\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__34010\,
            I => \N__34004\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__34007\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__6895\ : Odrv4
    port map (
            O => \N__34004\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__6894\ : InMux
    port map (
            O => \N__33999\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__6893\ : CascadeMux
    port map (
            O => \N__33996\,
            I => \N__33992\
        );

    \I__6892\ : InMux
    port map (
            O => \N__33995\,
            I => \N__33989\
        );

    \I__6891\ : InMux
    port map (
            O => \N__33992\,
            I => \N__33985\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__33989\,
            I => \N__33982\
        );

    \I__6889\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33979\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__33985\,
            I => \N__33974\
        );

    \I__6887\ : Span4Mux_h
    port map (
            O => \N__33982\,
            I => \N__33974\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__33979\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__6885\ : Odrv4
    port map (
            O => \N__33974\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__6884\ : InMux
    port map (
            O => \N__33969\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__6883\ : CascadeMux
    port map (
            O => \N__33966\,
            I => \N__33963\
        );

    \I__6882\ : InMux
    port map (
            O => \N__33963\,
            I => \N__33958\
        );

    \I__6881\ : CascadeMux
    port map (
            O => \N__33962\,
            I => \N__33955\
        );

    \I__6880\ : InMux
    port map (
            O => \N__33961\,
            I => \N__33952\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__33958\,
            I => \N__33949\
        );

    \I__6878\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33946\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__33952\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__6876\ : Odrv4
    port map (
            O => \N__33949\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__33946\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__6874\ : InMux
    port map (
            O => \N__33939\,
            I => \bfn_14_16_0_\
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__33936\,
            I => \N__33933\
        );

    \I__6872\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33930\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__33930\,
            I => \N__33926\
        );

    \I__6870\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33922\
        );

    \I__6869\ : Span4Mux_v
    port map (
            O => \N__33926\,
            I => \N__33919\
        );

    \I__6868\ : InMux
    port map (
            O => \N__33925\,
            I => \N__33916\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__33922\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__6866\ : Odrv4
    port map (
            O => \N__33919\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__33916\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__6864\ : CascadeMux
    port map (
            O => \N__33909\,
            I => \N__33906\
        );

    \I__6863\ : InMux
    port map (
            O => \N__33906\,
            I => \N__33903\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__33903\,
            I => \N__33898\
        );

    \I__6861\ : CascadeMux
    port map (
            O => \N__33902\,
            I => \N__33895\
        );

    \I__6860\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33892\
        );

    \I__6859\ : Span4Mux_h
    port map (
            O => \N__33898\,
            I => \N__33889\
        );

    \I__6858\ : InMux
    port map (
            O => \N__33895\,
            I => \N__33886\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__33892\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__6856\ : Odrv4
    port map (
            O => \N__33889\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__33886\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__6854\ : InMux
    port map (
            O => \N__33879\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__6853\ : CascadeMux
    port map (
            O => \N__33876\,
            I => \N__33873\
        );

    \I__6852\ : InMux
    port map (
            O => \N__33873\,
            I => \N__33869\
        );

    \I__6851\ : InMux
    port map (
            O => \N__33872\,
            I => \N__33866\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__33869\,
            I => \N__33860\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__33866\,
            I => \N__33860\
        );

    \I__6848\ : InMux
    port map (
            O => \N__33865\,
            I => \N__33857\
        );

    \I__6847\ : Span4Mux_v
    port map (
            O => \N__33860\,
            I => \N__33854\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__33857\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__6845\ : Odrv4
    port map (
            O => \N__33854\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__6844\ : InMux
    port map (
            O => \N__33849\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__6843\ : InMux
    port map (
            O => \N__33846\,
            I => \N__33839\
        );

    \I__6842\ : InMux
    port map (
            O => \N__33845\,
            I => \N__33839\
        );

    \I__6841\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33836\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__33839\,
            I => \N__33833\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__33836\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__33833\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__6837\ : InMux
    port map (
            O => \N__33828\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__6836\ : InMux
    port map (
            O => \N__33825\,
            I => \N__33818\
        );

    \I__6835\ : InMux
    port map (
            O => \N__33824\,
            I => \N__33818\
        );

    \I__6834\ : InMux
    port map (
            O => \N__33823\,
            I => \N__33815\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__33818\,
            I => \N__33812\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__33815\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__6831\ : Odrv4
    port map (
            O => \N__33812\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__6830\ : InMux
    port map (
            O => \N__33807\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__6829\ : CascadeMux
    port map (
            O => \N__33804\,
            I => \N__33800\
        );

    \I__6828\ : CascadeMux
    port map (
            O => \N__33803\,
            I => \N__33797\
        );

    \I__6827\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33791\
        );

    \I__6826\ : InMux
    port map (
            O => \N__33797\,
            I => \N__33791\
        );

    \I__6825\ : InMux
    port map (
            O => \N__33796\,
            I => \N__33788\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__33791\,
            I => \N__33785\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__33788\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__6822\ : Odrv4
    port map (
            O => \N__33785\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__6821\ : InMux
    port map (
            O => \N__33780\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__6820\ : CascadeMux
    port map (
            O => \N__33777\,
            I => \N__33773\
        );

    \I__6819\ : CascadeMux
    port map (
            O => \N__33776\,
            I => \N__33770\
        );

    \I__6818\ : InMux
    port map (
            O => \N__33773\,
            I => \N__33765\
        );

    \I__6817\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33765\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__33765\,
            I => \N__33761\
        );

    \I__6815\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33758\
        );

    \I__6814\ : Span4Mux_h
    port map (
            O => \N__33761\,
            I => \N__33755\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__33758\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__6812\ : Odrv4
    port map (
            O => \N__33755\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__6811\ : InMux
    port map (
            O => \N__33750\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__6810\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33741\
        );

    \I__6809\ : InMux
    port map (
            O => \N__33746\,
            I => \N__33741\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__33741\,
            I => \N__33737\
        );

    \I__6807\ : InMux
    port map (
            O => \N__33740\,
            I => \N__33734\
        );

    \I__6806\ : Span4Mux_h
    port map (
            O => \N__33737\,
            I => \N__33731\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__33734\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__6804\ : Odrv4
    port map (
            O => \N__33731\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__6803\ : InMux
    port map (
            O => \N__33726\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__6802\ : CascadeMux
    port map (
            O => \N__33723\,
            I => \N__33720\
        );

    \I__6801\ : InMux
    port map (
            O => \N__33720\,
            I => \N__33716\
        );

    \I__6800\ : InMux
    port map (
            O => \N__33719\,
            I => \N__33712\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__33716\,
            I => \N__33709\
        );

    \I__6798\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33706\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__33712\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__33709\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__33706\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__6794\ : InMux
    port map (
            O => \N__33699\,
            I => \bfn_14_15_0_\
        );

    \I__6793\ : InMux
    port map (
            O => \N__33696\,
            I => \N__33692\
        );

    \I__6792\ : InMux
    port map (
            O => \N__33695\,
            I => \N__33689\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__33692\,
            I => \N__33685\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__33689\,
            I => \N__33682\
        );

    \I__6789\ : InMux
    port map (
            O => \N__33688\,
            I => \N__33679\
        );

    \I__6788\ : Span4Mux_h
    port map (
            O => \N__33685\,
            I => \N__33676\
        );

    \I__6787\ : Odrv12
    port map (
            O => \N__33682\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__33679\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6785\ : Odrv4
    port map (
            O => \N__33676\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6784\ : InMux
    port map (
            O => \N__33669\,
            I => \bfn_14_13_0_\
        );

    \I__6783\ : InMux
    port map (
            O => \N__33666\,
            I => \N__33662\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__33665\,
            I => \N__33659\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__33662\,
            I => \N__33656\
        );

    \I__6780\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33653\
        );

    \I__6779\ : Span4Mux_v
    port map (
            O => \N__33656\,
            I => \N__33647\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__33653\,
            I => \N__33647\
        );

    \I__6777\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33644\
        );

    \I__6776\ : Span4Mux_h
    port map (
            O => \N__33647\,
            I => \N__33641\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__33644\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6774\ : Odrv4
    port map (
            O => \N__33641\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6773\ : InMux
    port map (
            O => \N__33636\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__6772\ : CascadeMux
    port map (
            O => \N__33633\,
            I => \N__33629\
        );

    \I__6771\ : CascadeMux
    port map (
            O => \N__33632\,
            I => \N__33626\
        );

    \I__6770\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33620\
        );

    \I__6769\ : InMux
    port map (
            O => \N__33626\,
            I => \N__33620\
        );

    \I__6768\ : InMux
    port map (
            O => \N__33625\,
            I => \N__33617\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__33620\,
            I => \N__33614\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__33617\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__6765\ : Odrv4
    port map (
            O => \N__33614\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__6764\ : InMux
    port map (
            O => \N__33609\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__6763\ : InMux
    port map (
            O => \N__33606\,
            I => \N__33599\
        );

    \I__6762\ : InMux
    port map (
            O => \N__33605\,
            I => \N__33599\
        );

    \I__6761\ : InMux
    port map (
            O => \N__33604\,
            I => \N__33596\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__33599\,
            I => \N__33593\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__33596\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__6758\ : Odrv4
    port map (
            O => \N__33593\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__6757\ : InMux
    port map (
            O => \N__33588\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__6756\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33578\
        );

    \I__6755\ : InMux
    port map (
            O => \N__33584\,
            I => \N__33578\
        );

    \I__6754\ : InMux
    port map (
            O => \N__33583\,
            I => \N__33575\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__33578\,
            I => \N__33572\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__33575\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__6751\ : Odrv4
    port map (
            O => \N__33572\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__6750\ : InMux
    port map (
            O => \N__33567\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__6749\ : CascadeMux
    port map (
            O => \N__33564\,
            I => \N__33560\
        );

    \I__6748\ : CascadeMux
    port map (
            O => \N__33563\,
            I => \N__33557\
        );

    \I__6747\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33551\
        );

    \I__6746\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33551\
        );

    \I__6745\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33548\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__33551\,
            I => \N__33545\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__33548\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__33545\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__6741\ : InMux
    port map (
            O => \N__33540\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__6740\ : CascadeMux
    port map (
            O => \N__33537\,
            I => \N__33534\
        );

    \I__6739\ : InMux
    port map (
            O => \N__33534\,
            I => \N__33530\
        );

    \I__6738\ : InMux
    port map (
            O => \N__33533\,
            I => \N__33526\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__33530\,
            I => \N__33523\
        );

    \I__6736\ : InMux
    port map (
            O => \N__33529\,
            I => \N__33520\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__33526\,
            I => \N__33517\
        );

    \I__6734\ : Span4Mux_h
    port map (
            O => \N__33523\,
            I => \N__33514\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__33520\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__6732\ : Odrv4
    port map (
            O => \N__33517\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__6731\ : Odrv4
    port map (
            O => \N__33514\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__6730\ : InMux
    port map (
            O => \N__33507\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__6729\ : InMux
    port map (
            O => \N__33504\,
            I => \N__33498\
        );

    \I__6728\ : InMux
    port map (
            O => \N__33503\,
            I => \N__33498\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__33498\,
            I => \N__33494\
        );

    \I__6726\ : InMux
    port map (
            O => \N__33497\,
            I => \N__33491\
        );

    \I__6725\ : Span4Mux_h
    port map (
            O => \N__33494\,
            I => \N__33488\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__33491\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__33488\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__6722\ : InMux
    port map (
            O => \N__33483\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__6721\ : CascadeMux
    port map (
            O => \N__33480\,
            I => \N__33477\
        );

    \I__6720\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33472\
        );

    \I__6719\ : CascadeMux
    port map (
            O => \N__33476\,
            I => \N__33469\
        );

    \I__6718\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33466\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__33472\,
            I => \N__33463\
        );

    \I__6716\ : InMux
    port map (
            O => \N__33469\,
            I => \N__33460\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__33466\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__33463\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__33460\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__6712\ : InMux
    port map (
            O => \N__33453\,
            I => \bfn_14_14_0_\
        );

    \I__6711\ : InMux
    port map (
            O => \N__33450\,
            I => \N__33447\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__33447\,
            I => \N__33444\
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__33444\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__33441\,
            I => \N__33436\
        );

    \I__6707\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33430\
        );

    \I__6706\ : CascadeMux
    port map (
            O => \N__33439\,
            I => \N__33427\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33436\,
            I => \N__33422\
        );

    \I__6704\ : InMux
    port map (
            O => \N__33435\,
            I => \N__33422\
        );

    \I__6703\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33419\
        );

    \I__6702\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33416\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__33430\,
            I => \N__33413\
        );

    \I__6700\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33410\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__33422\,
            I => \N__33405\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__33419\,
            I => \N__33405\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__33416\,
            I => \N__33402\
        );

    \I__6696\ : Span4Mux_h
    port map (
            O => \N__33413\,
            I => \N__33397\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__33410\,
            I => \N__33397\
        );

    \I__6694\ : Span4Mux_h
    port map (
            O => \N__33405\,
            I => \N__33394\
        );

    \I__6693\ : Odrv4
    port map (
            O => \N__33402\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__6692\ : Odrv4
    port map (
            O => \N__33397\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__6691\ : Odrv4
    port map (
            O => \N__33394\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__6690\ : CascadeMux
    port map (
            O => \N__33387\,
            I => \delay_measurement_inst.N_360_cascade_\
        );

    \I__6689\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33381\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__33381\,
            I => \N__33378\
        );

    \I__6687\ : Span4Mux_v
    port map (
            O => \N__33378\,
            I => \N__33373\
        );

    \I__6686\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33370\
        );

    \I__6685\ : InMux
    port map (
            O => \N__33376\,
            I => \N__33367\
        );

    \I__6684\ : Odrv4
    port map (
            O => \N__33373\,
            I => measured_delay_tr_9
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__33370\,
            I => measured_delay_tr_9
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__33367\,
            I => measured_delay_tr_9
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__33360\,
            I => \delay_measurement_inst.N_354_cascade_\
        );

    \I__6680\ : InMux
    port map (
            O => \N__33357\,
            I => \N__33353\
        );

    \I__6679\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33350\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__33353\,
            I => \N__33347\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__33350\,
            I => \N__33344\
        );

    \I__6676\ : Span4Mux_h
    port map (
            O => \N__33347\,
            I => \N__33340\
        );

    \I__6675\ : Span4Mux_v
    port map (
            O => \N__33344\,
            I => \N__33337\
        );

    \I__6674\ : InMux
    port map (
            O => \N__33343\,
            I => \N__33334\
        );

    \I__6673\ : Odrv4
    port map (
            O => \N__33340\,
            I => measured_delay_tr_10
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__33337\,
            I => measured_delay_tr_10
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__33334\,
            I => measured_delay_tr_10
        );

    \I__6670\ : InMux
    port map (
            O => \N__33327\,
            I => \N__33324\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__33324\,
            I => \N__33321\
        );

    \I__6668\ : Span4Mux_h
    port map (
            O => \N__33321\,
            I => \N__33316\
        );

    \I__6667\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33313\
        );

    \I__6666\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33310\
        );

    \I__6665\ : Odrv4
    port map (
            O => \N__33316\,
            I => measured_delay_tr_11
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__33313\,
            I => measured_delay_tr_11
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__33310\,
            I => measured_delay_tr_11
        );

    \I__6662\ : InMux
    port map (
            O => \N__33303\,
            I => \N__33299\
        );

    \I__6661\ : InMux
    port map (
            O => \N__33302\,
            I => \N__33296\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__33299\,
            I => \N__33293\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__33296\,
            I => \N__33290\
        );

    \I__6658\ : Span4Mux_h
    port map (
            O => \N__33293\,
            I => \N__33286\
        );

    \I__6657\ : Span4Mux_h
    port map (
            O => \N__33290\,
            I => \N__33283\
        );

    \I__6656\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33280\
        );

    \I__6655\ : Odrv4
    port map (
            O => \N__33286\,
            I => measured_delay_tr_12
        );

    \I__6654\ : Odrv4
    port map (
            O => \N__33283\,
            I => measured_delay_tr_12
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__33280\,
            I => measured_delay_tr_12
        );

    \I__6652\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33261\
        );

    \I__6651\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33261\
        );

    \I__6650\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33261\
        );

    \I__6649\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33261\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__33261\,
            I => \delay_measurement_inst.N_354\
        );

    \I__6647\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33254\
        );

    \I__6646\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33251\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__33254\,
            I => \N__33245\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__33251\,
            I => \N__33245\
        );

    \I__6643\ : CascadeMux
    port map (
            O => \N__33250\,
            I => \N__33242\
        );

    \I__6642\ : Span4Mux_h
    port map (
            O => \N__33245\,
            I => \N__33239\
        );

    \I__6641\ : InMux
    port map (
            O => \N__33242\,
            I => \N__33236\
        );

    \I__6640\ : Odrv4
    port map (
            O => \N__33239\,
            I => measured_delay_tr_13
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__33236\,
            I => measured_delay_tr_13
        );

    \I__6638\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33228\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__33228\,
            I => \N__33224\
        );

    \I__6636\ : InMux
    port map (
            O => \N__33227\,
            I => \N__33221\
        );

    \I__6635\ : Span12Mux_v
    port map (
            O => \N__33224\,
            I => \N__33218\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__33221\,
            I => \N__33215\
        );

    \I__6633\ : Span12Mux_h
    port map (
            O => \N__33218\,
            I => \N__33212\
        );

    \I__6632\ : Span4Mux_s2_h
    port map (
            O => \N__33215\,
            I => \N__33209\
        );

    \I__6631\ : Odrv12
    port map (
            O => \N__33212\,
            I => pwm_duty_input_1
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__33209\,
            I => pwm_duty_input_1
        );

    \I__6629\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33201\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__33201\,
            I => \N__33197\
        );

    \I__6627\ : InMux
    port map (
            O => \N__33200\,
            I => \N__33194\
        );

    \I__6626\ : Span12Mux_v
    port map (
            O => \N__33197\,
            I => \N__33191\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__33194\,
            I => \N__33188\
        );

    \I__6624\ : Span12Mux_h
    port map (
            O => \N__33191\,
            I => \N__33185\
        );

    \I__6623\ : Span4Mux_v
    port map (
            O => \N__33188\,
            I => \N__33182\
        );

    \I__6622\ : Odrv12
    port map (
            O => \N__33185\,
            I => pwm_duty_input_0
        );

    \I__6621\ : Odrv4
    port map (
            O => \N__33182\,
            I => pwm_duty_input_0
        );

    \I__6620\ : InMux
    port map (
            O => \N__33177\,
            I => \N__33174\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__33174\,
            I => \N__33171\
        );

    \I__6618\ : Span4Mux_v
    port map (
            O => \N__33171\,
            I => \N__33167\
        );

    \I__6617\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33164\
        );

    \I__6616\ : Span4Mux_h
    port map (
            O => \N__33167\,
            I => \N__33161\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__33164\,
            I => \N__33158\
        );

    \I__6614\ : Sp12to4
    port map (
            O => \N__33161\,
            I => \N__33155\
        );

    \I__6613\ : Span4Mux_v
    port map (
            O => \N__33158\,
            I => \N__33152\
        );

    \I__6612\ : Odrv12
    port map (
            O => \N__33155\,
            I => pwm_duty_input_2
        );

    \I__6611\ : Odrv4
    port map (
            O => \N__33152\,
            I => pwm_duty_input_2
        );

    \I__6610\ : InMux
    port map (
            O => \N__33147\,
            I => \N__33144\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__33144\,
            I => \N__33141\
        );

    \I__6608\ : Span12Mux_s8_h
    port map (
            O => \N__33141\,
            I => \N__33138\
        );

    \I__6607\ : Odrv12
    port map (
            O => \N__33138\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__6606\ : CascadeMux
    port map (
            O => \N__33135\,
            I => \phase_controller_inst1.stoper_tr.time_passed11_cascade_\
        );

    \I__6605\ : CascadeMux
    port map (
            O => \N__33132\,
            I => \N__33128\
        );

    \I__6604\ : CascadeMux
    port map (
            O => \N__33131\,
            I => \N__33124\
        );

    \I__6603\ : InMux
    port map (
            O => \N__33128\,
            I => \N__33121\
        );

    \I__6602\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33118\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33124\,
            I => \N__33115\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__33121\,
            I => \N__33110\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__33118\,
            I => \N__33110\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__33115\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__6597\ : Odrv4
    port map (
            O => \N__33110\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__6596\ : CascadeMux
    port map (
            O => \N__33105\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_\
        );

    \I__6595\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33098\
        );

    \I__6594\ : InMux
    port map (
            O => \N__33101\,
            I => \N__33095\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__33098\,
            I => \N__33092\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__33095\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\
        );

    \I__6591\ : Odrv4
    port map (
            O => \N__33092\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\
        );

    \I__6590\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33084\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__33084\,
            I => \N__33081\
        );

    \I__6588\ : Span4Mux_v
    port map (
            O => \N__33081\,
            I => \N__33078\
        );

    \I__6587\ : Odrv4
    port map (
            O => \N__33078\,
            I => delay_tr_input_c
        );

    \I__6586\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33072\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__33072\,
            I => delay_tr_d1
        );

    \I__6584\ : InMux
    port map (
            O => \N__33069\,
            I => \N__33063\
        );

    \I__6583\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33063\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__33063\,
            I => \N__33058\
        );

    \I__6581\ : InMux
    port map (
            O => \N__33062\,
            I => \N__33055\
        );

    \I__6580\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33052\
        );

    \I__6579\ : Span4Mux_v
    port map (
            O => \N__33058\,
            I => \N__33047\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__33055\,
            I => \N__33047\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__33052\,
            I => delay_tr_d2
        );

    \I__6576\ : Odrv4
    port map (
            O => \N__33047\,
            I => delay_tr_d2
        );

    \I__6575\ : InMux
    port map (
            O => \N__33042\,
            I => \N__33039\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__33039\,
            I => \N__33036\
        );

    \I__6573\ : Span4Mux_h
    port map (
            O => \N__33036\,
            I => \N__33033\
        );

    \I__6572\ : Span4Mux_h
    port map (
            O => \N__33033\,
            I => \N__33030\
        );

    \I__6571\ : Sp12to4
    port map (
            O => \N__33030\,
            I => \N__33027\
        );

    \I__6570\ : Odrv12
    port map (
            O => \N__33027\,
            I => il_min_comp1_c
        );

    \I__6569\ : CascadeMux
    port map (
            O => \N__33024\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__6568\ : IoInMux
    port map (
            O => \N__33021\,
            I => \N__33018\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__33018\,
            I => \N__33015\
        );

    \I__6566\ : Span4Mux_s1_v
    port map (
            O => \N__33015\,
            I => \N__33012\
        );

    \I__6565\ : Span4Mux_v
    port map (
            O => \N__33012\,
            I => \N__33009\
        );

    \I__6564\ : Span4Mux_v
    port map (
            O => \N__33009\,
            I => \N__33004\
        );

    \I__6563\ : InMux
    port map (
            O => \N__33008\,
            I => \N__32999\
        );

    \I__6562\ : InMux
    port map (
            O => \N__33007\,
            I => \N__32999\
        );

    \I__6561\ : Odrv4
    port map (
            O => \N__33004\,
            I => s1_phy_c
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__32999\,
            I => s1_phy_c
        );

    \I__6559\ : InMux
    port map (
            O => \N__32994\,
            I => \N__32990\
        );

    \I__6558\ : InMux
    port map (
            O => \N__32993\,
            I => \N__32987\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__32990\,
            I => \N__32982\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__32987\,
            I => \N__32982\
        );

    \I__6555\ : Span4Mux_h
    port map (
            O => \N__32982\,
            I => \N__32979\
        );

    \I__6554\ : Span4Mux_v
    port map (
            O => \N__32979\,
            I => \N__32975\
        );

    \I__6553\ : InMux
    port map (
            O => \N__32978\,
            I => \N__32972\
        );

    \I__6552\ : Odrv4
    port map (
            O => \N__32975\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__32972\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__6550\ : CEMux
    port map (
            O => \N__32967\,
            I => \N__32946\
        );

    \I__6549\ : CEMux
    port map (
            O => \N__32966\,
            I => \N__32946\
        );

    \I__6548\ : CEMux
    port map (
            O => \N__32965\,
            I => \N__32946\
        );

    \I__6547\ : CEMux
    port map (
            O => \N__32964\,
            I => \N__32946\
        );

    \I__6546\ : CEMux
    port map (
            O => \N__32963\,
            I => \N__32946\
        );

    \I__6545\ : CEMux
    port map (
            O => \N__32962\,
            I => \N__32946\
        );

    \I__6544\ : CEMux
    port map (
            O => \N__32961\,
            I => \N__32946\
        );

    \I__6543\ : GlobalMux
    port map (
            O => \N__32946\,
            I => \N__32943\
        );

    \I__6542\ : gio2CtrlBuf
    port map (
            O => \N__32943\,
            I => \current_shift_inst.timer_s1.N_185_i_g\
        );

    \I__6541\ : InMux
    port map (
            O => \N__32940\,
            I => \N__32936\
        );

    \I__6540\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32933\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__32936\,
            I => \N__32927\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__32933\,
            I => \N__32927\
        );

    \I__6537\ : InMux
    port map (
            O => \N__32932\,
            I => \N__32924\
        );

    \I__6536\ : Span4Mux_v
    port map (
            O => \N__32927\,
            I => \N__32918\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__32924\,
            I => \N__32918\
        );

    \I__6534\ : InMux
    port map (
            O => \N__32923\,
            I => \N__32915\
        );

    \I__6533\ : Odrv4
    port map (
            O => \N__32918\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__32915\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__6531\ : InMux
    port map (
            O => \N__32910\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__6530\ : InMux
    port map (
            O => \N__32907\,
            I => \N__32903\
        );

    \I__6529\ : InMux
    port map (
            O => \N__32906\,
            I => \N__32900\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__32903\,
            I => \N__32896\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__32900\,
            I => \N__32893\
        );

    \I__6526\ : InMux
    port map (
            O => \N__32899\,
            I => \N__32890\
        );

    \I__6525\ : Span4Mux_h
    port map (
            O => \N__32896\,
            I => \N__32886\
        );

    \I__6524\ : Span4Mux_v
    port map (
            O => \N__32893\,
            I => \N__32881\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__32890\,
            I => \N__32881\
        );

    \I__6522\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32878\
        );

    \I__6521\ : Odrv4
    port map (
            O => \N__32886\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__6520\ : Odrv4
    port map (
            O => \N__32881\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__32878\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__6518\ : InMux
    port map (
            O => \N__32871\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__6517\ : InMux
    port map (
            O => \N__32868\,
            I => \N__32864\
        );

    \I__6516\ : InMux
    port map (
            O => \N__32867\,
            I => \N__32860\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__32864\,
            I => \N__32857\
        );

    \I__6514\ : InMux
    port map (
            O => \N__32863\,
            I => \N__32853\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__32860\,
            I => \N__32850\
        );

    \I__6512\ : Sp12to4
    port map (
            O => \N__32857\,
            I => \N__32847\
        );

    \I__6511\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32844\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__32853\,
            I => \N__32841\
        );

    \I__6509\ : Span4Mux_h
    port map (
            O => \N__32850\,
            I => \N__32838\
        );

    \I__6508\ : Span12Mux_v
    port map (
            O => \N__32847\,
            I => \N__32831\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__32844\,
            I => \N__32831\
        );

    \I__6506\ : Span12Mux_v
    port map (
            O => \N__32841\,
            I => \N__32831\
        );

    \I__6505\ : Odrv4
    port map (
            O => \N__32838\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__6504\ : Odrv12
    port map (
            O => \N__32831\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__6503\ : InMux
    port map (
            O => \N__32826\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__32823\,
            I => \N__32820\
        );

    \I__6501\ : InMux
    port map (
            O => \N__32820\,
            I => \N__32813\
        );

    \I__6500\ : InMux
    port map (
            O => \N__32819\,
            I => \N__32813\
        );

    \I__6499\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32810\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__32813\,
            I => \N__32807\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__32810\,
            I => \N__32804\
        );

    \I__6496\ : Span4Mux_v
    port map (
            O => \N__32807\,
            I => \N__32800\
        );

    \I__6495\ : Span4Mux_h
    port map (
            O => \N__32804\,
            I => \N__32797\
        );

    \I__6494\ : InMux
    port map (
            O => \N__32803\,
            I => \N__32794\
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__32800\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__6492\ : Odrv4
    port map (
            O => \N__32797\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__32794\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__6490\ : InMux
    port map (
            O => \N__32787\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__6489\ : CascadeMux
    port map (
            O => \N__32784\,
            I => \N__32780\
        );

    \I__6488\ : InMux
    port map (
            O => \N__32783\,
            I => \N__32772\
        );

    \I__6487\ : InMux
    port map (
            O => \N__32780\,
            I => \N__32772\
        );

    \I__6486\ : InMux
    port map (
            O => \N__32779\,
            I => \N__32772\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__32772\,
            I => \N__32768\
        );

    \I__6484\ : InMux
    port map (
            O => \N__32771\,
            I => \N__32765\
        );

    \I__6483\ : Odrv4
    port map (
            O => \N__32768\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__32765\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__6481\ : InMux
    port map (
            O => \N__32760\,
            I => \bfn_13_18_0_\
        );

    \I__6480\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32753\
        );

    \I__6479\ : CascadeMux
    port map (
            O => \N__32756\,
            I => \N__32750\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__32753\,
            I => \N__32746\
        );

    \I__6477\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32741\
        );

    \I__6476\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32741\
        );

    \I__6475\ : Span12Mux_v
    port map (
            O => \N__32746\,
            I => \N__32735\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__32741\,
            I => \N__32735\
        );

    \I__6473\ : InMux
    port map (
            O => \N__32740\,
            I => \N__32732\
        );

    \I__6472\ : Odrv12
    port map (
            O => \N__32735\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__32732\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__6470\ : InMux
    port map (
            O => \N__32727\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__6469\ : InMux
    port map (
            O => \N__32724\,
            I => \N__32720\
        );

    \I__6468\ : CascadeMux
    port map (
            O => \N__32723\,
            I => \N__32717\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__32720\,
            I => \N__32713\
        );

    \I__6466\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32708\
        );

    \I__6465\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32708\
        );

    \I__6464\ : Span4Mux_h
    port map (
            O => \N__32713\,
            I => \N__32704\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__32708\,
            I => \N__32701\
        );

    \I__6462\ : InMux
    port map (
            O => \N__32707\,
            I => \N__32698\
        );

    \I__6461\ : Odrv4
    port map (
            O => \N__32704\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__32701\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__32698\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__6458\ : InMux
    port map (
            O => \N__32691\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__6457\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32684\
        );

    \I__6456\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32681\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__32684\,
            I => \N__32676\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__32681\,
            I => \N__32673\
        );

    \I__6453\ : InMux
    port map (
            O => \N__32680\,
            I => \N__32670\
        );

    \I__6452\ : InMux
    port map (
            O => \N__32679\,
            I => \N__32667\
        );

    \I__6451\ : Span4Mux_h
    port map (
            O => \N__32676\,
            I => \N__32664\
        );

    \I__6450\ : Span4Mux_v
    port map (
            O => \N__32673\,
            I => \N__32657\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__32670\,
            I => \N__32657\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__32667\,
            I => \N__32657\
        );

    \I__6447\ : Odrv4
    port map (
            O => \N__32664\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__6446\ : Odrv4
    port map (
            O => \N__32657\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__6445\ : InMux
    port map (
            O => \N__32652\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__6444\ : InMux
    port map (
            O => \N__32649\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__6443\ : InMux
    port map (
            O => \N__32646\,
            I => \N__32641\
        );

    \I__6442\ : InMux
    port map (
            O => \N__32645\,
            I => \N__32638\
        );

    \I__6441\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32635\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__32641\,
            I => \N__32630\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__32638\,
            I => \N__32630\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__32635\,
            I => \N__32627\
        );

    \I__6437\ : Span4Mux_v
    port map (
            O => \N__32630\,
            I => \N__32623\
        );

    \I__6436\ : Span4Mux_h
    port map (
            O => \N__32627\,
            I => \N__32620\
        );

    \I__6435\ : InMux
    port map (
            O => \N__32626\,
            I => \N__32617\
        );

    \I__6434\ : Odrv4
    port map (
            O => \N__32623\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__6433\ : Odrv4
    port map (
            O => \N__32620\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__32617\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__6431\ : InMux
    port map (
            O => \N__32610\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__6430\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32602\
        );

    \I__6429\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32599\
        );

    \I__6428\ : InMux
    port map (
            O => \N__32605\,
            I => \N__32596\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__32602\,
            I => \N__32591\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__32599\,
            I => \N__32591\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__32596\,
            I => \N__32588\
        );

    \I__6424\ : Span4Mux_v
    port map (
            O => \N__32591\,
            I => \N__32584\
        );

    \I__6423\ : Span4Mux_h
    port map (
            O => \N__32588\,
            I => \N__32581\
        );

    \I__6422\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32578\
        );

    \I__6421\ : Odrv4
    port map (
            O => \N__32584\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__6420\ : Odrv4
    port map (
            O => \N__32581\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__32578\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__6418\ : InMux
    port map (
            O => \N__32571\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__6417\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32562\
        );

    \I__6416\ : InMux
    port map (
            O => \N__32567\,
            I => \N__32559\
        );

    \I__6415\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32556\
        );

    \I__6414\ : InMux
    port map (
            O => \N__32565\,
            I => \N__32553\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__32562\,
            I => \N__32550\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__32559\,
            I => \N__32545\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__32556\,
            I => \N__32545\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__32553\,
            I => \N__32542\
        );

    \I__6409\ : Span4Mux_h
    port map (
            O => \N__32550\,
            I => \N__32539\
        );

    \I__6408\ : Span12Mux_v
    port map (
            O => \N__32545\,
            I => \N__32534\
        );

    \I__6407\ : Span12Mux_v
    port map (
            O => \N__32542\,
            I => \N__32534\
        );

    \I__6406\ : Odrv4
    port map (
            O => \N__32539\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__6405\ : Odrv12
    port map (
            O => \N__32534\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__6404\ : InMux
    port map (
            O => \N__32529\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__6403\ : InMux
    port map (
            O => \N__32526\,
            I => \N__32523\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__32523\,
            I => \N__32518\
        );

    \I__6401\ : InMux
    port map (
            O => \N__32522\,
            I => \N__32515\
        );

    \I__6400\ : InMux
    port map (
            O => \N__32521\,
            I => \N__32512\
        );

    \I__6399\ : Span4Mux_h
    port map (
            O => \N__32518\,
            I => \N__32506\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__32515\,
            I => \N__32506\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__32512\,
            I => \N__32503\
        );

    \I__6396\ : InMux
    port map (
            O => \N__32511\,
            I => \N__32500\
        );

    \I__6395\ : Span4Mux_v
    port map (
            O => \N__32506\,
            I => \N__32495\
        );

    \I__6394\ : Span4Mux_h
    port map (
            O => \N__32503\,
            I => \N__32495\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__32500\,
            I => \N__32492\
        );

    \I__6392\ : Odrv4
    port map (
            O => \N__32495\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__6391\ : Odrv12
    port map (
            O => \N__32492\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__6390\ : InMux
    port map (
            O => \N__32487\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__6389\ : InMux
    port map (
            O => \N__32484\,
            I => \N__32481\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__32481\,
            I => \N__32477\
        );

    \I__6387\ : CascadeMux
    port map (
            O => \N__32480\,
            I => \N__32474\
        );

    \I__6386\ : Sp12to4
    port map (
            O => \N__32477\,
            I => \N__32470\
        );

    \I__6385\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32465\
        );

    \I__6384\ : InMux
    port map (
            O => \N__32473\,
            I => \N__32465\
        );

    \I__6383\ : Span12Mux_v
    port map (
            O => \N__32470\,
            I => \N__32459\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__32465\,
            I => \N__32459\
        );

    \I__6381\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32456\
        );

    \I__6380\ : Odrv12
    port map (
            O => \N__32459\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__32456\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__6378\ : InMux
    port map (
            O => \N__32451\,
            I => \bfn_13_17_0_\
        );

    \I__6377\ : InMux
    port map (
            O => \N__32448\,
            I => \N__32443\
        );

    \I__6376\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32440\
        );

    \I__6375\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32437\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__32443\,
            I => \N__32432\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__32440\,
            I => \N__32432\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__32437\,
            I => \N__32429\
        );

    \I__6371\ : Span4Mux_v
    port map (
            O => \N__32432\,
            I => \N__32423\
        );

    \I__6370\ : Span4Mux_v
    port map (
            O => \N__32429\,
            I => \N__32423\
        );

    \I__6369\ : InMux
    port map (
            O => \N__32428\,
            I => \N__32420\
        );

    \I__6368\ : Odrv4
    port map (
            O => \N__32423\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__32420\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__6366\ : InMux
    port map (
            O => \N__32415\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__6365\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32408\
        );

    \I__6364\ : InMux
    port map (
            O => \N__32411\,
            I => \N__32405\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__32408\,
            I => \N__32401\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__32405\,
            I => \N__32398\
        );

    \I__6361\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32395\
        );

    \I__6360\ : Span4Mux_h
    port map (
            O => \N__32401\,
            I => \N__32391\
        );

    \I__6359\ : Span4Mux_v
    port map (
            O => \N__32398\,
            I => \N__32386\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__32395\,
            I => \N__32386\
        );

    \I__6357\ : InMux
    port map (
            O => \N__32394\,
            I => \N__32383\
        );

    \I__6356\ : Odrv4
    port map (
            O => \N__32391\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__32386\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__32383\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__6353\ : InMux
    port map (
            O => \N__32376\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__6352\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32370\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__32370\,
            I => \N__32366\
        );

    \I__6350\ : InMux
    port map (
            O => \N__32369\,
            I => \N__32363\
        );

    \I__6349\ : Span4Mux_h
    port map (
            O => \N__32366\,
            I => \N__32358\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__32363\,
            I => \N__32358\
        );

    \I__6347\ : Span4Mux_v
    port map (
            O => \N__32358\,
            I => \N__32353\
        );

    \I__6346\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32350\
        );

    \I__6345\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32347\
        );

    \I__6344\ : Odrv4
    port map (
            O => \N__32353\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__32350\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__32347\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__6341\ : InMux
    port map (
            O => \N__32340\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__6340\ : CascadeMux
    port map (
            O => \N__32337\,
            I => \N__32333\
        );

    \I__6339\ : CascadeMux
    port map (
            O => \N__32336\,
            I => \N__32329\
        );

    \I__6338\ : InMux
    port map (
            O => \N__32333\,
            I => \N__32326\
        );

    \I__6337\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32323\
        );

    \I__6336\ : InMux
    port map (
            O => \N__32329\,
            I => \N__32320\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__32326\,
            I => \N__32317\
        );

    \I__6334\ : LocalMux
    port map (
            O => \N__32323\,
            I => \N__32314\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__32320\,
            I => \N__32308\
        );

    \I__6332\ : Span4Mux_h
    port map (
            O => \N__32317\,
            I => \N__32308\
        );

    \I__6331\ : Span4Mux_h
    port map (
            O => \N__32314\,
            I => \N__32305\
        );

    \I__6330\ : InMux
    port map (
            O => \N__32313\,
            I => \N__32302\
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__32308\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__6328\ : Odrv4
    port map (
            O => \N__32305\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__32302\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__6326\ : InMux
    port map (
            O => \N__32295\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__6325\ : InMux
    port map (
            O => \N__32292\,
            I => \N__32288\
        );

    \I__6324\ : InMux
    port map (
            O => \N__32291\,
            I => \N__32284\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__32288\,
            I => \N__32281\
        );

    \I__6322\ : InMux
    port map (
            O => \N__32287\,
            I => \N__32278\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__32284\,
            I => \N__32275\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__32281\,
            I => \N__32272\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__32278\,
            I => \N__32269\
        );

    \I__6318\ : Span4Mux_v
    port map (
            O => \N__32275\,
            I => \N__32265\
        );

    \I__6317\ : Span4Mux_h
    port map (
            O => \N__32272\,
            I => \N__32260\
        );

    \I__6316\ : Span4Mux_h
    port map (
            O => \N__32269\,
            I => \N__32260\
        );

    \I__6315\ : InMux
    port map (
            O => \N__32268\,
            I => \N__32257\
        );

    \I__6314\ : Odrv4
    port map (
            O => \N__32265\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__6313\ : Odrv4
    port map (
            O => \N__32260\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__32257\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__6311\ : InMux
    port map (
            O => \N__32250\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__6310\ : InMux
    port map (
            O => \N__32247\,
            I => \N__32244\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__32244\,
            I => \N__32240\
        );

    \I__6308\ : InMux
    port map (
            O => \N__32243\,
            I => \N__32237\
        );

    \I__6307\ : Span4Mux_v
    port map (
            O => \N__32240\,
            I => \N__32231\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__32237\,
            I => \N__32231\
        );

    \I__6305\ : InMux
    port map (
            O => \N__32236\,
            I => \N__32228\
        );

    \I__6304\ : Span4Mux_v
    port map (
            O => \N__32231\,
            I => \N__32224\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__32228\,
            I => \N__32221\
        );

    \I__6302\ : InMux
    port map (
            O => \N__32227\,
            I => \N__32218\
        );

    \I__6301\ : Odrv4
    port map (
            O => \N__32224\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__6300\ : Odrv4
    port map (
            O => \N__32221\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__32218\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__6298\ : InMux
    port map (
            O => \N__32211\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__6297\ : CascadeMux
    port map (
            O => \N__32208\,
            I => \N__32205\
        );

    \I__6296\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32201\
        );

    \I__6295\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32198\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__32201\,
            I => \N__32194\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__32198\,
            I => \N__32191\
        );

    \I__6292\ : InMux
    port map (
            O => \N__32197\,
            I => \N__32188\
        );

    \I__6291\ : Span4Mux_v
    port map (
            O => \N__32194\,
            I => \N__32180\
        );

    \I__6290\ : Span4Mux_v
    port map (
            O => \N__32191\,
            I => \N__32180\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__32188\,
            I => \N__32180\
        );

    \I__6288\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32177\
        );

    \I__6287\ : Odrv4
    port map (
            O => \N__32180\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__32177\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__6285\ : InMux
    port map (
            O => \N__32172\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__6284\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32164\
        );

    \I__6283\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32161\
        );

    \I__6282\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32158\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__32164\,
            I => \N__32155\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__32161\,
            I => \N__32152\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__32158\,
            I => \N__32149\
        );

    \I__6278\ : Span4Mux_v
    port map (
            O => \N__32155\,
            I => \N__32145\
        );

    \I__6277\ : Span4Mux_v
    port map (
            O => \N__32152\,
            I => \N__32140\
        );

    \I__6276\ : Span4Mux_h
    port map (
            O => \N__32149\,
            I => \N__32140\
        );

    \I__6275\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32137\
        );

    \I__6274\ : Odrv4
    port map (
            O => \N__32145\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__6273\ : Odrv4
    port map (
            O => \N__32140\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__32137\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__6271\ : InMux
    port map (
            O => \N__32130\,
            I => \bfn_13_16_0_\
        );

    \I__6270\ : CascadeMux
    port map (
            O => \N__32127\,
            I => \N__32123\
        );

    \I__6269\ : InMux
    port map (
            O => \N__32126\,
            I => \N__32120\
        );

    \I__6268\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32116\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__32120\,
            I => \N__32113\
        );

    \I__6266\ : InMux
    port map (
            O => \N__32119\,
            I => \N__32110\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__32116\,
            I => \N__32105\
        );

    \I__6264\ : Span4Mux_v
    port map (
            O => \N__32113\,
            I => \N__32105\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__32110\,
            I => \N__32102\
        );

    \I__6262\ : Span4Mux_v
    port map (
            O => \N__32105\,
            I => \N__32096\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__32102\,
            I => \N__32096\
        );

    \I__6260\ : InMux
    port map (
            O => \N__32101\,
            I => \N__32093\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__32096\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__32093\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__6257\ : InMux
    port map (
            O => \N__32088\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__6256\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32081\
        );

    \I__6255\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32077\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__32081\,
            I => \N__32074\
        );

    \I__6253\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32071\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__32077\,
            I => \N__32068\
        );

    \I__6251\ : Span4Mux_v
    port map (
            O => \N__32074\,
            I => \N__32062\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__32071\,
            I => \N__32062\
        );

    \I__6249\ : Span4Mux_h
    port map (
            O => \N__32068\,
            I => \N__32059\
        );

    \I__6248\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32056\
        );

    \I__6247\ : Odrv4
    port map (
            O => \N__32062\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__6246\ : Odrv4
    port map (
            O => \N__32059\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__32056\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__6244\ : InMux
    port map (
            O => \N__32049\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__6243\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32042\
        );

    \I__6242\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32038\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__32042\,
            I => \N__32035\
        );

    \I__6240\ : InMux
    port map (
            O => \N__32041\,
            I => \N__32032\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__32038\,
            I => \N__32029\
        );

    \I__6238\ : Span4Mux_h
    port map (
            O => \N__32035\,
            I => \N__32026\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__32032\,
            I => \N__32023\
        );

    \I__6236\ : Span4Mux_h
    port map (
            O => \N__32029\,
            I => \N__32019\
        );

    \I__6235\ : Span4Mux_v
    port map (
            O => \N__32026\,
            I => \N__32014\
        );

    \I__6234\ : Span4Mux_h
    port map (
            O => \N__32023\,
            I => \N__32014\
        );

    \I__6233\ : InMux
    port map (
            O => \N__32022\,
            I => \N__32011\
        );

    \I__6232\ : Odrv4
    port map (
            O => \N__32019\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__6231\ : Odrv4
    port map (
            O => \N__32014\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__32011\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__6229\ : InMux
    port map (
            O => \N__32004\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__6228\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31993\
        );

    \I__6227\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31988\
        );

    \I__6226\ : InMux
    port map (
            O => \N__31999\,
            I => \N__31988\
        );

    \I__6225\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31983\
        );

    \I__6224\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31983\
        );

    \I__6223\ : InMux
    port map (
            O => \N__31996\,
            I => \N__31980\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__31993\,
            I => \N__31972\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__31988\,
            I => \N__31972\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__31983\,
            I => \N__31972\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__31980\,
            I => \N__31968\
        );

    \I__6218\ : InMux
    port map (
            O => \N__31979\,
            I => \N__31963\
        );

    \I__6217\ : Span4Mux_v
    port map (
            O => \N__31972\,
            I => \N__31960\
        );

    \I__6216\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31957\
        );

    \I__6215\ : Span4Mux_h
    port map (
            O => \N__31968\,
            I => \N__31954\
        );

    \I__6214\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31949\
        );

    \I__6213\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31949\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__31963\,
            I => measured_delay_tr_15
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__31960\,
            I => measured_delay_tr_15
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__31957\,
            I => measured_delay_tr_15
        );

    \I__6209\ : Odrv4
    port map (
            O => \N__31954\,
            I => measured_delay_tr_15
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__31949\,
            I => measured_delay_tr_15
        );

    \I__6207\ : InMux
    port map (
            O => \N__31938\,
            I => \N__31933\
        );

    \I__6206\ : InMux
    port map (
            O => \N__31937\,
            I => \N__31930\
        );

    \I__6205\ : InMux
    port map (
            O => \N__31936\,
            I => \N__31927\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__31933\,
            I => \N__31924\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__31930\,
            I => \N__31919\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__31927\,
            I => \N__31919\
        );

    \I__6201\ : Span4Mux_h
    port map (
            O => \N__31924\,
            I => \N__31914\
        );

    \I__6200\ : Span4Mux_h
    port map (
            O => \N__31919\,
            I => \N__31911\
        );

    \I__6199\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31908\
        );

    \I__6198\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31905\
        );

    \I__6197\ : Odrv4
    port map (
            O => \N__31914\,
            I => measured_delay_tr_14
        );

    \I__6196\ : Odrv4
    port map (
            O => \N__31911\,
            I => measured_delay_tr_14
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__31908\,
            I => measured_delay_tr_14
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__31905\,
            I => measured_delay_tr_14
        );

    \I__6193\ : CascadeMux
    port map (
            O => \N__31896\,
            I => \N__31892\
        );

    \I__6192\ : CascadeMux
    port map (
            O => \N__31895\,
            I => \N__31887\
        );

    \I__6191\ : InMux
    port map (
            O => \N__31892\,
            I => \N__31870\
        );

    \I__6190\ : InMux
    port map (
            O => \N__31891\,
            I => \N__31870\
        );

    \I__6189\ : InMux
    port map (
            O => \N__31890\,
            I => \N__31863\
        );

    \I__6188\ : InMux
    port map (
            O => \N__31887\,
            I => \N__31863\
        );

    \I__6187\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31863\
        );

    \I__6186\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31856\
        );

    \I__6185\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31856\
        );

    \I__6184\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31856\
        );

    \I__6183\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31847\
        );

    \I__6182\ : InMux
    port map (
            O => \N__31881\,
            I => \N__31847\
        );

    \I__6181\ : InMux
    port map (
            O => \N__31880\,
            I => \N__31847\
        );

    \I__6180\ : InMux
    port map (
            O => \N__31879\,
            I => \N__31847\
        );

    \I__6179\ : InMux
    port map (
            O => \N__31878\,
            I => \N__31838\
        );

    \I__6178\ : InMux
    port map (
            O => \N__31877\,
            I => \N__31838\
        );

    \I__6177\ : InMux
    port map (
            O => \N__31876\,
            I => \N__31838\
        );

    \I__6176\ : InMux
    port map (
            O => \N__31875\,
            I => \N__31838\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__31870\,
            I => \N__31833\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__31863\,
            I => \N__31833\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__31856\,
            I => \N__31830\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__31847\,
            I => \N__31827\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__31838\,
            I => \N__31824\
        );

    \I__6170\ : Span4Mux_h
    port map (
            O => \N__31833\,
            I => \N__31821\
        );

    \I__6169\ : Span4Mux_h
    port map (
            O => \N__31830\,
            I => \N__31814\
        );

    \I__6168\ : Span4Mux_v
    port map (
            O => \N__31827\,
            I => \N__31814\
        );

    \I__6167\ : Span4Mux_v
    port map (
            O => \N__31824\,
            I => \N__31814\
        );

    \I__6166\ : Odrv4
    port map (
            O => \N__31821\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__31814\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__6164\ : CascadeMux
    port map (
            O => \N__31809\,
            I => \N__31806\
        );

    \I__6163\ : InMux
    port map (
            O => \N__31806\,
            I => \N__31803\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__31803\,
            I => \delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14\
        );

    \I__6161\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31797\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__31797\,
            I => \N__31794\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__31794\,
            I => \N__31789\
        );

    \I__6158\ : InMux
    port map (
            O => \N__31793\,
            I => \N__31786\
        );

    \I__6157\ : InMux
    port map (
            O => \N__31792\,
            I => \N__31783\
        );

    \I__6156\ : Span4Mux_h
    port map (
            O => \N__31789\,
            I => \N__31780\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__31786\,
            I => \N__31777\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__31783\,
            I => \il_min_comp2_D2\
        );

    \I__6153\ : Odrv4
    port map (
            O => \N__31780\,
            I => \il_min_comp2_D2\
        );

    \I__6152\ : Odrv12
    port map (
            O => \N__31777\,
            I => \il_min_comp2_D2\
        );

    \I__6151\ : InMux
    port map (
            O => \N__31770\,
            I => \N__31767\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__31767\,
            I => \N__31764\
        );

    \I__6149\ : Span4Mux_h
    port map (
            O => \N__31764\,
            I => \N__31761\
        );

    \I__6148\ : Span4Mux_v
    port map (
            O => \N__31761\,
            I => \N__31756\
        );

    \I__6147\ : InMux
    port map (
            O => \N__31760\,
            I => \N__31753\
        );

    \I__6146\ : InMux
    port map (
            O => \N__31759\,
            I => \N__31750\
        );

    \I__6145\ : Odrv4
    port map (
            O => \N__31756\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__31753\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__31750\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__6142\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31740\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__31740\,
            I => \N__31736\
        );

    \I__6140\ : CascadeMux
    port map (
            O => \N__31739\,
            I => \N__31733\
        );

    \I__6139\ : Span4Mux_v
    port map (
            O => \N__31736\,
            I => \N__31730\
        );

    \I__6138\ : InMux
    port map (
            O => \N__31733\,
            I => \N__31727\
        );

    \I__6137\ : Span4Mux_v
    port map (
            O => \N__31730\,
            I => \N__31723\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__31727\,
            I => \N__31719\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__31726\,
            I => \N__31716\
        );

    \I__6134\ : Span4Mux_v
    port map (
            O => \N__31723\,
            I => \N__31713\
        );

    \I__6133\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31710\
        );

    \I__6132\ : Span4Mux_h
    port map (
            O => \N__31719\,
            I => \N__31707\
        );

    \I__6131\ : InMux
    port map (
            O => \N__31716\,
            I => \N__31704\
        );

    \I__6130\ : Span4Mux_v
    port map (
            O => \N__31713\,
            I => \N__31699\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__31710\,
            I => \N__31699\
        );

    \I__6128\ : Span4Mux_v
    port map (
            O => \N__31707\,
            I => \N__31692\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__31704\,
            I => \N__31692\
        );

    \I__6126\ : Span4Mux_h
    port map (
            O => \N__31699\,
            I => \N__31692\
        );

    \I__6125\ : Odrv4
    port map (
            O => \N__31692\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6124\ : InMux
    port map (
            O => \N__31689\,
            I => \N__31686\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__31686\,
            I => \N__31683\
        );

    \I__6122\ : Odrv4
    port map (
            O => \N__31683\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__6121\ : InMux
    port map (
            O => \N__31680\,
            I => \N__31676\
        );

    \I__6120\ : InMux
    port map (
            O => \N__31679\,
            I => \N__31673\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__31676\,
            I => \N__31669\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__31673\,
            I => \N__31666\
        );

    \I__6117\ : InMux
    port map (
            O => \N__31672\,
            I => \N__31663\
        );

    \I__6116\ : Span4Mux_v
    port map (
            O => \N__31669\,
            I => \N__31658\
        );

    \I__6115\ : Span4Mux_v
    port map (
            O => \N__31666\,
            I => \N__31658\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__31663\,
            I => \N__31654\
        );

    \I__6113\ : Span4Mux_h
    port map (
            O => \N__31658\,
            I => \N__31651\
        );

    \I__6112\ : InMux
    port map (
            O => \N__31657\,
            I => \N__31648\
        );

    \I__6111\ : Odrv4
    port map (
            O => \N__31654\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__31651\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__31648\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__6108\ : InMux
    port map (
            O => \N__31641\,
            I => \N__31638\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__31638\,
            I => \N__31635\
        );

    \I__6106\ : Span4Mux_v
    port map (
            O => \N__31635\,
            I => \N__31630\
        );

    \I__6105\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31625\
        );

    \I__6104\ : InMux
    port map (
            O => \N__31633\,
            I => \N__31625\
        );

    \I__6103\ : Sp12to4
    port map (
            O => \N__31630\,
            I => \N__31619\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__31625\,
            I => \N__31619\
        );

    \I__6101\ : InMux
    port map (
            O => \N__31624\,
            I => \N__31616\
        );

    \I__6100\ : Odrv12
    port map (
            O => \N__31619\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__31616\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__6098\ : InMux
    port map (
            O => \N__31611\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__6097\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31604\
        );

    \I__6096\ : InMux
    port map (
            O => \N__31607\,
            I => \N__31601\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__31604\,
            I => \N__31597\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__31601\,
            I => \N__31594\
        );

    \I__6093\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31591\
        );

    \I__6092\ : Span4Mux_h
    port map (
            O => \N__31597\,
            I => \N__31587\
        );

    \I__6091\ : Span4Mux_v
    port map (
            O => \N__31594\,
            I => \N__31584\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__31591\,
            I => \N__31581\
        );

    \I__6089\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31578\
        );

    \I__6088\ : Odrv4
    port map (
            O => \N__31587\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__6087\ : Odrv4
    port map (
            O => \N__31584\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__6086\ : Odrv12
    port map (
            O => \N__31581\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__31578\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__6084\ : InMux
    port map (
            O => \N__31569\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__6083\ : InMux
    port map (
            O => \N__31566\,
            I => \N__31563\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__31563\,
            I => \N__31559\
        );

    \I__6081\ : InMux
    port map (
            O => \N__31562\,
            I => \N__31556\
        );

    \I__6080\ : Span4Mux_v
    port map (
            O => \N__31559\,
            I => \N__31551\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__31556\,
            I => \N__31551\
        );

    \I__6078\ : Span4Mux_h
    port map (
            O => \N__31551\,
            I => \N__31546\
        );

    \I__6077\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31541\
        );

    \I__6076\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31541\
        );

    \I__6075\ : Odrv4
    port map (
            O => \N__31546\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__31541\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__6073\ : InMux
    port map (
            O => \N__31536\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__6072\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31530\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__31530\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__6070\ : InMux
    port map (
            O => \N__31527\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__6069\ : CascadeMux
    port map (
            O => \N__31524\,
            I => \N__31521\
        );

    \I__6068\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31518\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__31518\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__6066\ : CascadeMux
    port map (
            O => \N__31515\,
            I => \N__31512\
        );

    \I__6065\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31509\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__31509\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__6063\ : CascadeMux
    port map (
            O => \N__31506\,
            I => \N__31503\
        );

    \I__6062\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31500\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__31500\,
            I => \N__31497\
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__31497\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__6059\ : CascadeMux
    port map (
            O => \N__31494\,
            I => \N__31491\
        );

    \I__6058\ : InMux
    port map (
            O => \N__31491\,
            I => \N__31488\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__31488\,
            I => \N__31485\
        );

    \I__6056\ : Odrv4
    port map (
            O => \N__31485\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__6055\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31471\
        );

    \I__6054\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31471\
        );

    \I__6053\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31471\
        );

    \I__6052\ : InMux
    port map (
            O => \N__31479\,
            I => \N__31466\
        );

    \I__6051\ : InMux
    port map (
            O => \N__31478\,
            I => \N__31466\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__31471\,
            I => \N__31456\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__31466\,
            I => \N__31456\
        );

    \I__6048\ : InMux
    port map (
            O => \N__31465\,
            I => \N__31453\
        );

    \I__6047\ : InMux
    port map (
            O => \N__31464\,
            I => \N__31450\
        );

    \I__6046\ : InMux
    port map (
            O => \N__31463\,
            I => \N__31447\
        );

    \I__6045\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31442\
        );

    \I__6044\ : InMux
    port map (
            O => \N__31461\,
            I => \N__31442\
        );

    \I__6043\ : Span12Mux_h
    port map (
            O => \N__31456\,
            I => \N__31439\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__31453\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__31450\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__31447\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__31442\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__6038\ : Odrv12
    port map (
            O => \N__31439\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__6037\ : CascadeMux
    port map (
            O => \N__31428\,
            I => \N__31425\
        );

    \I__6036\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31422\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__31422\,
            I => \N__31419\
        );

    \I__6034\ : Odrv4
    port map (
            O => \N__31419\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__6033\ : InMux
    port map (
            O => \N__31416\,
            I => \N__31413\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__31413\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__6031\ : CascadeMux
    port map (
            O => \N__31410\,
            I => \N__31407\
        );

    \I__6030\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31404\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__31404\,
            I => \N__31401\
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__31401\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__6027\ : InMux
    port map (
            O => \N__31398\,
            I => \N__31395\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__31395\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__6025\ : CascadeMux
    port map (
            O => \N__31392\,
            I => \N__31389\
        );

    \I__6024\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31386\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__31386\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__6022\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31380\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__31380\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__6020\ : CascadeMux
    port map (
            O => \N__31377\,
            I => \N__31374\
        );

    \I__6019\ : InMux
    port map (
            O => \N__31374\,
            I => \N__31371\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__31371\,
            I => \N__31368\
        );

    \I__6017\ : Odrv4
    port map (
            O => \N__31368\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__6016\ : InMux
    port map (
            O => \N__31365\,
            I => \N__31362\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__31362\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__6014\ : CascadeMux
    port map (
            O => \N__31359\,
            I => \N__31356\
        );

    \I__6013\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31353\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__31353\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__6011\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31347\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__31347\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__6009\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31341\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__31341\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__31338\,
            I => \N__31335\
        );

    \I__6006\ : InMux
    port map (
            O => \N__31335\,
            I => \N__31332\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__31332\,
            I => \N__31329\
        );

    \I__6004\ : Odrv4
    port map (
            O => \N__31329\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__6003\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31323\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__31323\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__6001\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31317\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__31317\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__5999\ : CascadeMux
    port map (
            O => \N__31314\,
            I => \N__31311\
        );

    \I__5998\ : InMux
    port map (
            O => \N__31311\,
            I => \N__31308\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__31308\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__5996\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31302\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__31302\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__5994\ : CascadeMux
    port map (
            O => \N__31299\,
            I => \N__31296\
        );

    \I__5993\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31293\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__31293\,
            I => \N__31290\
        );

    \I__5991\ : Odrv4
    port map (
            O => \N__31290\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__5990\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31284\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__31284\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__5988\ : CascadeMux
    port map (
            O => \N__31281\,
            I => \N__31278\
        );

    \I__5987\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31275\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__31275\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__5985\ : InMux
    port map (
            O => \N__31272\,
            I => \N__31269\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__31269\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__5983\ : CascadeMux
    port map (
            O => \N__31266\,
            I => \N__31263\
        );

    \I__5982\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31260\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__31260\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__5980\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31254\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__31254\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__5978\ : CascadeMux
    port map (
            O => \N__31251\,
            I => \N__31248\
        );

    \I__5977\ : InMux
    port map (
            O => \N__31248\,
            I => \N__31245\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__31245\,
            I => \N__31242\
        );

    \I__5975\ : Odrv4
    port map (
            O => \N__31242\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__5974\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31236\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__31236\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__5972\ : CascadeMux
    port map (
            O => \N__31233\,
            I => \N__31230\
        );

    \I__5971\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31227\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__31227\,
            I => \N__31224\
        );

    \I__5969\ : Span4Mux_h
    port map (
            O => \N__31224\,
            I => \N__31221\
        );

    \I__5968\ : Odrv4
    port map (
            O => \N__31221\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__5967\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31215\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__31215\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__5965\ : InMux
    port map (
            O => \N__31212\,
            I => \N__31209\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__31209\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__31206\,
            I => \N__31203\
        );

    \I__5962\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31200\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31197\
        );

    \I__5960\ : Odrv4
    port map (
            O => \N__31197\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__5959\ : InMux
    port map (
            O => \N__31194\,
            I => \N__31191\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__31191\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__5957\ : CascadeMux
    port map (
            O => \N__31188\,
            I => \N__31183\
        );

    \I__5956\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31179\
        );

    \I__5955\ : InMux
    port map (
            O => \N__31186\,
            I => \N__31176\
        );

    \I__5954\ : InMux
    port map (
            O => \N__31183\,
            I => \N__31171\
        );

    \I__5953\ : InMux
    port map (
            O => \N__31182\,
            I => \N__31171\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__31179\,
            I => \N__31168\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__31176\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__31171\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__31168\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__5948\ : InMux
    port map (
            O => \N__31161\,
            I => \N__31155\
        );

    \I__5947\ : InMux
    port map (
            O => \N__31160\,
            I => \N__31152\
        );

    \I__5946\ : InMux
    port map (
            O => \N__31159\,
            I => \N__31147\
        );

    \I__5945\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31147\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__31155\,
            I => \N__31144\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__31152\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__31147\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__5941\ : Odrv4
    port map (
            O => \N__31144\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__5940\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31132\
        );

    \I__5939\ : InMux
    port map (
            O => \N__31136\,
            I => \N__31128\
        );

    \I__5938\ : InMux
    port map (
            O => \N__31135\,
            I => \N__31125\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__31132\,
            I => \N__31122\
        );

    \I__5936\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31119\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__31128\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__31125\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__5933\ : Odrv12
    port map (
            O => \N__31122\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__31119\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__5931\ : IoInMux
    port map (
            O => \N__31110\,
            I => \N__31107\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__31107\,
            I => \N__31104\
        );

    \I__5929\ : Span4Mux_s2_v
    port map (
            O => \N__31104\,
            I => \N__31101\
        );

    \I__5928\ : Span4Mux_v
    port map (
            O => \N__31101\,
            I => \N__31098\
        );

    \I__5927\ : Odrv4
    port map (
            O => \N__31098\,
            I => \current_shift_inst.timer_s1.N_185_i\
        );

    \I__5926\ : InMux
    port map (
            O => \N__31095\,
            I => \N__31090\
        );

    \I__5925\ : InMux
    port map (
            O => \N__31094\,
            I => \N__31087\
        );

    \I__5924\ : InMux
    port map (
            O => \N__31093\,
            I => \N__31084\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__31090\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__31087\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__31084\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__5920\ : InMux
    port map (
            O => \N__31077\,
            I => \N__31072\
        );

    \I__5919\ : InMux
    port map (
            O => \N__31076\,
            I => \N__31069\
        );

    \I__5918\ : InMux
    port map (
            O => \N__31075\,
            I => \N__31066\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__31072\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__31069\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__31066\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__5914\ : InMux
    port map (
            O => \N__31059\,
            I => \N__31056\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__31056\,
            I => \N__31053\
        );

    \I__5912\ : Span4Mux_h
    port map (
            O => \N__31053\,
            I => \N__31050\
        );

    \I__5911\ : Sp12to4
    port map (
            O => \N__31050\,
            I => \N__31047\
        );

    \I__5910\ : Odrv12
    port map (
            O => \N__31047\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__5909\ : InMux
    port map (
            O => \N__31044\,
            I => \N__31041\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__31041\,
            I => \phase_controller_inst2.start_timer_hc_RNO_0_0\
        );

    \I__5907\ : InMux
    port map (
            O => \N__31038\,
            I => \N__31035\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__31035\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__5905\ : CascadeMux
    port map (
            O => \N__31032\,
            I => \N__31029\
        );

    \I__5904\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31026\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__31026\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__5902\ : CascadeMux
    port map (
            O => \N__31023\,
            I => \N__31020\
        );

    \I__5901\ : InMux
    port map (
            O => \N__31020\,
            I => \N__31017\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__31017\,
            I => \N__31014\
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__31014\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__5898\ : InMux
    port map (
            O => \N__31011\,
            I => \N__31008\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__31008\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__5896\ : CascadeMux
    port map (
            O => \N__31005\,
            I => \N__31002\
        );

    \I__5895\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30999\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__30999\,
            I => \N__30996\
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__30996\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__5892\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30990\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__30990\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__5890\ : InMux
    port map (
            O => \N__30987\,
            I => \N__30984\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__30984\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__5888\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30978\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__30978\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__5886\ : InMux
    port map (
            O => \N__30975\,
            I => \N__30972\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__30972\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__5884\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30965\
        );

    \I__5883\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30962\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__30965\,
            I => \N__30959\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__30962\,
            I => \N__30956\
        );

    \I__5880\ : Span4Mux_h
    port map (
            O => \N__30959\,
            I => \N__30953\
        );

    \I__5879\ : Odrv12
    port map (
            O => \N__30956\,
            I => state_ns_i_a3_1
        );

    \I__5878\ : Odrv4
    port map (
            O => \N__30953\,
            I => state_ns_i_a3_1
        );

    \I__5877\ : InMux
    port map (
            O => \N__30948\,
            I => \N__30939\
        );

    \I__5876\ : InMux
    port map (
            O => \N__30947\,
            I => \N__30932\
        );

    \I__5875\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30932\
        );

    \I__5874\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30932\
        );

    \I__5873\ : InMux
    port map (
            O => \N__30944\,
            I => \N__30927\
        );

    \I__5872\ : InMux
    port map (
            O => \N__30943\,
            I => \N__30927\
        );

    \I__5871\ : CascadeMux
    port map (
            O => \N__30942\,
            I => \N__30912\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__30939\,
            I => \N__30904\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__30932\,
            I => \N__30899\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__30927\,
            I => \N__30899\
        );

    \I__5867\ : InMux
    port map (
            O => \N__30926\,
            I => \N__30884\
        );

    \I__5866\ : InMux
    port map (
            O => \N__30925\,
            I => \N__30884\
        );

    \I__5865\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30884\
        );

    \I__5864\ : InMux
    port map (
            O => \N__30923\,
            I => \N__30884\
        );

    \I__5863\ : InMux
    port map (
            O => \N__30922\,
            I => \N__30884\
        );

    \I__5862\ : InMux
    port map (
            O => \N__30921\,
            I => \N__30884\
        );

    \I__5861\ : InMux
    port map (
            O => \N__30920\,
            I => \N__30884\
        );

    \I__5860\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30871\
        );

    \I__5859\ : InMux
    port map (
            O => \N__30918\,
            I => \N__30871\
        );

    \I__5858\ : InMux
    port map (
            O => \N__30917\,
            I => \N__30871\
        );

    \I__5857\ : InMux
    port map (
            O => \N__30916\,
            I => \N__30871\
        );

    \I__5856\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30871\
        );

    \I__5855\ : InMux
    port map (
            O => \N__30912\,
            I => \N__30871\
        );

    \I__5854\ : InMux
    port map (
            O => \N__30911\,
            I => \N__30860\
        );

    \I__5853\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30860\
        );

    \I__5852\ : InMux
    port map (
            O => \N__30909\,
            I => \N__30860\
        );

    \I__5851\ : InMux
    port map (
            O => \N__30908\,
            I => \N__30860\
        );

    \I__5850\ : InMux
    port map (
            O => \N__30907\,
            I => \N__30860\
        );

    \I__5849\ : Span4Mux_v
    port map (
            O => \N__30904\,
            I => \N__30856\
        );

    \I__5848\ : Span4Mux_v
    port map (
            O => \N__30899\,
            I => \N__30853\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__30884\,
            I => \N__30846\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__30871\,
            I => \N__30846\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__30860\,
            I => \N__30846\
        );

    \I__5844\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30843\
        );

    \I__5843\ : Odrv4
    port map (
            O => \N__30856\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5842\ : Odrv4
    port map (
            O => \N__30853\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5841\ : Odrv4
    port map (
            O => \N__30846\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__30843\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5839\ : InMux
    port map (
            O => \N__30834\,
            I => \N__30831\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__30831\,
            I => \N__30826\
        );

    \I__5837\ : InMux
    port map (
            O => \N__30830\,
            I => \N__30823\
        );

    \I__5836\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30820\
        );

    \I__5835\ : Span4Mux_v
    port map (
            O => \N__30826\,
            I => \N__30817\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__30823\,
            I => \N__30812\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__30820\,
            I => \N__30812\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__30817\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__5831\ : Odrv4
    port map (
            O => \N__30812\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__5830\ : InMux
    port map (
            O => \N__30807\,
            I => \N__30804\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__30804\,
            I => \N__30801\
        );

    \I__5828\ : Span4Mux_h
    port map (
            O => \N__30801\,
            I => \N__30798\
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__30798\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__5826\ : InMux
    port map (
            O => \N__30795\,
            I => \N__30792\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__30792\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__5824\ : InMux
    port map (
            O => \N__30789\,
            I => \N__30786\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__30786\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__5822\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30780\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__30780\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__5820\ : InMux
    port map (
            O => \N__30777\,
            I => \N__30774\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__30774\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__5818\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30768\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__30768\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__5816\ : InMux
    port map (
            O => \N__30765\,
            I => \N__30762\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__30762\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__5814\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30756\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__30756\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__5812\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30750\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__30750\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__5810\ : InMux
    port map (
            O => \N__30747\,
            I => \N__30744\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__30744\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__5808\ : InMux
    port map (
            O => \N__30741\,
            I => \N__30738\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__30738\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__5806\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30732\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__30732\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__5804\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30726\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__30726\,
            I => \N__30723\
        );

    \I__5802\ : Span4Mux_h
    port map (
            O => \N__30723\,
            I => \N__30718\
        );

    \I__5801\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30715\
        );

    \I__5800\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30712\
        );

    \I__5799\ : Odrv4
    port map (
            O => \N__30718\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__30715\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__30712\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__5796\ : InMux
    port map (
            O => \N__30705\,
            I => \N__30702\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__30702\,
            I => \N__30699\
        );

    \I__5794\ : Span4Mux_v
    port map (
            O => \N__30699\,
            I => \N__30696\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__30696\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__30693\,
            I => \N__30683\
        );

    \I__5791\ : CascadeMux
    port map (
            O => \N__30692\,
            I => \N__30680\
        );

    \I__5790\ : CascadeMux
    port map (
            O => \N__30691\,
            I => \N__30661\
        );

    \I__5789\ : CascadeMux
    port map (
            O => \N__30690\,
            I => \N__30658\
        );

    \I__5788\ : CascadeMux
    port map (
            O => \N__30689\,
            I => \N__30655\
        );

    \I__5787\ : CascadeMux
    port map (
            O => \N__30688\,
            I => \N__30652\
        );

    \I__5786\ : CascadeMux
    port map (
            O => \N__30687\,
            I => \N__30649\
        );

    \I__5785\ : CascadeMux
    port map (
            O => \N__30686\,
            I => \N__30644\
        );

    \I__5784\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30641\
        );

    \I__5783\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30638\
        );

    \I__5782\ : InMux
    port map (
            O => \N__30679\,
            I => \N__30635\
        );

    \I__5781\ : CascadeMux
    port map (
            O => \N__30678\,
            I => \N__30632\
        );

    \I__5780\ : CascadeMux
    port map (
            O => \N__30677\,
            I => \N__30629\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__30676\,
            I => \N__30626\
        );

    \I__5778\ : CascadeMux
    port map (
            O => \N__30675\,
            I => \N__30616\
        );

    \I__5777\ : CascadeMux
    port map (
            O => \N__30674\,
            I => \N__30611\
        );

    \I__5776\ : InMux
    port map (
            O => \N__30673\,
            I => \N__30607\
        );

    \I__5775\ : CascadeMux
    port map (
            O => \N__30672\,
            I => \N__30599\
        );

    \I__5774\ : CascadeMux
    port map (
            O => \N__30671\,
            I => \N__30592\
        );

    \I__5773\ : CascadeMux
    port map (
            O => \N__30670\,
            I => \N__30589\
        );

    \I__5772\ : CascadeMux
    port map (
            O => \N__30669\,
            I => \N__30585\
        );

    \I__5771\ : CascadeMux
    port map (
            O => \N__30668\,
            I => \N__30582\
        );

    \I__5770\ : CascadeMux
    port map (
            O => \N__30667\,
            I => \N__30579\
        );

    \I__5769\ : CascadeMux
    port map (
            O => \N__30666\,
            I => \N__30576\
        );

    \I__5768\ : CascadeMux
    port map (
            O => \N__30665\,
            I => \N__30573\
        );

    \I__5767\ : CascadeMux
    port map (
            O => \N__30664\,
            I => \N__30570\
        );

    \I__5766\ : InMux
    port map (
            O => \N__30661\,
            I => \N__30563\
        );

    \I__5765\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30560\
        );

    \I__5764\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30555\
        );

    \I__5763\ : InMux
    port map (
            O => \N__30652\,
            I => \N__30555\
        );

    \I__5762\ : InMux
    port map (
            O => \N__30649\,
            I => \N__30548\
        );

    \I__5761\ : InMux
    port map (
            O => \N__30648\,
            I => \N__30548\
        );

    \I__5760\ : InMux
    port map (
            O => \N__30647\,
            I => \N__30548\
        );

    \I__5759\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30545\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__30641\,
            I => \N__30538\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__30638\,
            I => \N__30538\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__30635\,
            I => \N__30538\
        );

    \I__5755\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30531\
        );

    \I__5754\ : InMux
    port map (
            O => \N__30629\,
            I => \N__30531\
        );

    \I__5753\ : InMux
    port map (
            O => \N__30626\,
            I => \N__30531\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__30625\,
            I => \N__30528\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__30624\,
            I => \N__30525\
        );

    \I__5750\ : CascadeMux
    port map (
            O => \N__30623\,
            I => \N__30522\
        );

    \I__5749\ : CascadeMux
    port map (
            O => \N__30622\,
            I => \N__30519\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__30621\,
            I => \N__30516\
        );

    \I__5747\ : CascadeMux
    port map (
            O => \N__30620\,
            I => \N__30513\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__30619\,
            I => \N__30510\
        );

    \I__5745\ : InMux
    port map (
            O => \N__30616\,
            I => \N__30507\
        );

    \I__5744\ : InMux
    port map (
            O => \N__30615\,
            I => \N__30504\
        );

    \I__5743\ : InMux
    port map (
            O => \N__30614\,
            I => \N__30501\
        );

    \I__5742\ : InMux
    port map (
            O => \N__30611\,
            I => \N__30498\
        );

    \I__5741\ : CascadeMux
    port map (
            O => \N__30610\,
            I => \N__30495\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__30607\,
            I => \N__30489\
        );

    \I__5739\ : CascadeMux
    port map (
            O => \N__30606\,
            I => \N__30486\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__30605\,
            I => \N__30483\
        );

    \I__5737\ : CascadeMux
    port map (
            O => \N__30604\,
            I => \N__30479\
        );

    \I__5736\ : CascadeMux
    port map (
            O => \N__30603\,
            I => \N__30476\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__30602\,
            I => \N__30472\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30461\
        );

    \I__5733\ : CascadeMux
    port map (
            O => \N__30598\,
            I => \N__30455\
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__30597\,
            I => \N__30452\
        );

    \I__5731\ : CascadeMux
    port map (
            O => \N__30596\,
            I => \N__30449\
        );

    \I__5730\ : CascadeMux
    port map (
            O => \N__30595\,
            I => \N__30445\
        );

    \I__5729\ : InMux
    port map (
            O => \N__30592\,
            I => \N__30421\
        );

    \I__5728\ : InMux
    port map (
            O => \N__30589\,
            I => \N__30412\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30588\,
            I => \N__30412\
        );

    \I__5726\ : InMux
    port map (
            O => \N__30585\,
            I => \N__30412\
        );

    \I__5725\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30412\
        );

    \I__5724\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30403\
        );

    \I__5723\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30403\
        );

    \I__5722\ : InMux
    port map (
            O => \N__30573\,
            I => \N__30403\
        );

    \I__5721\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30403\
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__30569\,
            I => \N__30400\
        );

    \I__5719\ : CascadeMux
    port map (
            O => \N__30568\,
            I => \N__30397\
        );

    \I__5718\ : CascadeMux
    port map (
            O => \N__30567\,
            I => \N__30394\
        );

    \I__5717\ : CascadeMux
    port map (
            O => \N__30566\,
            I => \N__30390\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__30563\,
            I => \N__30375\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__30560\,
            I => \N__30375\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__30555\,
            I => \N__30375\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__30548\,
            I => \N__30375\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__30545\,
            I => \N__30375\
        );

    \I__5711\ : Span4Mux_v
    port map (
            O => \N__30538\,
            I => \N__30375\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__30531\,
            I => \N__30375\
        );

    \I__5709\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30366\
        );

    \I__5708\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30366\
        );

    \I__5707\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30366\
        );

    \I__5706\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30366\
        );

    \I__5705\ : InMux
    port map (
            O => \N__30516\,
            I => \N__30359\
        );

    \I__5704\ : InMux
    port map (
            O => \N__30513\,
            I => \N__30359\
        );

    \I__5703\ : InMux
    port map (
            O => \N__30510\,
            I => \N__30359\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__30507\,
            I => \N__30354\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__30504\,
            I => \N__30354\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__30501\,
            I => \N__30351\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__30498\,
            I => \N__30343\
        );

    \I__5698\ : InMux
    port map (
            O => \N__30495\,
            I => \N__30338\
        );

    \I__5697\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30338\
        );

    \I__5696\ : CascadeMux
    port map (
            O => \N__30493\,
            I => \N__30335\
        );

    \I__5695\ : CascadeMux
    port map (
            O => \N__30492\,
            I => \N__30329\
        );

    \I__5694\ : Span4Mux_h
    port map (
            O => \N__30489\,
            I => \N__30326\
        );

    \I__5693\ : InMux
    port map (
            O => \N__30486\,
            I => \N__30323\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30483\,
            I => \N__30316\
        );

    \I__5691\ : InMux
    port map (
            O => \N__30482\,
            I => \N__30316\
        );

    \I__5690\ : InMux
    port map (
            O => \N__30479\,
            I => \N__30316\
        );

    \I__5689\ : InMux
    port map (
            O => \N__30476\,
            I => \N__30309\
        );

    \I__5688\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30309\
        );

    \I__5687\ : InMux
    port map (
            O => \N__30472\,
            I => \N__30309\
        );

    \I__5686\ : InMux
    port map (
            O => \N__30471\,
            I => \N__30304\
        );

    \I__5685\ : InMux
    port map (
            O => \N__30470\,
            I => \N__30304\
        );

    \I__5684\ : CascadeMux
    port map (
            O => \N__30469\,
            I => \N__30301\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__30468\,
            I => \N__30298\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__30467\,
            I => \N__30295\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__30466\,
            I => \N__30292\
        );

    \I__5680\ : CascadeMux
    port map (
            O => \N__30465\,
            I => \N__30289\
        );

    \I__5679\ : CascadeMux
    port map (
            O => \N__30464\,
            I => \N__30286\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__30461\,
            I => \N__30269\
        );

    \I__5677\ : CascadeMux
    port map (
            O => \N__30460\,
            I => \N__30265\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__30459\,
            I => \N__30262\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__30458\,
            I => \N__30259\
        );

    \I__5674\ : InMux
    port map (
            O => \N__30455\,
            I => \N__30248\
        );

    \I__5673\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30248\
        );

    \I__5672\ : InMux
    port map (
            O => \N__30449\,
            I => \N__30248\
        );

    \I__5671\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30248\
        );

    \I__5670\ : InMux
    port map (
            O => \N__30445\,
            I => \N__30248\
        );

    \I__5669\ : CascadeMux
    port map (
            O => \N__30444\,
            I => \N__30245\
        );

    \I__5668\ : CascadeMux
    port map (
            O => \N__30443\,
            I => \N__30242\
        );

    \I__5667\ : CascadeMux
    port map (
            O => \N__30442\,
            I => \N__30239\
        );

    \I__5666\ : CascadeMux
    port map (
            O => \N__30441\,
            I => \N__30235\
        );

    \I__5665\ : CascadeMux
    port map (
            O => \N__30440\,
            I => \N__30232\
        );

    \I__5664\ : CascadeMux
    port map (
            O => \N__30439\,
            I => \N__30229\
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__30438\,
            I => \N__30226\
        );

    \I__5662\ : CascadeMux
    port map (
            O => \N__30437\,
            I => \N__30223\
        );

    \I__5661\ : CascadeMux
    port map (
            O => \N__30436\,
            I => \N__30220\
        );

    \I__5660\ : CascadeMux
    port map (
            O => \N__30435\,
            I => \N__30217\
        );

    \I__5659\ : CascadeMux
    port map (
            O => \N__30434\,
            I => \N__30214\
        );

    \I__5658\ : CascadeMux
    port map (
            O => \N__30433\,
            I => \N__30211\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__30432\,
            I => \N__30208\
        );

    \I__5656\ : CascadeMux
    port map (
            O => \N__30431\,
            I => \N__30205\
        );

    \I__5655\ : CascadeMux
    port map (
            O => \N__30430\,
            I => \N__30202\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__30429\,
            I => \N__30199\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__30428\,
            I => \N__30196\
        );

    \I__5652\ : CascadeMux
    port map (
            O => \N__30427\,
            I => \N__30193\
        );

    \I__5651\ : CascadeMux
    port map (
            O => \N__30426\,
            I => \N__30190\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__30425\,
            I => \N__30187\
        );

    \I__5649\ : CascadeMux
    port map (
            O => \N__30424\,
            I => \N__30183\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__30421\,
            I => \N__30176\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__30412\,
            I => \N__30176\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__30403\,
            I => \N__30176\
        );

    \I__5645\ : InMux
    port map (
            O => \N__30400\,
            I => \N__30171\
        );

    \I__5644\ : InMux
    port map (
            O => \N__30397\,
            I => \N__30171\
        );

    \I__5643\ : InMux
    port map (
            O => \N__30394\,
            I => \N__30164\
        );

    \I__5642\ : InMux
    port map (
            O => \N__30393\,
            I => \N__30164\
        );

    \I__5641\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30164\
        );

    \I__5640\ : Span4Mux_v
    port map (
            O => \N__30375\,
            I => \N__30157\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__30366\,
            I => \N__30157\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__30359\,
            I => \N__30157\
        );

    \I__5637\ : Span4Mux_h
    port map (
            O => \N__30354\,
            I => \N__30152\
        );

    \I__5636\ : Span4Mux_v
    port map (
            O => \N__30351\,
            I => \N__30152\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__30350\,
            I => \N__30149\
        );

    \I__5634\ : CascadeMux
    port map (
            O => \N__30349\,
            I => \N__30146\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__30348\,
            I => \N__30142\
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__30347\,
            I => \N__30138\
        );

    \I__5631\ : CascadeMux
    port map (
            O => \N__30346\,
            I => \N__30135\
        );

    \I__5630\ : Span4Mux_v
    port map (
            O => \N__30343\,
            I => \N__30130\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__30338\,
            I => \N__30130\
        );

    \I__5628\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30127\
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__30334\,
            I => \N__30124\
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__30333\,
            I => \N__30121\
        );

    \I__5625\ : InMux
    port map (
            O => \N__30332\,
            I => \N__30118\
        );

    \I__5624\ : InMux
    port map (
            O => \N__30329\,
            I => \N__30115\
        );

    \I__5623\ : Span4Mux_v
    port map (
            O => \N__30326\,
            I => \N__30104\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__30323\,
            I => \N__30104\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__30316\,
            I => \N__30104\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__30309\,
            I => \N__30104\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__30304\,
            I => \N__30104\
        );

    \I__5618\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30099\
        );

    \I__5617\ : InMux
    port map (
            O => \N__30298\,
            I => \N__30099\
        );

    \I__5616\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30090\
        );

    \I__5615\ : InMux
    port map (
            O => \N__30292\,
            I => \N__30090\
        );

    \I__5614\ : InMux
    port map (
            O => \N__30289\,
            I => \N__30090\
        );

    \I__5613\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30090\
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__30285\,
            I => \N__30087\
        );

    \I__5611\ : CascadeMux
    port map (
            O => \N__30284\,
            I => \N__30084\
        );

    \I__5610\ : CascadeMux
    port map (
            O => \N__30283\,
            I => \N__30081\
        );

    \I__5609\ : CascadeMux
    port map (
            O => \N__30282\,
            I => \N__30078\
        );

    \I__5608\ : CascadeMux
    port map (
            O => \N__30281\,
            I => \N__30075\
        );

    \I__5607\ : CascadeMux
    port map (
            O => \N__30280\,
            I => \N__30072\
        );

    \I__5606\ : CascadeMux
    port map (
            O => \N__30279\,
            I => \N__30069\
        );

    \I__5605\ : CascadeMux
    port map (
            O => \N__30278\,
            I => \N__30066\
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__30277\,
            I => \N__30063\
        );

    \I__5603\ : CascadeMux
    port map (
            O => \N__30276\,
            I => \N__30060\
        );

    \I__5602\ : CascadeMux
    port map (
            O => \N__30275\,
            I => \N__30057\
        );

    \I__5601\ : CascadeMux
    port map (
            O => \N__30274\,
            I => \N__30054\
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__30273\,
            I => \N__30051\
        );

    \I__5599\ : CascadeMux
    port map (
            O => \N__30272\,
            I => \N__30048\
        );

    \I__5598\ : Span4Mux_v
    port map (
            O => \N__30269\,
            I => \N__30045\
        );

    \I__5597\ : InMux
    port map (
            O => \N__30268\,
            I => \N__30036\
        );

    \I__5596\ : InMux
    port map (
            O => \N__30265\,
            I => \N__30036\
        );

    \I__5595\ : InMux
    port map (
            O => \N__30262\,
            I => \N__30036\
        );

    \I__5594\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30036\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__30248\,
            I => \N__30033\
        );

    \I__5592\ : InMux
    port map (
            O => \N__30245\,
            I => \N__30024\
        );

    \I__5591\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30024\
        );

    \I__5590\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30024\
        );

    \I__5589\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30024\
        );

    \I__5588\ : InMux
    port map (
            O => \N__30235\,
            I => \N__30015\
        );

    \I__5587\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30015\
        );

    \I__5586\ : InMux
    port map (
            O => \N__30229\,
            I => \N__30015\
        );

    \I__5585\ : InMux
    port map (
            O => \N__30226\,
            I => \N__30015\
        );

    \I__5584\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30006\
        );

    \I__5583\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30006\
        );

    \I__5582\ : InMux
    port map (
            O => \N__30217\,
            I => \N__30006\
        );

    \I__5581\ : InMux
    port map (
            O => \N__30214\,
            I => \N__30006\
        );

    \I__5580\ : InMux
    port map (
            O => \N__30211\,
            I => \N__29997\
        );

    \I__5579\ : InMux
    port map (
            O => \N__30208\,
            I => \N__29997\
        );

    \I__5578\ : InMux
    port map (
            O => \N__30205\,
            I => \N__29997\
        );

    \I__5577\ : InMux
    port map (
            O => \N__30202\,
            I => \N__29997\
        );

    \I__5576\ : InMux
    port map (
            O => \N__30199\,
            I => \N__29988\
        );

    \I__5575\ : InMux
    port map (
            O => \N__30196\,
            I => \N__29988\
        );

    \I__5574\ : InMux
    port map (
            O => \N__30193\,
            I => \N__29988\
        );

    \I__5573\ : InMux
    port map (
            O => \N__30190\,
            I => \N__29988\
        );

    \I__5572\ : InMux
    port map (
            O => \N__30187\,
            I => \N__29981\
        );

    \I__5571\ : InMux
    port map (
            O => \N__30186\,
            I => \N__29981\
        );

    \I__5570\ : InMux
    port map (
            O => \N__30183\,
            I => \N__29981\
        );

    \I__5569\ : Span4Mux_v
    port map (
            O => \N__30176\,
            I => \N__29974\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__30171\,
            I => \N__29974\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__30164\,
            I => \N__29974\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__30157\,
            I => \N__29969\
        );

    \I__5565\ : Span4Mux_h
    port map (
            O => \N__30152\,
            I => \N__29969\
        );

    \I__5564\ : InMux
    port map (
            O => \N__30149\,
            I => \N__29960\
        );

    \I__5563\ : InMux
    port map (
            O => \N__30146\,
            I => \N__29960\
        );

    \I__5562\ : InMux
    port map (
            O => \N__30145\,
            I => \N__29960\
        );

    \I__5561\ : InMux
    port map (
            O => \N__30142\,
            I => \N__29960\
        );

    \I__5560\ : InMux
    port map (
            O => \N__30141\,
            I => \N__29953\
        );

    \I__5559\ : InMux
    port map (
            O => \N__30138\,
            I => \N__29953\
        );

    \I__5558\ : InMux
    port map (
            O => \N__30135\,
            I => \N__29953\
        );

    \I__5557\ : Span4Mux_h
    port map (
            O => \N__30130\,
            I => \N__29948\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__30127\,
            I => \N__29948\
        );

    \I__5555\ : InMux
    port map (
            O => \N__30124\,
            I => \N__29945\
        );

    \I__5554\ : InMux
    port map (
            O => \N__30121\,
            I => \N__29942\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__30118\,
            I => \N__29937\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__30115\,
            I => \N__29937\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__30104\,
            I => \N__29930\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__30099\,
            I => \N__29930\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__30090\,
            I => \N__29930\
        );

    \I__5548\ : InMux
    port map (
            O => \N__30087\,
            I => \N__29921\
        );

    \I__5547\ : InMux
    port map (
            O => \N__30084\,
            I => \N__29921\
        );

    \I__5546\ : InMux
    port map (
            O => \N__30081\,
            I => \N__29921\
        );

    \I__5545\ : InMux
    port map (
            O => \N__30078\,
            I => \N__29921\
        );

    \I__5544\ : InMux
    port map (
            O => \N__30075\,
            I => \N__29912\
        );

    \I__5543\ : InMux
    port map (
            O => \N__30072\,
            I => \N__29912\
        );

    \I__5542\ : InMux
    port map (
            O => \N__30069\,
            I => \N__29912\
        );

    \I__5541\ : InMux
    port map (
            O => \N__30066\,
            I => \N__29912\
        );

    \I__5540\ : InMux
    port map (
            O => \N__30063\,
            I => \N__29903\
        );

    \I__5539\ : InMux
    port map (
            O => \N__30060\,
            I => \N__29903\
        );

    \I__5538\ : InMux
    port map (
            O => \N__30057\,
            I => \N__29903\
        );

    \I__5537\ : InMux
    port map (
            O => \N__30054\,
            I => \N__29903\
        );

    \I__5536\ : InMux
    port map (
            O => \N__30051\,
            I => \N__29898\
        );

    \I__5535\ : InMux
    port map (
            O => \N__30048\,
            I => \N__29898\
        );

    \I__5534\ : Span4Mux_v
    port map (
            O => \N__30045\,
            I => \N__29879\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__30036\,
            I => \N__29879\
        );

    \I__5532\ : Span4Mux_h
    port map (
            O => \N__30033\,
            I => \N__29879\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__30024\,
            I => \N__29879\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__30015\,
            I => \N__29879\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__30006\,
            I => \N__29879\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__29997\,
            I => \N__29879\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__29988\,
            I => \N__29879\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__29981\,
            I => \N__29879\
        );

    \I__5525\ : Span4Mux_h
    port map (
            O => \N__29974\,
            I => \N__29870\
        );

    \I__5524\ : Span4Mux_v
    port map (
            O => \N__29969\,
            I => \N__29870\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__29960\,
            I => \N__29870\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__29953\,
            I => \N__29870\
        );

    \I__5521\ : Odrv4
    port map (
            O => \N__29948\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__29945\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__29942\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5518\ : Odrv12
    port map (
            O => \N__29937\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5517\ : Odrv4
    port map (
            O => \N__29930\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__29921\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__29912\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__29903\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__29898\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__29879\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5511\ : Odrv4
    port map (
            O => \N__29870\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__29847\,
            I => \N__29838\
        );

    \I__5509\ : CascadeMux
    port map (
            O => \N__29846\,
            I => \N__29829\
        );

    \I__5508\ : InMux
    port map (
            O => \N__29845\,
            I => \N__29825\
        );

    \I__5507\ : CascadeMux
    port map (
            O => \N__29844\,
            I => \N__29804\
        );

    \I__5506\ : InMux
    port map (
            O => \N__29843\,
            I => \N__29796\
        );

    \I__5505\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29793\
        );

    \I__5504\ : InMux
    port map (
            O => \N__29841\,
            I => \N__29784\
        );

    \I__5503\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29784\
        );

    \I__5502\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29784\
        );

    \I__5501\ : InMux
    port map (
            O => \N__29836\,
            I => \N__29784\
        );

    \I__5500\ : InMux
    port map (
            O => \N__29835\,
            I => \N__29777\
        );

    \I__5499\ : InMux
    port map (
            O => \N__29834\,
            I => \N__29777\
        );

    \I__5498\ : InMux
    port map (
            O => \N__29833\,
            I => \N__29768\
        );

    \I__5497\ : InMux
    port map (
            O => \N__29832\,
            I => \N__29768\
        );

    \I__5496\ : InMux
    port map (
            O => \N__29829\,
            I => \N__29768\
        );

    \I__5495\ : InMux
    port map (
            O => \N__29828\,
            I => \N__29768\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__29825\,
            I => \N__29764\
        );

    \I__5493\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29761\
        );

    \I__5492\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29756\
        );

    \I__5491\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29756\
        );

    \I__5490\ : InMux
    port map (
            O => \N__29821\,
            I => \N__29747\
        );

    \I__5489\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29747\
        );

    \I__5488\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29747\
        );

    \I__5487\ : InMux
    port map (
            O => \N__29818\,
            I => \N__29747\
        );

    \I__5486\ : InMux
    port map (
            O => \N__29817\,
            I => \N__29740\
        );

    \I__5485\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29740\
        );

    \I__5484\ : InMux
    port map (
            O => \N__29815\,
            I => \N__29740\
        );

    \I__5483\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29737\
        );

    \I__5482\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29722\
        );

    \I__5481\ : InMux
    port map (
            O => \N__29812\,
            I => \N__29722\
        );

    \I__5480\ : InMux
    port map (
            O => \N__29811\,
            I => \N__29722\
        );

    \I__5479\ : InMux
    port map (
            O => \N__29810\,
            I => \N__29722\
        );

    \I__5478\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29719\
        );

    \I__5477\ : InMux
    port map (
            O => \N__29808\,
            I => \N__29710\
        );

    \I__5476\ : InMux
    port map (
            O => \N__29807\,
            I => \N__29710\
        );

    \I__5475\ : InMux
    port map (
            O => \N__29804\,
            I => \N__29710\
        );

    \I__5474\ : InMux
    port map (
            O => \N__29803\,
            I => \N__29710\
        );

    \I__5473\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29693\
        );

    \I__5472\ : InMux
    port map (
            O => \N__29801\,
            I => \N__29687\
        );

    \I__5471\ : InMux
    port map (
            O => \N__29800\,
            I => \N__29682\
        );

    \I__5470\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29682\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__29796\,
            I => \N__29675\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__29793\,
            I => \N__29675\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__29784\,
            I => \N__29675\
        );

    \I__5466\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29670\
        );

    \I__5465\ : InMux
    port map (
            O => \N__29782\,
            I => \N__29670\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__29777\,
            I => \N__29665\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__29768\,
            I => \N__29665\
        );

    \I__5462\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29662\
        );

    \I__5461\ : Span4Mux_h
    port map (
            O => \N__29764\,
            I => \N__29651\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__29761\,
            I => \N__29651\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__29756\,
            I => \N__29651\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__29747\,
            I => \N__29651\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__29740\,
            I => \N__29651\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__29737\,
            I => \N__29648\
        );

    \I__5455\ : InMux
    port map (
            O => \N__29736\,
            I => \N__29639\
        );

    \I__5454\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29639\
        );

    \I__5453\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29639\
        );

    \I__5452\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29639\
        );

    \I__5451\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29634\
        );

    \I__5450\ : InMux
    port map (
            O => \N__29731\,
            I => \N__29634\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__29722\,
            I => \N__29631\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__29719\,
            I => \N__29625\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__29710\,
            I => \N__29625\
        );

    \I__5446\ : InMux
    port map (
            O => \N__29709\,
            I => \N__29618\
        );

    \I__5445\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29618\
        );

    \I__5444\ : InMux
    port map (
            O => \N__29707\,
            I => \N__29618\
        );

    \I__5443\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29609\
        );

    \I__5442\ : InMux
    port map (
            O => \N__29705\,
            I => \N__29609\
        );

    \I__5441\ : InMux
    port map (
            O => \N__29704\,
            I => \N__29609\
        );

    \I__5440\ : InMux
    port map (
            O => \N__29703\,
            I => \N__29609\
        );

    \I__5439\ : InMux
    port map (
            O => \N__29702\,
            I => \N__29600\
        );

    \I__5438\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29600\
        );

    \I__5437\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29600\
        );

    \I__5436\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29600\
        );

    \I__5435\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29595\
        );

    \I__5434\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29595\
        );

    \I__5433\ : CascadeMux
    port map (
            O => \N__29696\,
            I => \N__29592\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__29693\,
            I => \N__29588\
        );

    \I__5431\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29585\
        );

    \I__5430\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29582\
        );

    \I__5429\ : InMux
    port map (
            O => \N__29690\,
            I => \N__29576\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__29687\,
            I => \N__29573\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__29682\,
            I => \N__29570\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__29675\,
            I => \N__29563\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__29670\,
            I => \N__29563\
        );

    \I__5424\ : Span4Mux_v
    port map (
            O => \N__29665\,
            I => \N__29563\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__29662\,
            I => \N__29550\
        );

    \I__5422\ : Span4Mux_v
    port map (
            O => \N__29651\,
            I => \N__29550\
        );

    \I__5421\ : Span4Mux_h
    port map (
            O => \N__29648\,
            I => \N__29550\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__29639\,
            I => \N__29550\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__29634\,
            I => \N__29550\
        );

    \I__5418\ : Span4Mux_h
    port map (
            O => \N__29631\,
            I => \N__29550\
        );

    \I__5417\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29547\
        );

    \I__5416\ : Span4Mux_v
    port map (
            O => \N__29625\,
            I => \N__29536\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__29618\,
            I => \N__29536\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__29609\,
            I => \N__29536\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__29600\,
            I => \N__29536\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__29595\,
            I => \N__29536\
        );

    \I__5411\ : InMux
    port map (
            O => \N__29592\,
            I => \N__29529\
        );

    \I__5410\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29529\
        );

    \I__5409\ : Span4Mux_h
    port map (
            O => \N__29588\,
            I => \N__29524\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__29585\,
            I => \N__29524\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__29582\,
            I => \N__29521\
        );

    \I__5406\ : InMux
    port map (
            O => \N__29581\,
            I => \N__29516\
        );

    \I__5405\ : InMux
    port map (
            O => \N__29580\,
            I => \N__29516\
        );

    \I__5404\ : InMux
    port map (
            O => \N__29579\,
            I => \N__29513\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__29576\,
            I => \N__29504\
        );

    \I__5402\ : Span4Mux_v
    port map (
            O => \N__29573\,
            I => \N__29504\
        );

    \I__5401\ : Span4Mux_v
    port map (
            O => \N__29570\,
            I => \N__29504\
        );

    \I__5400\ : Span4Mux_v
    port map (
            O => \N__29563\,
            I => \N__29504\
        );

    \I__5399\ : Span4Mux_v
    port map (
            O => \N__29550\,
            I => \N__29501\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__29547\,
            I => \N__29496\
        );

    \I__5397\ : Span4Mux_v
    port map (
            O => \N__29536\,
            I => \N__29496\
        );

    \I__5396\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29491\
        );

    \I__5395\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29491\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__29529\,
            I => \N__29484\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__29524\,
            I => \N__29484\
        );

    \I__5392\ : Span4Mux_h
    port map (
            O => \N__29521\,
            I => \N__29484\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__29516\,
            I => \N__29481\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__29513\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5389\ : Odrv4
    port map (
            O => \N__29504\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__29501\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__29496\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__29491\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5385\ : Odrv4
    port map (
            O => \N__29484\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5384\ : Odrv4
    port map (
            O => \N__29481\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5383\ : InMux
    port map (
            O => \N__29466\,
            I => \N__29461\
        );

    \I__5382\ : InMux
    port map (
            O => \N__29465\,
            I => \N__29458\
        );

    \I__5381\ : InMux
    port map (
            O => \N__29464\,
            I => \N__29455\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__29461\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__29458\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__29455\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__5377\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29445\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__29445\,
            I => \N__29442\
        );

    \I__5375\ : Span4Mux_h
    port map (
            O => \N__29442\,
            I => \N__29439\
        );

    \I__5374\ : Span4Mux_v
    port map (
            O => \N__29439\,
            I => \N__29436\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__29436\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\
        );

    \I__5372\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29430\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__29430\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__5370\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29424\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__29424\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__5368\ : InMux
    port map (
            O => \N__29421\,
            I => \N__29418\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__29418\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__5366\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29412\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__29412\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__5364\ : InMux
    port map (
            O => \N__29409\,
            I => \N__29406\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__29406\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__5362\ : InMux
    port map (
            O => \N__29403\,
            I => \N__29400\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__29400\,
            I => \N__29396\
        );

    \I__5360\ : InMux
    port map (
            O => \N__29399\,
            I => \N__29393\
        );

    \I__5359\ : Span4Mux_s1_v
    port map (
            O => \N__29396\,
            I => \N__29387\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__29393\,
            I => \N__29387\
        );

    \I__5357\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29384\
        );

    \I__5356\ : Span4Mux_v
    port map (
            O => \N__29387\,
            I => \N__29380\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__29384\,
            I => \N__29377\
        );

    \I__5354\ : InMux
    port map (
            O => \N__29383\,
            I => \N__29374\
        );

    \I__5353\ : Span4Mux_h
    port map (
            O => \N__29380\,
            I => \N__29370\
        );

    \I__5352\ : Span4Mux_h
    port map (
            O => \N__29377\,
            I => \N__29365\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__29374\,
            I => \N__29365\
        );

    \I__5350\ : InMux
    port map (
            O => \N__29373\,
            I => \N__29362\
        );

    \I__5349\ : Sp12to4
    port map (
            O => \N__29370\,
            I => \N__29359\
        );

    \I__5348\ : Span4Mux_v
    port map (
            O => \N__29365\,
            I => \N__29356\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__29362\,
            I => \N__29353\
        );

    \I__5346\ : Span12Mux_v
    port map (
            O => \N__29359\,
            I => \N__29350\
        );

    \I__5345\ : Sp12to4
    port map (
            O => \N__29356\,
            I => \N__29347\
        );

    \I__5344\ : Span4Mux_v
    port map (
            O => \N__29353\,
            I => \N__29344\
        );

    \I__5343\ : Span12Mux_v
    port map (
            O => \N__29350\,
            I => \N__29341\
        );

    \I__5342\ : Span12Mux_h
    port map (
            O => \N__29347\,
            I => \N__29338\
        );

    \I__5341\ : Sp12to4
    port map (
            O => \N__29344\,
            I => \N__29335\
        );

    \I__5340\ : Span12Mux_h
    port map (
            O => \N__29341\,
            I => \N__29330\
        );

    \I__5339\ : Span12Mux_v
    port map (
            O => \N__29338\,
            I => \N__29330\
        );

    \I__5338\ : Span12Mux_h
    port map (
            O => \N__29335\,
            I => \N__29327\
        );

    \I__5337\ : Odrv12
    port map (
            O => \N__29330\,
            I => start_stop_c
        );

    \I__5336\ : Odrv12
    port map (
            O => \N__29327\,
            I => start_stop_c
        );

    \I__5335\ : CEMux
    port map (
            O => \N__29322\,
            I => \N__29317\
        );

    \I__5334\ : CEMux
    port map (
            O => \N__29321\,
            I => \N__29313\
        );

    \I__5333\ : CEMux
    port map (
            O => \N__29320\,
            I => \N__29310\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__29317\,
            I => \N__29307\
        );

    \I__5331\ : CEMux
    port map (
            O => \N__29316\,
            I => \N__29304\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__29313\,
            I => \N__29301\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__29310\,
            I => \N__29298\
        );

    \I__5328\ : Span4Mux_h
    port map (
            O => \N__29307\,
            I => \N__29295\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__29304\,
            I => \N__29292\
        );

    \I__5326\ : Span4Mux_h
    port map (
            O => \N__29301\,
            I => \N__29289\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__29298\,
            I => \N__29286\
        );

    \I__5324\ : Span4Mux_v
    port map (
            O => \N__29295\,
            I => \N__29281\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__29292\,
            I => \N__29281\
        );

    \I__5322\ : Sp12to4
    port map (
            O => \N__29289\,
            I => \N__29277\
        );

    \I__5321\ : Span4Mux_v
    port map (
            O => \N__29286\,
            I => \N__29274\
        );

    \I__5320\ : Span4Mux_v
    port map (
            O => \N__29281\,
            I => \N__29271\
        );

    \I__5319\ : CEMux
    port map (
            O => \N__29280\,
            I => \N__29268\
        );

    \I__5318\ : Odrv12
    port map (
            O => \N__29277\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__5317\ : Odrv4
    port map (
            O => \N__29274\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__29271\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__29268\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__5314\ : InMux
    port map (
            O => \N__29259\,
            I => \N__29256\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__29256\,
            I => \N__29253\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__29253\,
            I => \N__29248\
        );

    \I__5311\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29245\
        );

    \I__5310\ : InMux
    port map (
            O => \N__29251\,
            I => \N__29242\
        );

    \I__5309\ : Odrv4
    port map (
            O => \N__29248\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__29245\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__29242\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__5306\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29232\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__29232\,
            I => \N__29229\
        );

    \I__5304\ : Span4Mux_v
    port map (
            O => \N__29229\,
            I => \N__29226\
        );

    \I__5303\ : Span4Mux_h
    port map (
            O => \N__29226\,
            I => \N__29223\
        );

    \I__5302\ : Odrv4
    port map (
            O => \N__29223\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__5301\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29217\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__29217\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__5299\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29208\
        );

    \I__5298\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29205\
        );

    \I__5297\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29200\
        );

    \I__5296\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29200\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__29208\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__29205\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__29200\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__5292\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29190\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__29190\,
            I => \N__29186\
        );

    \I__5290\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29183\
        );

    \I__5289\ : Span4Mux_h
    port map (
            O => \N__29186\,
            I => \N__29176\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__29183\,
            I => \N__29176\
        );

    \I__5287\ : InMux
    port map (
            O => \N__29182\,
            I => \N__29171\
        );

    \I__5286\ : InMux
    port map (
            O => \N__29181\,
            I => \N__29171\
        );

    \I__5285\ : Span4Mux_h
    port map (
            O => \N__29176\,
            I => \N__29168\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__29171\,
            I => \N__29165\
        );

    \I__5283\ : Odrv4
    port map (
            O => \N__29168\,
            I => \phase_controller_inst2.stoper_tr.time_passed11\
        );

    \I__5282\ : Odrv12
    port map (
            O => \N__29165\,
            I => \phase_controller_inst2.stoper_tr.time_passed11\
        );

    \I__5281\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29153\
        );

    \I__5280\ : InMux
    port map (
            O => \N__29159\,
            I => \N__29153\
        );

    \I__5279\ : InMux
    port map (
            O => \N__29158\,
            I => \N__29149\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__29153\,
            I => \N__29144\
        );

    \I__5277\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29141\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__29149\,
            I => \N__29138\
        );

    \I__5275\ : InMux
    port map (
            O => \N__29148\,
            I => \N__29133\
        );

    \I__5274\ : InMux
    port map (
            O => \N__29147\,
            I => \N__29133\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__29144\,
            I => \N__29130\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N__29127\
        );

    \I__5271\ : Span4Mux_v
    port map (
            O => \N__29138\,
            I => \N__29122\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__29133\,
            I => \N__29122\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__29130\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__29127\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5267\ : Odrv4
    port map (
            O => \N__29122\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__5266\ : CascadeMux
    port map (
            O => \N__29115\,
            I => \N__29112\
        );

    \I__5265\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29105\
        );

    \I__5264\ : InMux
    port map (
            O => \N__29111\,
            I => \N__29105\
        );

    \I__5263\ : CascadeMux
    port map (
            O => \N__29110\,
            I => \N__29095\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__29105\,
            I => \N__29091\
        );

    \I__5261\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29088\
        );

    \I__5260\ : InMux
    port map (
            O => \N__29103\,
            I => \N__29068\
        );

    \I__5259\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29068\
        );

    \I__5258\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29068\
        );

    \I__5257\ : InMux
    port map (
            O => \N__29100\,
            I => \N__29068\
        );

    \I__5256\ : InMux
    port map (
            O => \N__29099\,
            I => \N__29068\
        );

    \I__5255\ : InMux
    port map (
            O => \N__29098\,
            I => \N__29068\
        );

    \I__5254\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29068\
        );

    \I__5253\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29065\
        );

    \I__5252\ : Span4Mux_v
    port map (
            O => \N__29091\,
            I => \N__29060\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__29088\,
            I => \N__29060\
        );

    \I__5250\ : CascadeMux
    port map (
            O => \N__29087\,
            I => \N__29055\
        );

    \I__5249\ : CascadeMux
    port map (
            O => \N__29086\,
            I => \N__29052\
        );

    \I__5248\ : CascadeMux
    port map (
            O => \N__29085\,
            I => \N__29049\
        );

    \I__5247\ : CascadeMux
    port map (
            O => \N__29084\,
            I => \N__29043\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__29083\,
            I => \N__29040\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29034\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__29065\,
            I => \N__29029\
        );

    \I__5243\ : Span4Mux_h
    port map (
            O => \N__29060\,
            I => \N__29029\
        );

    \I__5242\ : InMux
    port map (
            O => \N__29059\,
            I => \N__29026\
        );

    \I__5241\ : InMux
    port map (
            O => \N__29058\,
            I => \N__29023\
        );

    \I__5240\ : InMux
    port map (
            O => \N__29055\,
            I => \N__29010\
        );

    \I__5239\ : InMux
    port map (
            O => \N__29052\,
            I => \N__29010\
        );

    \I__5238\ : InMux
    port map (
            O => \N__29049\,
            I => \N__29010\
        );

    \I__5237\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29010\
        );

    \I__5236\ : InMux
    port map (
            O => \N__29047\,
            I => \N__29010\
        );

    \I__5235\ : InMux
    port map (
            O => \N__29046\,
            I => \N__29010\
        );

    \I__5234\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29003\
        );

    \I__5233\ : InMux
    port map (
            O => \N__29040\,
            I => \N__29003\
        );

    \I__5232\ : InMux
    port map (
            O => \N__29039\,
            I => \N__29003\
        );

    \I__5231\ : InMux
    port map (
            O => \N__29038\,
            I => \N__28998\
        );

    \I__5230\ : InMux
    port map (
            O => \N__29037\,
            I => \N__28998\
        );

    \I__5229\ : Span4Mux_h
    port map (
            O => \N__29034\,
            I => \N__28993\
        );

    \I__5228\ : Span4Mux_h
    port map (
            O => \N__29029\,
            I => \N__28993\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__29026\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__29023\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__29010\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__29003\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__28998\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5222\ : Odrv4
    port map (
            O => \N__28993\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__5221\ : CascadeMux
    port map (
            O => \N__28980\,
            I => \N__28975\
        );

    \I__5220\ : CascadeMux
    port map (
            O => \N__28979\,
            I => \N__28972\
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__28978\,
            I => \N__28969\
        );

    \I__5218\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28956\
        );

    \I__5217\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28956\
        );

    \I__5216\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28956\
        );

    \I__5215\ : CascadeMux
    port map (
            O => \N__28968\,
            I => \N__28953\
        );

    \I__5214\ : CascadeMux
    port map (
            O => \N__28967\,
            I => \N__28950\
        );

    \I__5213\ : CascadeMux
    port map (
            O => \N__28966\,
            I => \N__28947\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__28965\,
            I => \N__28938\
        );

    \I__5211\ : InMux
    port map (
            O => \N__28964\,
            I => \N__28928\
        );

    \I__5210\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28928\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__28956\,
            I => \N__28924\
        );

    \I__5208\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28913\
        );

    \I__5207\ : InMux
    port map (
            O => \N__28950\,
            I => \N__28913\
        );

    \I__5206\ : InMux
    port map (
            O => \N__28947\,
            I => \N__28913\
        );

    \I__5205\ : InMux
    port map (
            O => \N__28946\,
            I => \N__28913\
        );

    \I__5204\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28913\
        );

    \I__5203\ : InMux
    port map (
            O => \N__28944\,
            I => \N__28906\
        );

    \I__5202\ : InMux
    port map (
            O => \N__28943\,
            I => \N__28906\
        );

    \I__5201\ : InMux
    port map (
            O => \N__28942\,
            I => \N__28906\
        );

    \I__5200\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28891\
        );

    \I__5199\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28891\
        );

    \I__5198\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28891\
        );

    \I__5197\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28891\
        );

    \I__5196\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28891\
        );

    \I__5195\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28891\
        );

    \I__5194\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28891\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__28928\,
            I => \N__28888\
        );

    \I__5192\ : CascadeMux
    port map (
            O => \N__28927\,
            I => \N__28884\
        );

    \I__5191\ : Span4Mux_v
    port map (
            O => \N__28924\,
            I => \N__28878\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__28913\,
            I => \N__28878\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__28906\,
            I => \N__28875\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__28891\,
            I => \N__28870\
        );

    \I__5187\ : Span4Mux_h
    port map (
            O => \N__28888\,
            I => \N__28870\
        );

    \I__5186\ : InMux
    port map (
            O => \N__28887\,
            I => \N__28867\
        );

    \I__5185\ : InMux
    port map (
            O => \N__28884\,
            I => \N__28861\
        );

    \I__5184\ : InMux
    port map (
            O => \N__28883\,
            I => \N__28861\
        );

    \I__5183\ : Span4Mux_h
    port map (
            O => \N__28878\,
            I => \N__28858\
        );

    \I__5182\ : Span4Mux_h
    port map (
            O => \N__28875\,
            I => \N__28855\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__28870\,
            I => \N__28850\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__28867\,
            I => \N__28850\
        );

    \I__5179\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28847\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__28861\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__28858\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__28855\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__5175\ : Odrv4
    port map (
            O => \N__28850\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__28847\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__28836\,
            I => \N__28833\
        );

    \I__5172\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28797\
        );

    \I__5171\ : InMux
    port map (
            O => \N__28832\,
            I => \N__28797\
        );

    \I__5170\ : InMux
    port map (
            O => \N__28831\,
            I => \N__28797\
        );

    \I__5169\ : InMux
    port map (
            O => \N__28830\,
            I => \N__28797\
        );

    \I__5168\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28797\
        );

    \I__5167\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28797\
        );

    \I__5166\ : InMux
    port map (
            O => \N__28827\,
            I => \N__28797\
        );

    \I__5165\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28797\
        );

    \I__5164\ : InMux
    port map (
            O => \N__28825\,
            I => \N__28790\
        );

    \I__5163\ : InMux
    port map (
            O => \N__28824\,
            I => \N__28790\
        );

    \I__5162\ : InMux
    port map (
            O => \N__28823\,
            I => \N__28790\
        );

    \I__5161\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28785\
        );

    \I__5160\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28785\
        );

    \I__5159\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28770\
        );

    \I__5158\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28770\
        );

    \I__5157\ : InMux
    port map (
            O => \N__28818\,
            I => \N__28770\
        );

    \I__5156\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28770\
        );

    \I__5155\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28770\
        );

    \I__5154\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28770\
        );

    \I__5153\ : InMux
    port map (
            O => \N__28814\,
            I => \N__28770\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__28797\,
            I => \N__28764\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__28790\,
            I => \N__28761\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__28785\,
            I => \N__28758\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__28770\,
            I => \N__28755\
        );

    \I__5148\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28752\
        );

    \I__5147\ : InMux
    port map (
            O => \N__28768\,
            I => \N__28746\
        );

    \I__5146\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28746\
        );

    \I__5145\ : Span4Mux_h
    port map (
            O => \N__28764\,
            I => \N__28743\
        );

    \I__5144\ : Span4Mux_h
    port map (
            O => \N__28761\,
            I => \N__28740\
        );

    \I__5143\ : Span12Mux_v
    port map (
            O => \N__28758\,
            I => \N__28737\
        );

    \I__5142\ : Span4Mux_h
    port map (
            O => \N__28755\,
            I => \N__28732\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__28752\,
            I => \N__28732\
        );

    \I__5140\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28729\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__28746\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__28743\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__28740\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__5136\ : Odrv12
    port map (
            O => \N__28737\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__28732\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__28729\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__5133\ : InMux
    port map (
            O => \N__28716\,
            I => \N__28713\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__28713\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__5131\ : InMux
    port map (
            O => \N__28710\,
            I => \N__28707\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__28707\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__5129\ : InMux
    port map (
            O => \N__28704\,
            I => \N__28700\
        );

    \I__5128\ : CascadeMux
    port map (
            O => \N__28703\,
            I => \N__28695\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__28700\,
            I => \N__28688\
        );

    \I__5126\ : InMux
    port map (
            O => \N__28699\,
            I => \N__28677\
        );

    \I__5125\ : InMux
    port map (
            O => \N__28698\,
            I => \N__28677\
        );

    \I__5124\ : InMux
    port map (
            O => \N__28695\,
            I => \N__28677\
        );

    \I__5123\ : InMux
    port map (
            O => \N__28694\,
            I => \N__28677\
        );

    \I__5122\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28672\
        );

    \I__5121\ : InMux
    port map (
            O => \N__28692\,
            I => \N__28672\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__28691\,
            I => \N__28668\
        );

    \I__5119\ : Span4Mux_h
    port map (
            O => \N__28688\,
            I => \N__28664\
        );

    \I__5118\ : InMux
    port map (
            O => \N__28687\,
            I => \N__28659\
        );

    \I__5117\ : InMux
    port map (
            O => \N__28686\,
            I => \N__28659\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__28677\,
            I => \N__28654\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__28672\,
            I => \N__28654\
        );

    \I__5114\ : InMux
    port map (
            O => \N__28671\,
            I => \N__28647\
        );

    \I__5113\ : InMux
    port map (
            O => \N__28668\,
            I => \N__28647\
        );

    \I__5112\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28647\
        );

    \I__5111\ : Odrv4
    port map (
            O => \N__28664\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__28659\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__5109\ : Odrv4
    port map (
            O => \N__28654\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__28647\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__5107\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28635\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__28635\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\
        );

    \I__5105\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28629\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__28629\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__28626\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\
        );

    \I__5102\ : InMux
    port map (
            O => \N__28623\,
            I => \N__28620\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__28620\,
            I => \N__28616\
        );

    \I__5100\ : InMux
    port map (
            O => \N__28619\,
            I => \N__28613\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__28616\,
            I => \phase_controller_inst1.stoper_tr.N_257\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__28613\,
            I => \phase_controller_inst1.stoper_tr.N_257\
        );

    \I__5097\ : CascadeMux
    port map (
            O => \N__28608\,
            I => \phase_controller_inst1.stoper_tr.N_257_cascade_\
        );

    \I__5096\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28599\
        );

    \I__5095\ : InMux
    port map (
            O => \N__28604\,
            I => \N__28599\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28594\
        );

    \I__5093\ : InMux
    port map (
            O => \N__28598\,
            I => \N__28589\
        );

    \I__5092\ : InMux
    port map (
            O => \N__28597\,
            I => \N__28589\
        );

    \I__5091\ : Odrv4
    port map (
            O => \N__28594\,
            I => \phase_controller_inst1.stoper_tr.N_240\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__28589\,
            I => \phase_controller_inst1.stoper_tr.N_240\
        );

    \I__5089\ : InMux
    port map (
            O => \N__28584\,
            I => \N__28578\
        );

    \I__5088\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28578\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__28578\,
            I => \N__28574\
        );

    \I__5086\ : InMux
    port map (
            O => \N__28577\,
            I => \N__28571\
        );

    \I__5085\ : Odrv12
    port map (
            O => \N__28574\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__28571\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__5083\ : InMux
    port map (
            O => \N__28566\,
            I => \N__28563\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__28563\,
            I => \N__28560\
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__28560\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\
        );

    \I__5080\ : InMux
    port map (
            O => \N__28557\,
            I => \N__28554\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__28554\,
            I => \N__28551\
        );

    \I__5078\ : Span4Mux_v
    port map (
            O => \N__28551\,
            I => \N__28548\
        );

    \I__5077\ : Odrv4
    port map (
            O => \N__28548\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__5076\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28541\
        );

    \I__5075\ : InMux
    port map (
            O => \N__28544\,
            I => \N__28538\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__28541\,
            I => \N__28535\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__28538\,
            I => \N__28532\
        );

    \I__5072\ : Odrv4
    port map (
            O => \N__28535\,
            I => \current_shift_inst.un4_control_input_0_31\
        );

    \I__5071\ : Odrv12
    port map (
            O => \N__28532\,
            I => \current_shift_inst.un4_control_input_0_31\
        );

    \I__5070\ : IoInMux
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28521\
        );

    \I__5068\ : Odrv12
    port map (
            O => \N__28521\,
            I => \delay_measurement_inst.delay_tr_timer.N_463_i\
        );

    \I__5067\ : InMux
    port map (
            O => \N__28518\,
            I => \N__28514\
        );

    \I__5066\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28511\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__28514\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__28511\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__5063\ : InMux
    port map (
            O => \N__28506\,
            I => \N__28502\
        );

    \I__5062\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28498\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__28502\,
            I => \N__28495\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28501\,
            I => \N__28492\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__28498\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__5058\ : Odrv4
    port map (
            O => \N__28495\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__28492\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__5056\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28482\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__28482\,
            I => \N__28478\
        );

    \I__5054\ : InMux
    port map (
            O => \N__28481\,
            I => \N__28475\
        );

    \I__5053\ : Sp12to4
    port map (
            O => \N__28478\,
            I => \N__28469\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__28475\,
            I => \N__28469\
        );

    \I__5051\ : InMux
    port map (
            O => \N__28474\,
            I => \N__28466\
        );

    \I__5050\ : Odrv12
    port map (
            O => \N__28469\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__28466\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__5048\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28458\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__28458\,
            I => \N__28455\
        );

    \I__5046\ : Span4Mux_h
    port map (
            O => \N__28455\,
            I => \N__28452\
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__28452\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\
        );

    \I__5044\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28446\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__28446\,
            I => \N__28443\
        );

    \I__5042\ : Span4Mux_v
    port map (
            O => \N__28443\,
            I => \N__28440\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__28440\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__5040\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__28434\,
            I => \N__28430\
        );

    \I__5038\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28427\
        );

    \I__5037\ : Sp12to4
    port map (
            O => \N__28430\,
            I => \N__28421\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__28427\,
            I => \N__28421\
        );

    \I__5035\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28418\
        );

    \I__5034\ : Odrv12
    port map (
            O => \N__28421\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__28418\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__5032\ : InMux
    port map (
            O => \N__28413\,
            I => \N__28410\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__28410\,
            I => \N__28407\
        );

    \I__5030\ : Odrv4
    port map (
            O => \N__28407\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__5029\ : InMux
    port map (
            O => \N__28404\,
            I => \N__28401\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__28401\,
            I => \N__28396\
        );

    \I__5027\ : InMux
    port map (
            O => \N__28400\,
            I => \N__28391\
        );

    \I__5026\ : InMux
    port map (
            O => \N__28399\,
            I => \N__28391\
        );

    \I__5025\ : Odrv4
    port map (
            O => \N__28396\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__28391\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__5023\ : InMux
    port map (
            O => \N__28386\,
            I => \N__28383\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__28383\,
            I => \N__28380\
        );

    \I__5021\ : Span4Mux_h
    port map (
            O => \N__28380\,
            I => \N__28377\
        );

    \I__5020\ : Odrv4
    port map (
            O => \N__28377\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__5019\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28371\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__28371\,
            I => \N__28367\
        );

    \I__5017\ : InMux
    port map (
            O => \N__28370\,
            I => \N__28364\
        );

    \I__5016\ : Sp12to4
    port map (
            O => \N__28367\,
            I => \N__28358\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__28364\,
            I => \N__28358\
        );

    \I__5014\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28355\
        );

    \I__5013\ : Odrv12
    port map (
            O => \N__28358\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__28355\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5011\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28347\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__28347\,
            I => \N__28344\
        );

    \I__5009\ : Odrv12
    port map (
            O => \N__28344\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\
        );

    \I__5008\ : InMux
    port map (
            O => \N__28341\,
            I => \N__28338\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__28338\,
            I => \N__28334\
        );

    \I__5006\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28331\
        );

    \I__5005\ : Sp12to4
    port map (
            O => \N__28334\,
            I => \N__28325\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__28331\,
            I => \N__28325\
        );

    \I__5003\ : InMux
    port map (
            O => \N__28330\,
            I => \N__28322\
        );

    \I__5002\ : Odrv12
    port map (
            O => \N__28325\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__28322\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__5000\ : InMux
    port map (
            O => \N__28317\,
            I => \N__28314\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__28314\,
            I => \N__28311\
        );

    \I__4998\ : Odrv4
    port map (
            O => \N__28311\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\
        );

    \I__4997\ : InMux
    port map (
            O => \N__28308\,
            I => \N__28305\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__28305\,
            I => \N__28301\
        );

    \I__4995\ : InMux
    port map (
            O => \N__28304\,
            I => \N__28298\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__28301\,
            I => \N__28294\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__28298\,
            I => \N__28291\
        );

    \I__4992\ : InMux
    port map (
            O => \N__28297\,
            I => \N__28288\
        );

    \I__4991\ : Odrv4
    port map (
            O => \N__28294\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__4990\ : Odrv12
    port map (
            O => \N__28291\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__28288\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__4988\ : InMux
    port map (
            O => \N__28281\,
            I => \N__28278\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__28278\,
            I => \N__28275\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__28275\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\
        );

    \I__4985\ : InMux
    port map (
            O => \N__28272\,
            I => \N__28269\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__28269\,
            I => \N__28265\
        );

    \I__4983\ : InMux
    port map (
            O => \N__28268\,
            I => \N__28262\
        );

    \I__4982\ : Span4Mux_v
    port map (
            O => \N__28265\,
            I => \N__28258\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__28262\,
            I => \N__28255\
        );

    \I__4980\ : InMux
    port map (
            O => \N__28261\,
            I => \N__28252\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__28258\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__4978\ : Odrv12
    port map (
            O => \N__28255\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__28252\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__4976\ : InMux
    port map (
            O => \N__28245\,
            I => \N__28242\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__28242\,
            I => \N__28239\
        );

    \I__4974\ : Odrv4
    port map (
            O => \N__28239\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\
        );

    \I__4973\ : InMux
    port map (
            O => \N__28236\,
            I => \N__28233\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__28233\,
            I => \N__28230\
        );

    \I__4971\ : Odrv4
    port map (
            O => \N__28230\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\
        );

    \I__4970\ : CascadeMux
    port map (
            O => \N__28227\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\
        );

    \I__4969\ : InMux
    port map (
            O => \N__28224\,
            I => \N__28221\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__28221\,
            I => \N__28218\
        );

    \I__4967\ : Span4Mux_h
    port map (
            O => \N__28218\,
            I => \N__28215\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__28215\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__4965\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28209\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__28209\,
            I => \N__28206\
        );

    \I__4963\ : Span4Mux_v
    port map (
            O => \N__28206\,
            I => \N__28201\
        );

    \I__4962\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28198\
        );

    \I__4961\ : InMux
    port map (
            O => \N__28204\,
            I => \N__28195\
        );

    \I__4960\ : Odrv4
    port map (
            O => \N__28201\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__28198\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__28195\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__4957\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28185\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__28185\,
            I => \N__28182\
        );

    \I__4955\ : Span12Mux_v
    port map (
            O => \N__28182\,
            I => \N__28179\
        );

    \I__4954\ : Odrv12
    port map (
            O => \N__28179\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__4953\ : InMux
    port map (
            O => \N__28176\,
            I => \N__28173\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__4951\ : Span4Mux_v
    port map (
            O => \N__28170\,
            I => \N__28167\
        );

    \I__4950\ : Odrv4
    port map (
            O => \N__28167\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__4949\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28161\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__28161\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__4947\ : InMux
    port map (
            O => \N__28158\,
            I => \N__28155\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__28155\,
            I => \N__28152\
        );

    \I__4945\ : Span4Mux_h
    port map (
            O => \N__28152\,
            I => \N__28149\
        );

    \I__4944\ : Span4Mux_v
    port map (
            O => \N__28149\,
            I => \N__28146\
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__28146\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__4942\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28134\
        );

    \I__4941\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28134\
        );

    \I__4940\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28134\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__28134\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__4938\ : InMux
    port map (
            O => \N__28131\,
            I => \N__28128\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__28128\,
            I => \N__28125\
        );

    \I__4936\ : Odrv4
    port map (
            O => \N__28125\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__4935\ : InMux
    port map (
            O => \N__28122\,
            I => \N__28119\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28115\
        );

    \I__4933\ : InMux
    port map (
            O => \N__28118\,
            I => \N__28112\
        );

    \I__4932\ : Span4Mux_v
    port map (
            O => \N__28115\,
            I => \N__28106\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__28112\,
            I => \N__28106\
        );

    \I__4930\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28103\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__28106\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__28103\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__4927\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28095\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__28095\,
            I => \N__28092\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__28092\,
            I => \N__28089\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__28089\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__4923\ : InMux
    port map (
            O => \N__28086\,
            I => \N__28083\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__28083\,
            I => \N__28079\
        );

    \I__4921\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28076\
        );

    \I__4920\ : Span4Mux_v
    port map (
            O => \N__28079\,
            I => \N__28070\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__28076\,
            I => \N__28070\
        );

    \I__4918\ : InMux
    port map (
            O => \N__28075\,
            I => \N__28067\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__28070\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__28067\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__4915\ : InMux
    port map (
            O => \N__28062\,
            I => \N__28059\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__28059\,
            I => \N__28056\
        );

    \I__4913\ : Span4Mux_h
    port map (
            O => \N__28056\,
            I => \N__28053\
        );

    \I__4912\ : Odrv4
    port map (
            O => \N__28053\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\
        );

    \I__4911\ : InMux
    port map (
            O => \N__28050\,
            I => \N__28047\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__28047\,
            I => \N__28043\
        );

    \I__4909\ : InMux
    port map (
            O => \N__28046\,
            I => \N__28040\
        );

    \I__4908\ : Span4Mux_v
    port map (
            O => \N__28043\,
            I => \N__28034\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__28040\,
            I => \N__28034\
        );

    \I__4906\ : InMux
    port map (
            O => \N__28039\,
            I => \N__28031\
        );

    \I__4905\ : Odrv4
    port map (
            O => \N__28034\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__28031\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__4903\ : InMux
    port map (
            O => \N__28026\,
            I => \N__28023\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__28023\,
            I => \N__28020\
        );

    \I__4901\ : Span4Mux_h
    port map (
            O => \N__28020\,
            I => \N__28017\
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__28017\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__4899\ : InMux
    port map (
            O => \N__28014\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__4898\ : InMux
    port map (
            O => \N__28011\,
            I => \N__28008\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__28008\,
            I => \N__28005\
        );

    \I__4896\ : Odrv12
    port map (
            O => \N__28005\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__4895\ : InMux
    port map (
            O => \N__28002\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__4894\ : InMux
    port map (
            O => \N__27999\,
            I => \N__27992\
        );

    \I__4893\ : InMux
    port map (
            O => \N__27998\,
            I => \N__27992\
        );

    \I__4892\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27989\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__27992\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__27989\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__4889\ : InMux
    port map (
            O => \N__27984\,
            I => \bfn_11_17_0_\
        );

    \I__4888\ : InMux
    port map (
            O => \N__27981\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__4887\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27975\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__27975\,
            I => \N__27970\
        );

    \I__4885\ : InMux
    port map (
            O => \N__27974\,
            I => \N__27965\
        );

    \I__4884\ : InMux
    port map (
            O => \N__27973\,
            I => \N__27965\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__27970\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__27965\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__4881\ : InMux
    port map (
            O => \N__27960\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__4880\ : InMux
    port map (
            O => \N__27957\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__4879\ : InMux
    port map (
            O => \N__27954\,
            I => \N__27951\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__27951\,
            I => \N__27947\
        );

    \I__4877\ : InMux
    port map (
            O => \N__27950\,
            I => \N__27944\
        );

    \I__4876\ : Span4Mux_v
    port map (
            O => \N__27947\,
            I => \N__27938\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__27944\,
            I => \N__27938\
        );

    \I__4874\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27935\
        );

    \I__4873\ : Odrv4
    port map (
            O => \N__27938\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__27935\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__4871\ : InMux
    port map (
            O => \N__27930\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__4870\ : InMux
    port map (
            O => \N__27927\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__4869\ : InMux
    port map (
            O => \N__27924\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__4868\ : InMux
    port map (
            O => \N__27921\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__4867\ : InMux
    port map (
            O => \N__27918\,
            I => \N__27915\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__27915\,
            I => \N__27912\
        );

    \I__4865\ : Odrv4
    port map (
            O => \N__27912\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__4864\ : InMux
    port map (
            O => \N__27909\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__4863\ : InMux
    port map (
            O => \N__27906\,
            I => \N__27903\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__27903\,
            I => \N__27900\
        );

    \I__4861\ : Odrv4
    port map (
            O => \N__27900\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__4860\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27894\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__27894\,
            I => \N__27890\
        );

    \I__4858\ : InMux
    port map (
            O => \N__27893\,
            I => \N__27887\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__27890\,
            I => \N__27882\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__27887\,
            I => \N__27882\
        );

    \I__4855\ : Span4Mux_v
    port map (
            O => \N__27882\,
            I => \N__27878\
        );

    \I__4854\ : InMux
    port map (
            O => \N__27881\,
            I => \N__27875\
        );

    \I__4853\ : Odrv4
    port map (
            O => \N__27878\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__27875\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__4851\ : InMux
    port map (
            O => \N__27870\,
            I => \bfn_11_16_0_\
        );

    \I__4850\ : InMux
    port map (
            O => \N__27867\,
            I => \N__27864\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__27864\,
            I => \N__27859\
        );

    \I__4848\ : InMux
    port map (
            O => \N__27863\,
            I => \N__27854\
        );

    \I__4847\ : InMux
    port map (
            O => \N__27862\,
            I => \N__27854\
        );

    \I__4846\ : Odrv12
    port map (
            O => \N__27859\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__27854\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__4844\ : InMux
    port map (
            O => \N__27849\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__4843\ : InMux
    port map (
            O => \N__27846\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__4842\ : InMux
    port map (
            O => \N__27843\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__4841\ : InMux
    port map (
            O => \N__27840\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__4840\ : InMux
    port map (
            O => \N__27837\,
            I => \N__27831\
        );

    \I__4839\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27831\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__27831\,
            I => \N__27828\
        );

    \I__4837\ : Span4Mux_v
    port map (
            O => \N__27828\,
            I => \N__27824\
        );

    \I__4836\ : InMux
    port map (
            O => \N__27827\,
            I => \N__27821\
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__27824\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__27821\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__4833\ : InMux
    port map (
            O => \N__27816\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__4832\ : InMux
    port map (
            O => \N__27813\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__4831\ : InMux
    port map (
            O => \N__27810\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__4830\ : InMux
    port map (
            O => \N__27807\,
            I => \N__27803\
        );

    \I__4829\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27800\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__27803\,
            I => \N__27797\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__27800\,
            I => \N__27794\
        );

    \I__4826\ : Span4Mux_v
    port map (
            O => \N__27797\,
            I => \N__27790\
        );

    \I__4825\ : Span4Mux_v
    port map (
            O => \N__27794\,
            I => \N__27787\
        );

    \I__4824\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27784\
        );

    \I__4823\ : Odrv4
    port map (
            O => \N__27790\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__4822\ : Odrv4
    port map (
            O => \N__27787\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__27784\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__4820\ : InMux
    port map (
            O => \N__27777\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__4819\ : InMux
    port map (
            O => \N__27774\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__4818\ : InMux
    port map (
            O => \N__27771\,
            I => \N__27768\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__27768\,
            I => \N__27765\
        );

    \I__4816\ : Span4Mux_h
    port map (
            O => \N__27765\,
            I => \N__27760\
        );

    \I__4815\ : InMux
    port map (
            O => \N__27764\,
            I => \N__27757\
        );

    \I__4814\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27754\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__27760\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__27757\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__27754\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__4810\ : InMux
    port map (
            O => \N__27747\,
            I => \bfn_11_15_0_\
        );

    \I__4809\ : InMux
    port map (
            O => \N__27744\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__4808\ : InMux
    port map (
            O => \N__27741\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__4807\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27735\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27732\
        );

    \I__4805\ : Span4Mux_v
    port map (
            O => \N__27732\,
            I => \N__27727\
        );

    \I__4804\ : InMux
    port map (
            O => \N__27731\,
            I => \N__27724\
        );

    \I__4803\ : InMux
    port map (
            O => \N__27730\,
            I => \N__27721\
        );

    \I__4802\ : Odrv4
    port map (
            O => \N__27727\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__27724\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__27721\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__4799\ : InMux
    port map (
            O => \N__27714\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__4798\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27708\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__27708\,
            I => \N__27704\
        );

    \I__4796\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27701\
        );

    \I__4795\ : Span4Mux_v
    port map (
            O => \N__27704\,
            I => \N__27696\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__27701\,
            I => \N__27696\
        );

    \I__4793\ : Span4Mux_v
    port map (
            O => \N__27696\,
            I => \N__27692\
        );

    \I__4792\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27689\
        );

    \I__4791\ : Odrv4
    port map (
            O => \N__27692\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__27689\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__4789\ : InMux
    port map (
            O => \N__27684\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__4788\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27678\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__27678\,
            I => \N__27675\
        );

    \I__4786\ : Span4Mux_v
    port map (
            O => \N__27675\,
            I => \N__27672\
        );

    \I__4785\ : Span4Mux_h
    port map (
            O => \N__27672\,
            I => \N__27669\
        );

    \I__4784\ : Span4Mux_v
    port map (
            O => \N__27669\,
            I => \N__27666\
        );

    \I__4783\ : Odrv4
    port map (
            O => \N__27666\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__27663\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__4781\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27657\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__27657\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__27654\,
            I => \N__27649\
        );

    \I__4778\ : InMux
    port map (
            O => \N__27653\,
            I => \N__27646\
        );

    \I__4777\ : InMux
    port map (
            O => \N__27652\,
            I => \N__27643\
        );

    \I__4776\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27640\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__27646\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__27643\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__27640\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__4772\ : InMux
    port map (
            O => \N__27633\,
            I => \N__27630\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__27630\,
            I => \N__27627\
        );

    \I__4770\ : Span4Mux_v
    port map (
            O => \N__27627\,
            I => \N__27622\
        );

    \I__4769\ : InMux
    port map (
            O => \N__27626\,
            I => \N__27617\
        );

    \I__4768\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27617\
        );

    \I__4767\ : Odrv4
    port map (
            O => \N__27622\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__27617\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__4765\ : InMux
    port map (
            O => \N__27612\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__4764\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27606\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__27606\,
            I => \N__27603\
        );

    \I__4762\ : Span4Mux_v
    port map (
            O => \N__27603\,
            I => \N__27598\
        );

    \I__4761\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27593\
        );

    \I__4760\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27593\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__27598\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__27593\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__4757\ : InMux
    port map (
            O => \N__27588\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__4756\ : InMux
    port map (
            O => \N__27585\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__27582\,
            I => \N__27579\
        );

    \I__4754\ : InMux
    port map (
            O => \N__27579\,
            I => \N__27576\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__27576\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__4752\ : CascadeMux
    port map (
            O => \N__27573\,
            I => \N__27570\
        );

    \I__4751\ : InMux
    port map (
            O => \N__27570\,
            I => \N__27567\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__27567\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__4749\ : CascadeMux
    port map (
            O => \N__27564\,
            I => \N__27561\
        );

    \I__4748\ : InMux
    port map (
            O => \N__27561\,
            I => \N__27558\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__27558\,
            I => \N__27555\
        );

    \I__4746\ : Odrv4
    port map (
            O => \N__27555\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__4745\ : CascadeMux
    port map (
            O => \N__27552\,
            I => \N__27549\
        );

    \I__4744\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27546\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__27546\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__27543\,
            I => \N__27540\
        );

    \I__4741\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27537\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__27537\,
            I => \N__27534\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__27534\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__27531\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__4737\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27525\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__27525\,
            I => \N__27522\
        );

    \I__4735\ : Span4Mux_h
    port map (
            O => \N__27522\,
            I => \N__27519\
        );

    \I__4734\ : Span4Mux_v
    port map (
            O => \N__27519\,
            I => \N__27516\
        );

    \I__4733\ : Odrv4
    port map (
            O => \N__27516\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__27513\,
            I => \N__27510\
        );

    \I__4731\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27507\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__27507\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__4729\ : InMux
    port map (
            O => \N__27504\,
            I => \N__27501\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__27501\,
            I => \N__27498\
        );

    \I__4727\ : Span4Mux_h
    port map (
            O => \N__27498\,
            I => \N__27494\
        );

    \I__4726\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27491\
        );

    \I__4725\ : Odrv4
    port map (
            O => \N__27494\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__27491\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__4723\ : InMux
    port map (
            O => \N__27486\,
            I => \N__27483\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__27483\,
            I => \N__27480\
        );

    \I__4721\ : Span4Mux_h
    port map (
            O => \N__27480\,
            I => \N__27477\
        );

    \I__4720\ : Sp12to4
    port map (
            O => \N__27477\,
            I => \N__27474\
        );

    \I__4719\ : Span12Mux_s10_v
    port map (
            O => \N__27474\,
            I => \N__27469\
        );

    \I__4718\ : CascadeMux
    port map (
            O => \N__27473\,
            I => \N__27466\
        );

    \I__4717\ : CascadeMux
    port map (
            O => \N__27472\,
            I => \N__27463\
        );

    \I__4716\ : Span12Mux_v
    port map (
            O => \N__27469\,
            I => \N__27459\
        );

    \I__4715\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27456\
        );

    \I__4714\ : InMux
    port map (
            O => \N__27463\,
            I => \N__27453\
        );

    \I__4713\ : InMux
    port map (
            O => \N__27462\,
            I => \N__27450\
        );

    \I__4712\ : Odrv12
    port map (
            O => \N__27459\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__27456\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__27453\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__27450\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4708\ : InMux
    port map (
            O => \N__27441\,
            I => \N__27436\
        );

    \I__4707\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27433\
        );

    \I__4706\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27430\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__27436\,
            I => \N__27427\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__27433\,
            I => \N__27424\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__27430\,
            I => \N__27421\
        );

    \I__4702\ : Span4Mux_v
    port map (
            O => \N__27427\,
            I => \N__27418\
        );

    \I__4701\ : Span4Mux_h
    port map (
            O => \N__27424\,
            I => \N__27415\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__27421\,
            I => \il_max_comp2_D2\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__27418\,
            I => \il_max_comp2_D2\
        );

    \I__4698\ : Odrv4
    port map (
            O => \N__27415\,
            I => \il_max_comp2_D2\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__27408\,
            I => \N__27405\
        );

    \I__4696\ : InMux
    port map (
            O => \N__27405\,
            I => \N__27402\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__27402\,
            I => \N__27399\
        );

    \I__4694\ : Span4Mux_h
    port map (
            O => \N__27399\,
            I => \N__27396\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__27396\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__27393\,
            I => \N__27390\
        );

    \I__4691\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27387\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__27387\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__4689\ : CascadeMux
    port map (
            O => \N__27384\,
            I => \N__27381\
        );

    \I__4688\ : InMux
    port map (
            O => \N__27381\,
            I => \N__27378\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__27378\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__4686\ : CascadeMux
    port map (
            O => \N__27375\,
            I => \N__27372\
        );

    \I__4685\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27369\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__27369\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__4683\ : CascadeMux
    port map (
            O => \N__27366\,
            I => \N__27363\
        );

    \I__4682\ : InMux
    port map (
            O => \N__27363\,
            I => \N__27360\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__27360\,
            I => \N__27357\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__27357\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__4679\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27351\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__27351\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\
        );

    \I__4677\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27345\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__27345\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\
        );

    \I__4675\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27339\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__27339\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__4673\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27333\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__27333\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\
        );

    \I__4671\ : InMux
    port map (
            O => \N__27330\,
            I => \N__27327\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__27327\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__4669\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27321\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__27321\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__4667\ : InMux
    port map (
            O => \N__27318\,
            I => \N__27315\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__27315\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\
        );

    \I__4665\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27309\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__27309\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__4663\ : InMux
    port map (
            O => \N__27306\,
            I => \N__27303\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__27303\,
            I => \N__27300\
        );

    \I__4661\ : Odrv4
    port map (
            O => \N__27300\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__4660\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27294\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__27294\,
            I => \N__27291\
        );

    \I__4658\ : Span4Mux_h
    port map (
            O => \N__27291\,
            I => \N__27288\
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__27288\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__4656\ : InMux
    port map (
            O => \N__27285\,
            I => \N__27282\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__27282\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\
        );

    \I__4654\ : InMux
    port map (
            O => \N__27279\,
            I => \N__27276\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__27276\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__4652\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27270\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__27270\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\
        );

    \I__4650\ : InMux
    port map (
            O => \N__27267\,
            I => \N__27264\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__27264\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\
        );

    \I__4648\ : InMux
    port map (
            O => \N__27261\,
            I => \N__27258\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__27258\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__4646\ : InMux
    port map (
            O => \N__27255\,
            I => \N__27252\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__27252\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\
        );

    \I__4644\ : InMux
    port map (
            O => \N__27249\,
            I => \N__27246\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__27246\,
            I => \N__27243\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__27243\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\
        );

    \I__4641\ : InMux
    port map (
            O => \N__27240\,
            I => \N__27237\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__27237\,
            I => \N__27234\
        );

    \I__4639\ : Odrv4
    port map (
            O => \N__27234\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\
        );

    \I__4638\ : InMux
    port map (
            O => \N__27231\,
            I => \N__27228\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__27228\,
            I => \N__27225\
        );

    \I__4636\ : Span4Mux_v
    port map (
            O => \N__27225\,
            I => \N__27222\
        );

    \I__4635\ : Odrv4
    port map (
            O => \N__27222\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__4634\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27216\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__27216\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__4632\ : CascadeMux
    port map (
            O => \N__27213\,
            I => \N__27210\
        );

    \I__4631\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__27207\,
            I => \N__27204\
        );

    \I__4629\ : Span4Mux_v
    port map (
            O => \N__27204\,
            I => \N__27201\
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__27201\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__4627\ : InMux
    port map (
            O => \N__27198\,
            I => \N__27195\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__27195\,
            I => \N__27192\
        );

    \I__4625\ : Span4Mux_v
    port map (
            O => \N__27192\,
            I => \N__27189\
        );

    \I__4624\ : Odrv4
    port map (
            O => \N__27189\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__4623\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__27183\,
            I => \N__27180\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__27180\,
            I => \N__27177\
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__27177\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__4619\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__27171\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__27168\,
            I => \N__27165\
        );

    \I__4616\ : InMux
    port map (
            O => \N__27165\,
            I => \N__27162\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__27162\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__4614\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27156\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__27156\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__4612\ : CascadeMux
    port map (
            O => \N__27153\,
            I => \N__27150\
        );

    \I__4611\ : InMux
    port map (
            O => \N__27150\,
            I => \N__27147\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__27147\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__27144\,
            I => \N__27141\
        );

    \I__4608\ : InMux
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__27138\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__4606\ : InMux
    port map (
            O => \N__27135\,
            I => \N__27132\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__27132\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__4604\ : InMux
    port map (
            O => \N__27129\,
            I => \N__27126\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__27126\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__4602\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27120\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__27120\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__4600\ : InMux
    port map (
            O => \N__27117\,
            I => \N__27114\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__27114\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__4598\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27108\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__27108\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__4596\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27102\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__27102\,
            I => \N__27099\
        );

    \I__4594\ : Span4Mux_v
    port map (
            O => \N__27099\,
            I => \N__27096\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__27096\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\
        );

    \I__4592\ : InMux
    port map (
            O => \N__27093\,
            I => \N__27074\
        );

    \I__4591\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27071\
        );

    \I__4590\ : InMux
    port map (
            O => \N__27091\,
            I => \N__27054\
        );

    \I__4589\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27054\
        );

    \I__4588\ : InMux
    port map (
            O => \N__27089\,
            I => \N__27054\
        );

    \I__4587\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27054\
        );

    \I__4586\ : InMux
    port map (
            O => \N__27087\,
            I => \N__27054\
        );

    \I__4585\ : InMux
    port map (
            O => \N__27086\,
            I => \N__27054\
        );

    \I__4584\ : InMux
    port map (
            O => \N__27085\,
            I => \N__27054\
        );

    \I__4583\ : InMux
    port map (
            O => \N__27084\,
            I => \N__27054\
        );

    \I__4582\ : InMux
    port map (
            O => \N__27083\,
            I => \N__27041\
        );

    \I__4581\ : InMux
    port map (
            O => \N__27082\,
            I => \N__27041\
        );

    \I__4580\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27041\
        );

    \I__4579\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27041\
        );

    \I__4578\ : InMux
    port map (
            O => \N__27079\,
            I => \N__27041\
        );

    \I__4577\ : InMux
    port map (
            O => \N__27078\,
            I => \N__27041\
        );

    \I__4576\ : InMux
    port map (
            O => \N__27077\,
            I => \N__27038\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__27074\,
            I => \N__27033\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__27071\,
            I => \N__27033\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__27054\,
            I => \N__27030\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__27041\,
            I => \N__27027\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__27038\,
            I => \N__27014\
        );

    \I__4570\ : Span4Mux_v
    port map (
            O => \N__27033\,
            I => \N__27011\
        );

    \I__4569\ : Span4Mux_v
    port map (
            O => \N__27030\,
            I => \N__27006\
        );

    \I__4568\ : Span4Mux_v
    port map (
            O => \N__27027\,
            I => \N__27006\
        );

    \I__4567\ : InMux
    port map (
            O => \N__27026\,
            I => \N__26997\
        );

    \I__4566\ : InMux
    port map (
            O => \N__27025\,
            I => \N__26997\
        );

    \I__4565\ : InMux
    port map (
            O => \N__27024\,
            I => \N__26997\
        );

    \I__4564\ : InMux
    port map (
            O => \N__27023\,
            I => \N__26997\
        );

    \I__4563\ : InMux
    port map (
            O => \N__27022\,
            I => \N__26986\
        );

    \I__4562\ : InMux
    port map (
            O => \N__27021\,
            I => \N__26986\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27020\,
            I => \N__26986\
        );

    \I__4560\ : InMux
    port map (
            O => \N__27019\,
            I => \N__26986\
        );

    \I__4559\ : InMux
    port map (
            O => \N__27018\,
            I => \N__26986\
        );

    \I__4558\ : InMux
    port map (
            O => \N__27017\,
            I => \N__26983\
        );

    \I__4557\ : Odrv4
    port map (
            O => \N__27014\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__4556\ : Odrv4
    port map (
            O => \N__27011\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__4555\ : Odrv4
    port map (
            O => \N__27006\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__26997\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__26986\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__26983\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__4551\ : CascadeMux
    port map (
            O => \N__26970\,
            I => \N__26966\
        );

    \I__4550\ : InMux
    port map (
            O => \N__26969\,
            I => \N__26963\
        );

    \I__4549\ : InMux
    port map (
            O => \N__26966\,
            I => \N__26960\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__26963\,
            I => \N__26955\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__26960\,
            I => \N__26955\
        );

    \I__4546\ : Span12Mux_v
    port map (
            O => \N__26955\,
            I => \N__26952\
        );

    \I__4545\ : Odrv12
    port map (
            O => \N__26952\,
            I => \current_shift_inst.N_1819_i\
        );

    \I__4544\ : InMux
    port map (
            O => \N__26949\,
            I => \N__26946\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__26946\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__26943\,
            I => \N__26940\
        );

    \I__4541\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26937\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__26937\,
            I => \N__26934\
        );

    \I__4539\ : Span4Mux_v
    port map (
            O => \N__26934\,
            I => \N__26931\
        );

    \I__4538\ : Odrv4
    port map (
            O => \N__26931\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__4537\ : InMux
    port map (
            O => \N__26928\,
            I => \N__26925\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__26925\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__4535\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26919\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__26919\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__4533\ : InMux
    port map (
            O => \N__26916\,
            I => \N__26913\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__26913\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__4531\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26907\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__26904\,
            I => \N__26901\
        );

    \I__4528\ : Odrv4
    port map (
            O => \N__26901\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\
        );

    \I__4527\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__26895\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__4525\ : InMux
    port map (
            O => \N__26892\,
            I => \N__26889\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__26889\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__4523\ : CascadeMux
    port map (
            O => \N__26886\,
            I => \N__26883\
        );

    \I__4522\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26880\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__26880\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__4520\ : InMux
    port map (
            O => \N__26877\,
            I => \N__26874\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__26874\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__4518\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26868\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__26868\,
            I => \N__26865\
        );

    \I__4516\ : Span12Mux_v
    port map (
            O => \N__26865\,
            I => \N__26862\
        );

    \I__4515\ : Odrv12
    port map (
            O => \N__26862\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\
        );

    \I__4514\ : InMux
    port map (
            O => \N__26859\,
            I => \N__26856\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__26856\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__4512\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26850\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__26850\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__4510\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26844\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__26844\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__4508\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26838\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__26838\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__4506\ : InMux
    port map (
            O => \N__26835\,
            I => \N__26832\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__26832\,
            I => \N__26829\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__26829\,
            I => \N__26826\
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__26826\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\
        );

    \I__4502\ : InMux
    port map (
            O => \N__26823\,
            I => \N__26820\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__26820\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__4500\ : InMux
    port map (
            O => \N__26817\,
            I => \N__26814\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__26814\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__4498\ : InMux
    port map (
            O => \N__26811\,
            I => \N__26808\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__26808\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__4496\ : InMux
    port map (
            O => \N__26805\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__4495\ : CascadeMux
    port map (
            O => \N__26802\,
            I => \N__26799\
        );

    \I__4494\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26796\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__26796\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__26793\,
            I => \N__26790\
        );

    \I__4491\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26787\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__26787\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__26784\,
            I => \N__26781\
        );

    \I__4488\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26778\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__26778\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__4486\ : InMux
    port map (
            O => \N__26775\,
            I => \N__26772\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__26772\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__4484\ : CascadeMux
    port map (
            O => \N__26769\,
            I => \N__26766\
        );

    \I__4483\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26763\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__26763\,
            I => \N__26759\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__26762\,
            I => \N__26756\
        );

    \I__4480\ : Span4Mux_v
    port map (
            O => \N__26759\,
            I => \N__26751\
        );

    \I__4479\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26748\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__26755\,
            I => \N__26745\
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__26754\,
            I => \N__26742\
        );

    \I__4476\ : Span4Mux_v
    port map (
            O => \N__26751\,
            I => \N__26739\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__26748\,
            I => \N__26736\
        );

    \I__4474\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26733\
        );

    \I__4473\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26730\
        );

    \I__4472\ : Odrv4
    port map (
            O => \N__26739\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__4471\ : Odrv4
    port map (
            O => \N__26736\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__26733\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__26730\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__4468\ : InMux
    port map (
            O => \N__26721\,
            I => \N__26718\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__26718\,
            I => \N__26715\
        );

    \I__4466\ : Span4Mux_v
    port map (
            O => \N__26715\,
            I => \N__26712\
        );

    \I__4465\ : Odrv4
    port map (
            O => \N__26712\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__4464\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26706\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__26706\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__4462\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26700\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__26700\,
            I => \N__26697\
        );

    \I__4460\ : Span4Mux_v
    port map (
            O => \N__26697\,
            I => \N__26691\
        );

    \I__4459\ : InMux
    port map (
            O => \N__26696\,
            I => \N__26684\
        );

    \I__4458\ : InMux
    port map (
            O => \N__26695\,
            I => \N__26684\
        );

    \I__4457\ : InMux
    port map (
            O => \N__26694\,
            I => \N__26684\
        );

    \I__4456\ : Odrv4
    port map (
            O => \N__26691\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__26684\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__4454\ : InMux
    port map (
            O => \N__26679\,
            I => \N__26676\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__26676\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__4452\ : InMux
    port map (
            O => \N__26673\,
            I => \N__26670\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__26670\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__26667\,
            I => \N__26664\
        );

    \I__4449\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26661\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__26661\,
            I => \N__26658\
        );

    \I__4447\ : Odrv4
    port map (
            O => \N__26658\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__4446\ : InMux
    port map (
            O => \N__26655\,
            I => \N__26651\
        );

    \I__4445\ : InMux
    port map (
            O => \N__26654\,
            I => \N__26648\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__26651\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__26648\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4442\ : InMux
    port map (
            O => \N__26643\,
            I => \N__26640\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__26640\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__4440\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26633\
        );

    \I__4439\ : InMux
    port map (
            O => \N__26636\,
            I => \N__26630\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__26633\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__26630\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__4436\ : InMux
    port map (
            O => \N__26625\,
            I => \N__26622\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__26622\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__4434\ : InMux
    port map (
            O => \N__26619\,
            I => \N__26615\
        );

    \I__4433\ : InMux
    port map (
            O => \N__26618\,
            I => \N__26612\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__26615\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__26612\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__4430\ : InMux
    port map (
            O => \N__26607\,
            I => \N__26604\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__26604\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__26601\,
            I => \N__26598\
        );

    \I__4427\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26595\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__26595\,
            I => \N__26592\
        );

    \I__4425\ : Odrv12
    port map (
            O => \N__26592\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__4424\ : InMux
    port map (
            O => \N__26589\,
            I => \N__26586\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__26586\,
            I => \N__26582\
        );

    \I__4422\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26579\
        );

    \I__4421\ : Span4Mux_h
    port map (
            O => \N__26582\,
            I => \N__26576\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__26579\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__4419\ : Odrv4
    port map (
            O => \N__26576\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__4418\ : InMux
    port map (
            O => \N__26571\,
            I => \N__26568\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__26568\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\
        );

    \I__4416\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26561\
        );

    \I__4415\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26558\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__26561\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__26558\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__4412\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26550\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__26550\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\
        );

    \I__4410\ : InMux
    port map (
            O => \N__26547\,
            I => \N__26543\
        );

    \I__4409\ : InMux
    port map (
            O => \N__26546\,
            I => \N__26540\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__26543\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__26540\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__4406\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26532\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__26532\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\
        );

    \I__4404\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26525\
        );

    \I__4403\ : InMux
    port map (
            O => \N__26528\,
            I => \N__26522\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__26525\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__26522\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__4400\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26514\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__26514\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\
        );

    \I__4398\ : CascadeMux
    port map (
            O => \N__26511\,
            I => \N__26508\
        );

    \I__4397\ : InMux
    port map (
            O => \N__26508\,
            I => \N__26505\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__26505\,
            I => \N__26502\
        );

    \I__4395\ : Odrv4
    port map (
            O => \N__26502\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__4394\ : CascadeMux
    port map (
            O => \N__26499\,
            I => \N__26496\
        );

    \I__4393\ : InMux
    port map (
            O => \N__26496\,
            I => \N__26492\
        );

    \I__4392\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26489\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__26492\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__26489\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4389\ : InMux
    port map (
            O => \N__26484\,
            I => \N__26481\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__26481\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__4387\ : InMux
    port map (
            O => \N__26478\,
            I => \N__26474\
        );

    \I__4386\ : InMux
    port map (
            O => \N__26477\,
            I => \N__26471\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__26474\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__26471\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4383\ : InMux
    port map (
            O => \N__26466\,
            I => \N__26463\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__26463\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__4381\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26456\
        );

    \I__4380\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26453\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__26456\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__26453\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4377\ : CascadeMux
    port map (
            O => \N__26448\,
            I => \N__26445\
        );

    \I__4376\ : InMux
    port map (
            O => \N__26445\,
            I => \N__26442\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__26442\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__4374\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26436\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__26436\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__4372\ : InMux
    port map (
            O => \N__26433\,
            I => \N__26429\
        );

    \I__4371\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26426\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__26429\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__26426\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__26421\,
            I => \N__26418\
        );

    \I__4367\ : InMux
    port map (
            O => \N__26418\,
            I => \N__26415\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__26415\,
            I => \N__26412\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__26412\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__4364\ : InMux
    port map (
            O => \N__26409\,
            I => \N__26406\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__26406\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__4362\ : InMux
    port map (
            O => \N__26403\,
            I => \N__26399\
        );

    \I__4361\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26396\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__26399\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__26396\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4358\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26388\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__26388\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__4356\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26381\
        );

    \I__4355\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26378\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__26381\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__26378\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4352\ : InMux
    port map (
            O => \N__26373\,
            I => \N__26370\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__26370\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__26367\,
            I => \N__26364\
        );

    \I__4349\ : InMux
    port map (
            O => \N__26364\,
            I => \N__26361\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__26361\,
            I => \N__26358\
        );

    \I__4347\ : Span4Mux_h
    port map (
            O => \N__26358\,
            I => \N__26355\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__26355\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__4345\ : InMux
    port map (
            O => \N__26352\,
            I => \N__26348\
        );

    \I__4344\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26345\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__26348\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__26345\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4341\ : InMux
    port map (
            O => \N__26340\,
            I => \N__26337\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__26337\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__4339\ : InMux
    port map (
            O => \N__26334\,
            I => \N__26330\
        );

    \I__4338\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26327\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__26330\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__26327\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4335\ : InMux
    port map (
            O => \N__26322\,
            I => \N__26319\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__26319\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__26316\,
            I => \N__26312\
        );

    \I__4332\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26308\
        );

    \I__4331\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26305\
        );

    \I__4330\ : InMux
    port map (
            O => \N__26311\,
            I => \N__26302\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__26308\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__26305\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__26302\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4326\ : InMux
    port map (
            O => \N__26295\,
            I => \N__26292\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__26292\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__4324\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26285\
        );

    \I__4323\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26282\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__26285\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__26282\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4320\ : InMux
    port map (
            O => \N__26277\,
            I => \N__26274\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__26274\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__26271\,
            I => \N__26268\
        );

    \I__4317\ : InMux
    port map (
            O => \N__26268\,
            I => \N__26264\
        );

    \I__4316\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26261\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__26264\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__26261\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4313\ : InMux
    port map (
            O => \N__26256\,
            I => \N__26253\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__26253\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__4311\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26246\
        );

    \I__4310\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26243\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__26246\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__26243\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__4307\ : InMux
    port map (
            O => \N__26238\,
            I => \N__26235\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__26235\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__4305\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26229\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__26229\,
            I => \N__26226\
        );

    \I__4303\ : Span4Mux_v
    port map (
            O => \N__26226\,
            I => \N__26223\
        );

    \I__4302\ : Odrv4
    port map (
            O => \N__26223\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__4301\ : InMux
    port map (
            O => \N__26220\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__4300\ : InMux
    port map (
            O => \N__26217\,
            I => \N__26214\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__26214\,
            I => \N__26211\
        );

    \I__4298\ : Sp12to4
    port map (
            O => \N__26211\,
            I => \N__26208\
        );

    \I__4297\ : Odrv12
    port map (
            O => \N__26208\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__4296\ : InMux
    port map (
            O => \N__26205\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__4295\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26199\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__26199\,
            I => \N__26196\
        );

    \I__4293\ : Sp12to4
    port map (
            O => \N__26196\,
            I => \N__26193\
        );

    \I__4292\ : Odrv12
    port map (
            O => \N__26193\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__4291\ : InMux
    port map (
            O => \N__26190\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__4290\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26184\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__26184\,
            I => \N__26181\
        );

    \I__4288\ : Odrv4
    port map (
            O => \N__26181\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__4287\ : InMux
    port map (
            O => \N__26178\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__4286\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26172\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__26172\,
            I => \N__26169\
        );

    \I__4284\ : Span4Mux_v
    port map (
            O => \N__26169\,
            I => \N__26166\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__26166\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__4282\ : InMux
    port map (
            O => \N__26163\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__4281\ : InMux
    port map (
            O => \N__26160\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__26157\,
            I => \N__26154\
        );

    \I__4279\ : InMux
    port map (
            O => \N__26154\,
            I => \N__26151\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__26151\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__4277\ : IoInMux
    port map (
            O => \N__26148\,
            I => \N__26145\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__26145\,
            I => \N__26142\
        );

    \I__4275\ : Odrv12
    port map (
            O => \N__26142\,
            I => s3_phy_c
        );

    \I__4274\ : InMux
    port map (
            O => \N__26139\,
            I => \N__26136\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__26136\,
            I => \N__26133\
        );

    \I__4272\ : Span4Mux_v
    port map (
            O => \N__26133\,
            I => \N__26130\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__26130\,
            I => \current_shift_inst.un38_control_input_0_s1_17\
        );

    \I__4270\ : InMux
    port map (
            O => \N__26127\,
            I => \current_shift_inst.un38_control_input_cry_16_s1\
        );

    \I__4269\ : InMux
    port map (
            O => \N__26124\,
            I => \N__26121\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__26121\,
            I => \N__26118\
        );

    \I__4267\ : Span4Mux_v
    port map (
            O => \N__26118\,
            I => \N__26115\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__26115\,
            I => \current_shift_inst.un38_control_input_0_s1_18\
        );

    \I__4265\ : InMux
    port map (
            O => \N__26112\,
            I => \current_shift_inst.un38_control_input_cry_17_s1\
        );

    \I__4264\ : InMux
    port map (
            O => \N__26109\,
            I => \N__26106\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__26106\,
            I => \N__26103\
        );

    \I__4262\ : Span4Mux_v
    port map (
            O => \N__26103\,
            I => \N__26100\
        );

    \I__4261\ : Span4Mux_h
    port map (
            O => \N__26100\,
            I => \N__26097\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__26097\,
            I => \current_shift_inst.un38_control_input_0_s1_19\
        );

    \I__4259\ : InMux
    port map (
            O => \N__26094\,
            I => \current_shift_inst.un38_control_input_cry_18_s1\
        );

    \I__4258\ : InMux
    port map (
            O => \N__26091\,
            I => \N__26088\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__26088\,
            I => \N__26085\
        );

    \I__4256\ : Span4Mux_v
    port map (
            O => \N__26085\,
            I => \N__26082\
        );

    \I__4255\ : Odrv4
    port map (
            O => \N__26082\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__4254\ : InMux
    port map (
            O => \N__26079\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__4253\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26073\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__26073\,
            I => \N__26070\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__26070\,
            I => \N__26067\
        );

    \I__4250\ : Odrv4
    port map (
            O => \N__26067\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__4249\ : InMux
    port map (
            O => \N__26064\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__4248\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26058\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__26058\,
            I => \N__26055\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__26055\,
            I => \N__26052\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__26052\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__4244\ : InMux
    port map (
            O => \N__26049\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__4243\ : InMux
    port map (
            O => \N__26046\,
            I => \N__26043\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__26043\,
            I => \N__26040\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__26040\,
            I => \N__26037\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__26037\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__4239\ : InMux
    port map (
            O => \N__26034\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__4238\ : InMux
    port map (
            O => \N__26031\,
            I => \N__26028\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__26028\,
            I => \N__26025\
        );

    \I__4236\ : Span4Mux_v
    port map (
            O => \N__26025\,
            I => \N__26022\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__26022\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__4234\ : InMux
    port map (
            O => \N__26019\,
            I => \bfn_9_22_0_\
        );

    \I__4233\ : InMux
    port map (
            O => \N__26016\,
            I => \N__26013\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__26013\,
            I => \N__26010\
        );

    \I__4231\ : Span4Mux_v
    port map (
            O => \N__26010\,
            I => \N__26007\
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__26007\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__4229\ : InMux
    port map (
            O => \N__26004\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__4228\ : InMux
    port map (
            O => \N__26001\,
            I => \N__25998\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__25998\,
            I => \N__25995\
        );

    \I__4226\ : Odrv12
    port map (
            O => \N__25995\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\
        );

    \I__4225\ : InMux
    port map (
            O => \N__25992\,
            I => \N__25989\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__25989\,
            I => \N__25986\
        );

    \I__4223\ : Span4Mux_v
    port map (
            O => \N__25986\,
            I => \N__25983\
        );

    \I__4222\ : Odrv4
    port map (
            O => \N__25983\,
            I => \current_shift_inst.un38_control_input_0_s1_9\
        );

    \I__4221\ : InMux
    port map (
            O => \N__25980\,
            I => \current_shift_inst.un38_control_input_cry_8_s1\
        );

    \I__4220\ : InMux
    port map (
            O => \N__25977\,
            I => \N__25974\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__25974\,
            I => \N__25971\
        );

    \I__4218\ : Odrv4
    port map (
            O => \N__25971\,
            I => \current_shift_inst.un38_control_input_0_s1_10\
        );

    \I__4217\ : InMux
    port map (
            O => \N__25968\,
            I => \current_shift_inst.un38_control_input_cry_9_s1\
        );

    \I__4216\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25962\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__25962\,
            I => \N__25959\
        );

    \I__4214\ : Span4Mux_v
    port map (
            O => \N__25959\,
            I => \N__25956\
        );

    \I__4213\ : Odrv4
    port map (
            O => \N__25956\,
            I => \current_shift_inst.un38_control_input_0_s1_11\
        );

    \I__4212\ : InMux
    port map (
            O => \N__25953\,
            I => \current_shift_inst.un38_control_input_cry_10_s1\
        );

    \I__4211\ : InMux
    port map (
            O => \N__25950\,
            I => \N__25947\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__25947\,
            I => \N__25944\
        );

    \I__4209\ : Span4Mux_v
    port map (
            O => \N__25944\,
            I => \N__25941\
        );

    \I__4208\ : Odrv4
    port map (
            O => \N__25941\,
            I => \current_shift_inst.un38_control_input_0_s1_12\
        );

    \I__4207\ : InMux
    port map (
            O => \N__25938\,
            I => \current_shift_inst.un38_control_input_cry_11_s1\
        );

    \I__4206\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25932\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__25932\,
            I => \N__25929\
        );

    \I__4204\ : Odrv4
    port map (
            O => \N__25929\,
            I => \current_shift_inst.un38_control_input_0_s1_13\
        );

    \I__4203\ : InMux
    port map (
            O => \N__25926\,
            I => \current_shift_inst.un38_control_input_cry_12_s1\
        );

    \I__4202\ : InMux
    port map (
            O => \N__25923\,
            I => \N__25920\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__25920\,
            I => \N__25917\
        );

    \I__4200\ : Span4Mux_h
    port map (
            O => \N__25917\,
            I => \N__25914\
        );

    \I__4199\ : Span4Mux_v
    port map (
            O => \N__25914\,
            I => \N__25911\
        );

    \I__4198\ : Odrv4
    port map (
            O => \N__25911\,
            I => \current_shift_inst.un38_control_input_0_s1_14\
        );

    \I__4197\ : InMux
    port map (
            O => \N__25908\,
            I => \current_shift_inst.un38_control_input_cry_13_s1\
        );

    \I__4196\ : InMux
    port map (
            O => \N__25905\,
            I => \N__25902\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__25902\,
            I => \N__25899\
        );

    \I__4194\ : Span4Mux_h
    port map (
            O => \N__25899\,
            I => \N__25896\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__25896\,
            I => \current_shift_inst.un38_control_input_0_s1_15\
        );

    \I__4192\ : InMux
    port map (
            O => \N__25893\,
            I => \current_shift_inst.un38_control_input_cry_14_s1\
        );

    \I__4191\ : InMux
    port map (
            O => \N__25890\,
            I => \N__25887\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__25887\,
            I => \N__25884\
        );

    \I__4189\ : Span4Mux_v
    port map (
            O => \N__25884\,
            I => \N__25881\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__25881\,
            I => \current_shift_inst.un38_control_input_0_s1_16\
        );

    \I__4187\ : InMux
    port map (
            O => \N__25878\,
            I => \bfn_9_21_0_\
        );

    \I__4186\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25872\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__25872\,
            I => \N__25869\
        );

    \I__4184\ : Span4Mux_h
    port map (
            O => \N__25869\,
            I => \N__25866\
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__25866\,
            I => \current_shift_inst.un38_control_input_0_s1_6\
        );

    \I__4182\ : InMux
    port map (
            O => \N__25863\,
            I => \current_shift_inst.un38_control_input_cry_5_s1\
        );

    \I__4181\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25857\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__25857\,
            I => \current_shift_inst.un38_control_input_0_s1_7\
        );

    \I__4179\ : InMux
    port map (
            O => \N__25854\,
            I => \current_shift_inst.un38_control_input_cry_6_s1\
        );

    \I__4178\ : InMux
    port map (
            O => \N__25851\,
            I => \N__25848\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__25848\,
            I => \N__25845\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__25845\,
            I => \N__25842\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__25842\,
            I => \current_shift_inst.un38_control_input_0_s1_8\
        );

    \I__4174\ : InMux
    port map (
            O => \N__25839\,
            I => \bfn_9_20_0_\
        );

    \I__4173\ : InMux
    port map (
            O => \N__25836\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__4172\ : InMux
    port map (
            O => \N__25833\,
            I => \N__25830\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__25830\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5\
        );

    \I__4170\ : InMux
    port map (
            O => \N__25827\,
            I => \N__25824\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__25824\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__25821\,
            I => \N__25818\
        );

    \I__4167\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25815\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__25815\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13\
        );

    \I__4165\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__25809\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14\
        );

    \I__4163\ : CascadeMux
    port map (
            O => \N__25806\,
            I => \N__25803\
        );

    \I__4162\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25800\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__25800\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15\
        );

    \I__4160\ : InMux
    port map (
            O => \N__25797\,
            I => \N__25794\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__25794\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17\
        );

    \I__4158\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25788\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__25788\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18\
        );

    \I__4156\ : InMux
    port map (
            O => \N__25785\,
            I => \N__25782\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__25782\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19\
        );

    \I__4154\ : InMux
    port map (
            O => \N__25779\,
            I => \N__25776\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__25776\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2\
        );

    \I__4152\ : InMux
    port map (
            O => \N__25773\,
            I => \N__25770\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__25770\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3\
        );

    \I__4150\ : InMux
    port map (
            O => \N__25767\,
            I => \N__25764\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__25764\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9\
        );

    \I__4148\ : InMux
    port map (
            O => \N__25761\,
            I => \N__25758\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__25758\,
            I => \N__25755\
        );

    \I__4146\ : Span4Mux_h
    port map (
            O => \N__25755\,
            I => \N__25752\
        );

    \I__4145\ : Odrv4
    port map (
            O => \N__25752\,
            I => \il_max_comp2_D1\
        );

    \I__4144\ : InMux
    port map (
            O => \N__25749\,
            I => \N__25746\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__25746\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7\
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__25743\,
            I => \N__25740\
        );

    \I__4141\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25737\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__25737\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8\
        );

    \I__4139\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25731\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__25731\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4\
        );

    \I__4137\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25725\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__25725\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10\
        );

    \I__4135\ : CascadeMux
    port map (
            O => \N__25722\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__4134\ : InMux
    port map (
            O => \N__25719\,
            I => \N__25716\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__25716\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11\
        );

    \I__4132\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25710\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__25710\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12\
        );

    \I__4130\ : InMux
    port map (
            O => \N__25707\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__4129\ : InMux
    port map (
            O => \N__25704\,
            I => \N__25701\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__25701\,
            I => \N__25698\
        );

    \I__4127\ : Span4Mux_v
    port map (
            O => \N__25698\,
            I => \N__25695\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__25695\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__4125\ : InMux
    port map (
            O => \N__25692\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__4124\ : InMux
    port map (
            O => \N__25689\,
            I => \N__25686\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__25686\,
            I => \N__25683\
        );

    \I__4122\ : Odrv12
    port map (
            O => \N__25683\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__4121\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25677\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__25677\,
            I => \N__25674\
        );

    \I__4119\ : Odrv12
    port map (
            O => \N__25674\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__4118\ : InMux
    port map (
            O => \N__25671\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__4117\ : InMux
    port map (
            O => \N__25668\,
            I => \N__25665\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__25665\,
            I => \N__25662\
        );

    \I__4115\ : Span4Mux_h
    port map (
            O => \N__25662\,
            I => \N__25659\
        );

    \I__4114\ : Span4Mux_v
    port map (
            O => \N__25659\,
            I => \N__25656\
        );

    \I__4113\ : Odrv4
    port map (
            O => \N__25656\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__4112\ : InMux
    port map (
            O => \N__25653\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__4111\ : InMux
    port map (
            O => \N__25650\,
            I => \N__25647\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__25647\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__4109\ : InMux
    port map (
            O => \N__25644\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__4108\ : InMux
    port map (
            O => \N__25641\,
            I => \N__25638\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__25638\,
            I => \N__25635\
        );

    \I__4106\ : Odrv12
    port map (
            O => \N__25635\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__4105\ : InMux
    port map (
            O => \N__25632\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__4104\ : InMux
    port map (
            O => \N__25629\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__4103\ : InMux
    port map (
            O => \N__25626\,
            I => \N__25623\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__25623\,
            I => \N__25620\
        );

    \I__4101\ : Span4Mux_h
    port map (
            O => \N__25620\,
            I => \N__25617\
        );

    \I__4100\ : Span4Mux_v
    port map (
            O => \N__25617\,
            I => \N__25614\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__25614\,
            I => \current_shift_inst.control_input_1_axb_25\
        );

    \I__4098\ : IoInMux
    port map (
            O => \N__25611\,
            I => \N__25608\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__25608\,
            I => \N__25605\
        );

    \I__4096\ : Odrv12
    port map (
            O => \N__25605\,
            I => s4_phy_c
        );

    \I__4095\ : InMux
    port map (
            O => \N__25602\,
            I => \N__25599\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__4093\ : Odrv4
    port map (
            O => \N__25596\,
            I => \il_max_comp1_D1\
        );

    \I__4092\ : InMux
    port map (
            O => \N__25593\,
            I => \N__25590\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__25590\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\
        );

    \I__4090\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25584\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__25584\,
            I => \N__25581\
        );

    \I__4088\ : Odrv12
    port map (
            O => \N__25581\,
            I => \current_shift_inst.un38_control_input_0_s0_17\
        );

    \I__4087\ : InMux
    port map (
            O => \N__25578\,
            I => \current_shift_inst.un38_control_input_cry_16_s0\
        );

    \I__4086\ : InMux
    port map (
            O => \N__25575\,
            I => \N__25572\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__25572\,
            I => \N__25569\
        );

    \I__4084\ : Odrv12
    port map (
            O => \N__25569\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\
        );

    \I__4083\ : InMux
    port map (
            O => \N__25566\,
            I => \N__25563\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__25563\,
            I => \N__25560\
        );

    \I__4081\ : Span4Mux_v
    port map (
            O => \N__25560\,
            I => \N__25557\
        );

    \I__4080\ : Odrv4
    port map (
            O => \N__25557\,
            I => \current_shift_inst.un38_control_input_0_s0_18\
        );

    \I__4079\ : InMux
    port map (
            O => \N__25554\,
            I => \current_shift_inst.un38_control_input_cry_17_s0\
        );

    \I__4078\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25548\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__25548\,
            I => \N__25545\
        );

    \I__4076\ : Odrv12
    port map (
            O => \N__25545\,
            I => \current_shift_inst.un38_control_input_0_s0_19\
        );

    \I__4075\ : InMux
    port map (
            O => \N__25542\,
            I => \current_shift_inst.un38_control_input_cry_18_s0\
        );

    \I__4074\ : InMux
    port map (
            O => \N__25539\,
            I => \N__25536\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__25536\,
            I => \N__25533\
        );

    \I__4072\ : Odrv12
    port map (
            O => \N__25533\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__4071\ : InMux
    port map (
            O => \N__25530\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__4070\ : InMux
    port map (
            O => \N__25527\,
            I => \N__25524\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__25524\,
            I => \N__25521\
        );

    \I__4068\ : Span4Mux_v
    port map (
            O => \N__25521\,
            I => \N__25518\
        );

    \I__4067\ : Odrv4
    port map (
            O => \N__25518\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__4066\ : InMux
    port map (
            O => \N__25515\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__4065\ : InMux
    port map (
            O => \N__25512\,
            I => \N__25509\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__25509\,
            I => \N__25506\
        );

    \I__4063\ : Span4Mux_h
    port map (
            O => \N__25506\,
            I => \N__25503\
        );

    \I__4062\ : Span4Mux_v
    port map (
            O => \N__25503\,
            I => \N__25500\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__25500\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__4060\ : InMux
    port map (
            O => \N__25497\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__4059\ : InMux
    port map (
            O => \N__25494\,
            I => \N__25491\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__25491\,
            I => \N__25488\
        );

    \I__4057\ : Odrv12
    port map (
            O => \N__25488\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__4056\ : InMux
    port map (
            O => \N__25485\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__4055\ : InMux
    port map (
            O => \N__25482\,
            I => \N__25479\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__4053\ : Span4Mux_v
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__25473\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__4051\ : InMux
    port map (
            O => \N__25470\,
            I => \bfn_8_22_0_\
        );

    \I__4050\ : InMux
    port map (
            O => \N__25467\,
            I => \N__25464\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__25464\,
            I => \N__25461\
        );

    \I__4048\ : Span4Mux_v
    port map (
            O => \N__25461\,
            I => \N__25458\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__25458\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__4046\ : InMux
    port map (
            O => \N__25455\,
            I => \N__25452\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__25452\,
            I => \N__25449\
        );

    \I__4044\ : Odrv12
    port map (
            O => \N__25449\,
            I => \current_shift_inst.un38_control_input_0_s0_9\
        );

    \I__4043\ : InMux
    port map (
            O => \N__25446\,
            I => \current_shift_inst.un38_control_input_cry_8_s0\
        );

    \I__4042\ : InMux
    port map (
            O => \N__25443\,
            I => \N__25440\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__25437\,
            I => \current_shift_inst.un38_control_input_0_s0_10\
        );

    \I__4039\ : InMux
    port map (
            O => \N__25434\,
            I => \current_shift_inst.un38_control_input_cry_9_s0\
        );

    \I__4038\ : InMux
    port map (
            O => \N__25431\,
            I => \N__25428\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__25428\,
            I => \N__25425\
        );

    \I__4036\ : Odrv12
    port map (
            O => \N__25425\,
            I => \current_shift_inst.un38_control_input_0_s0_11\
        );

    \I__4035\ : InMux
    port map (
            O => \N__25422\,
            I => \current_shift_inst.un38_control_input_cry_10_s0\
        );

    \I__4034\ : InMux
    port map (
            O => \N__25419\,
            I => \N__25416\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__25416\,
            I => \N__25413\
        );

    \I__4032\ : Odrv12
    port map (
            O => \N__25413\,
            I => \current_shift_inst.un38_control_input_0_s0_12\
        );

    \I__4031\ : InMux
    port map (
            O => \N__25410\,
            I => \current_shift_inst.un38_control_input_cry_11_s0\
        );

    \I__4030\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25404\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__25401\,
            I => \current_shift_inst.un38_control_input_0_s0_13\
        );

    \I__4027\ : InMux
    port map (
            O => \N__25398\,
            I => \current_shift_inst.un38_control_input_cry_12_s0\
        );

    \I__4026\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25392\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__25392\,
            I => \N__25389\
        );

    \I__4024\ : Span4Mux_v
    port map (
            O => \N__25389\,
            I => \N__25386\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__25386\,
            I => \current_shift_inst.un38_control_input_0_s0_14\
        );

    \I__4022\ : InMux
    port map (
            O => \N__25383\,
            I => \current_shift_inst.un38_control_input_cry_13_s0\
        );

    \I__4021\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25377\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__25377\,
            I => \N__25374\
        );

    \I__4019\ : Odrv12
    port map (
            O => \N__25374\,
            I => \current_shift_inst.un38_control_input_0_s0_15\
        );

    \I__4018\ : InMux
    port map (
            O => \N__25371\,
            I => \current_shift_inst.un38_control_input_cry_14_s0\
        );

    \I__4017\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25365\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__25365\,
            I => \N__25362\
        );

    \I__4015\ : Span4Mux_v
    port map (
            O => \N__25362\,
            I => \N__25359\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__25359\,
            I => \current_shift_inst.un38_control_input_0_s0_16\
        );

    \I__4013\ : InMux
    port map (
            O => \N__25356\,
            I => \bfn_8_21_0_\
        );

    \I__4012\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25350\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__25350\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__4010\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25344\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__25344\,
            I => \N__25341\
        );

    \I__4008\ : Odrv4
    port map (
            O => \N__25341\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__4007\ : InMux
    port map (
            O => \N__25338\,
            I => \N__25335\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__25335\,
            I => \N__25332\
        );

    \I__4005\ : Odrv4
    port map (
            O => \N__25332\,
            I => \current_shift_inst.un38_control_input_0_s0_6\
        );

    \I__4004\ : InMux
    port map (
            O => \N__25329\,
            I => \current_shift_inst.un38_control_input_cry_5_s0\
        );

    \I__4003\ : InMux
    port map (
            O => \N__25326\,
            I => \N__25323\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__25323\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\
        );

    \I__4001\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25317\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__25317\,
            I => \current_shift_inst.un38_control_input_0_s0_7\
        );

    \I__3999\ : InMux
    port map (
            O => \N__25314\,
            I => \current_shift_inst.un38_control_input_cry_6_s0\
        );

    \I__3998\ : InMux
    port map (
            O => \N__25311\,
            I => \N__25308\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__25308\,
            I => \N__25305\
        );

    \I__3996\ : Span4Mux_v
    port map (
            O => \N__25305\,
            I => \N__25302\
        );

    \I__3995\ : Odrv4
    port map (
            O => \N__25302\,
            I => \current_shift_inst.un38_control_input_0_s0_8\
        );

    \I__3994\ : InMux
    port map (
            O => \N__25299\,
            I => \bfn_8_20_0_\
        );

    \I__3993\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25293\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__25293\,
            I => \N__25290\
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__25290\,
            I => \current_shift_inst.control_input_1_axb_18\
        );

    \I__3990\ : InMux
    port map (
            O => \N__25287\,
            I => \N__25284\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__25284\,
            I => \N__25281\
        );

    \I__3988\ : Odrv4
    port map (
            O => \N__25281\,
            I => \current_shift_inst.control_input_1_axb_19\
        );

    \I__3987\ : InMux
    port map (
            O => \N__25278\,
            I => \N__25275\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__25275\,
            I => \current_shift_inst.control_input_1_axb_24\
        );

    \I__3985\ : InMux
    port map (
            O => \N__25272\,
            I => \N__25269\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__25269\,
            I => \N__25266\
        );

    \I__3983\ : Span4Mux_h
    port map (
            O => \N__25266\,
            I => \N__25263\
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__25263\,
            I => \current_shift_inst.control_input_1_axb_9\
        );

    \I__3981\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25257\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__25257\,
            I => \N__25254\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__25254\,
            I => \N__25251\
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__25251\,
            I => \current_shift_inst.control_input_1_axb_1\
        );

    \I__3977\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25245\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__25245\,
            I => \N__25242\
        );

    \I__3975\ : Odrv4
    port map (
            O => \N__25242\,
            I => \current_shift_inst.control_input_1_axb_17\
        );

    \I__3974\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25236\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__25236\,
            I => \N__25233\
        );

    \I__3972\ : Span4Mux_v
    port map (
            O => \N__25233\,
            I => \N__25230\
        );

    \I__3971\ : Odrv4
    port map (
            O => \N__25230\,
            I => \current_shift_inst.control_input_1_axb_4\
        );

    \I__3970\ : InMux
    port map (
            O => \N__25227\,
            I => \N__25224\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__25224\,
            I => \N__25221\
        );

    \I__3968\ : Span4Mux_v
    port map (
            O => \N__25221\,
            I => \N__25218\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__25218\,
            I => \current_shift_inst.control_input_1_axb_7\
        );

    \I__3966\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25212\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__25212\,
            I => \current_shift_inst.control_input_1_axb_16\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__25209\,
            I => \N__25206\
        );

    \I__3963\ : InMux
    port map (
            O => \N__25206\,
            I => \N__25203\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__25203\,
            I => \current_shift_inst.control_input_1_axb_11\
        );

    \I__3961\ : InMux
    port map (
            O => \N__25200\,
            I => \N__25197\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__25197\,
            I => \current_shift_inst.control_input_1_axb_8\
        );

    \I__3959\ : InMux
    port map (
            O => \N__25194\,
            I => \N__25191\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__25191\,
            I => \N__25188\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__25188\,
            I => \current_shift_inst.control_input_1_axb_20\
        );

    \I__3956\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25182\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__25182\,
            I => \N__25179\
        );

    \I__3954\ : Span4Mux_h
    port map (
            O => \N__25179\,
            I => \N__25176\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__25176\,
            I => \current_shift_inst.control_input_1_axb_0\
        );

    \I__3952\ : InMux
    port map (
            O => \N__25173\,
            I => \N__25170\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__25170\,
            I => \current_shift_inst.control_input_1_axb_3\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__25167\,
            I => \N__25164\
        );

    \I__3949\ : InMux
    port map (
            O => \N__25164\,
            I => \N__25161\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__25161\,
            I => \N__25158\
        );

    \I__3947\ : Odrv12
    port map (
            O => \N__25158\,
            I => \phase_controller_inst2.start_timer_tr_0_sqmuxa\
        );

    \I__3946\ : InMux
    port map (
            O => \N__25155\,
            I => \N__25152\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__25152\,
            I => \current_shift_inst.control_input_1_axb_2\
        );

    \I__3944\ : InMux
    port map (
            O => \N__25149\,
            I => \N__25146\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__25146\,
            I => \current_shift_inst.control_input_1_axb_6\
        );

    \I__3942\ : InMux
    port map (
            O => \N__25143\,
            I => \N__25140\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__25140\,
            I => \current_shift_inst.control_input_1_axb_5\
        );

    \I__3940\ : InMux
    port map (
            O => \N__25137\,
            I => \N__25134\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__25134\,
            I => \current_shift_inst.control_input_1_axb_14\
        );

    \I__3938\ : InMux
    port map (
            O => \N__25131\,
            I => \N__25128\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__25128\,
            I => \current_shift_inst.control_input_1_axb_13\
        );

    \I__3936\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25122\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__25122\,
            I => \current_shift_inst.control_input_1_axb_12\
        );

    \I__3934\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25116\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__25116\,
            I => \current_shift_inst.control_input_1_axb_15\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25110\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__25110\,
            I => \current_shift_inst.control_input_1_axb_10\
        );

    \I__3930\ : InMux
    port map (
            O => \N__25107\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__25104\,
            I => \N__25101\
        );

    \I__3928\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25098\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__25098\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16\
        );

    \I__3926\ : InMux
    port map (
            O => \N__25095\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__3925\ : InMux
    port map (
            O => \N__25092\,
            I => \bfn_8_13_0_\
        );

    \I__3924\ : InMux
    port map (
            O => \N__25089\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__3923\ : InMux
    port map (
            O => \N__25086\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__3922\ : InMux
    port map (
            O => \N__25083\,
            I => \N__25080\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__25080\,
            I => \N__25077\
        );

    \I__3920\ : Odrv4
    port map (
            O => \N__25077\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0\
        );

    \I__3919\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25071\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__25071\,
            I => \N__25068\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__25068\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__3916\ : InMux
    port map (
            O => \N__25065\,
            I => \N__25062\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__25062\,
            I => \current_shift_inst.control_input_1_axb_22\
        );

    \I__3914\ : InMux
    port map (
            O => \N__25059\,
            I => \N__25056\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__25056\,
            I => \current_shift_inst.control_input_1_axb_21\
        );

    \I__3912\ : InMux
    port map (
            O => \N__25053\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__3911\ : InMux
    port map (
            O => \N__25050\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__3910\ : InMux
    port map (
            O => \N__25047\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__3909\ : InMux
    port map (
            O => \N__25044\,
            I => \bfn_8_12_0_\
        );

    \I__3908\ : InMux
    port map (
            O => \N__25041\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__3907\ : InMux
    port map (
            O => \N__25038\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__3906\ : InMux
    port map (
            O => \N__25035\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__3905\ : InMux
    port map (
            O => \N__25032\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__3904\ : InMux
    port map (
            O => \N__25029\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__3903\ : InMux
    port map (
            O => \N__25026\,
            I => \N__25023\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__25023\,
            I => \N__25020\
        );

    \I__3901\ : Odrv4
    port map (
            O => \N__25020\,
            I => \il_min_comp2_D1\
        );

    \I__3900\ : InMux
    port map (
            O => \N__25017\,
            I => \N__25012\
        );

    \I__3899\ : InMux
    port map (
            O => \N__25016\,
            I => \N__25009\
        );

    \I__3898\ : InMux
    port map (
            O => \N__25015\,
            I => \N__25006\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__25012\,
            I => \N__25003\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__25009\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__25006\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__25003\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__3893\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24992\
        );

    \I__3892\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24989\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__24992\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__24989\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3889\ : InMux
    port map (
            O => \N__24984\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__3888\ : InMux
    port map (
            O => \N__24981\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__3887\ : InMux
    port map (
            O => \N__24978\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__3886\ : InMux
    port map (
            O => \N__24975\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__3885\ : CascadeMux
    port map (
            O => \N__24972\,
            I => \N__24968\
        );

    \I__3884\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24965\
        );

    \I__3883\ : InMux
    port map (
            O => \N__24968\,
            I => \N__24962\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__24965\,
            I => \N__24959\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__24962\,
            I => \N__24956\
        );

    \I__3880\ : Span4Mux_h
    port map (
            O => \N__24959\,
            I => \N__24953\
        );

    \I__3879\ : Span4Mux_h
    port map (
            O => \N__24956\,
            I => \N__24950\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__24953\,
            I => \current_shift_inst.control_inputZ0Z_23\
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__24950\,
            I => \current_shift_inst.control_inputZ0Z_23\
        );

    \I__3876\ : InMux
    port map (
            O => \N__24945\,
            I => \current_shift_inst.control_input_1_cry_22\
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__24942\,
            I => \N__24938\
        );

    \I__3874\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24935\
        );

    \I__3873\ : InMux
    port map (
            O => \N__24938\,
            I => \N__24932\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__24935\,
            I => \N__24927\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__24932\,
            I => \N__24927\
        );

    \I__3870\ : Odrv12
    port map (
            O => \N__24927\,
            I => \current_shift_inst.control_inputZ0Z_24\
        );

    \I__3869\ : InMux
    port map (
            O => \N__24924\,
            I => \bfn_7_16_0_\
        );

    \I__3868\ : InMux
    port map (
            O => \N__24921\,
            I => \current_shift_inst.control_input_1_cry_24\
        );

    \I__3867\ : CascadeMux
    port map (
            O => \N__24918\,
            I => \N__24910\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__24917\,
            I => \N__24906\
        );

    \I__3865\ : CascadeMux
    port map (
            O => \N__24916\,
            I => \N__24902\
        );

    \I__3864\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24899\
        );

    \I__3863\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24884\
        );

    \I__3862\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24884\
        );

    \I__3861\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24884\
        );

    \I__3860\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24884\
        );

    \I__3859\ : InMux
    port map (
            O => \N__24906\,
            I => \N__24884\
        );

    \I__3858\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24884\
        );

    \I__3857\ : InMux
    port map (
            O => \N__24902\,
            I => \N__24884\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__24899\,
            I => \N__24879\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__24884\,
            I => \N__24879\
        );

    \I__3854\ : Span4Mux_h
    port map (
            O => \N__24879\,
            I => \N__24876\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__24876\,
            I => \current_shift_inst.control_inputZ0Z_25\
        );

    \I__3852\ : CEMux
    port map (
            O => \N__24873\,
            I => \N__24868\
        );

    \I__3851\ : CEMux
    port map (
            O => \N__24872\,
            I => \N__24863\
        );

    \I__3850\ : CEMux
    port map (
            O => \N__24871\,
            I => \N__24858\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__24868\,
            I => \N__24853\
        );

    \I__3848\ : CEMux
    port map (
            O => \N__24867\,
            I => \N__24850\
        );

    \I__3847\ : CEMux
    port map (
            O => \N__24866\,
            I => \N__24847\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__24863\,
            I => \N__24842\
        );

    \I__3845\ : CEMux
    port map (
            O => \N__24862\,
            I => \N__24839\
        );

    \I__3844\ : CEMux
    port map (
            O => \N__24861\,
            I => \N__24836\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__24858\,
            I => \N__24833\
        );

    \I__3842\ : CEMux
    port map (
            O => \N__24857\,
            I => \N__24830\
        );

    \I__3841\ : CEMux
    port map (
            O => \N__24856\,
            I => \N__24827\
        );

    \I__3840\ : Span4Mux_h
    port map (
            O => \N__24853\,
            I => \N__24816\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__24850\,
            I => \N__24816\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__24847\,
            I => \N__24813\
        );

    \I__3837\ : CEMux
    port map (
            O => \N__24846\,
            I => \N__24809\
        );

    \I__3836\ : CEMux
    port map (
            O => \N__24845\,
            I => \N__24806\
        );

    \I__3835\ : Span4Mux_v
    port map (
            O => \N__24842\,
            I => \N__24800\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__24839\,
            I => \N__24800\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__24836\,
            I => \N__24797\
        );

    \I__3832\ : Span4Mux_v
    port map (
            O => \N__24833\,
            I => \N__24790\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__24830\,
            I => \N__24790\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__24827\,
            I => \N__24790\
        );

    \I__3829\ : CEMux
    port map (
            O => \N__24826\,
            I => \N__24787\
        );

    \I__3828\ : CEMux
    port map (
            O => \N__24825\,
            I => \N__24782\
        );

    \I__3827\ : CEMux
    port map (
            O => \N__24824\,
            I => \N__24779\
        );

    \I__3826\ : CEMux
    port map (
            O => \N__24823\,
            I => \N__24776\
        );

    \I__3825\ : CEMux
    port map (
            O => \N__24822\,
            I => \N__24771\
        );

    \I__3824\ : CEMux
    port map (
            O => \N__24821\,
            I => \N__24767\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__24816\,
            I => \N__24763\
        );

    \I__3822\ : Span4Mux_h
    port map (
            O => \N__24813\,
            I => \N__24760\
        );

    \I__3821\ : CEMux
    port map (
            O => \N__24812\,
            I => \N__24757\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24752\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__24806\,
            I => \N__24752\
        );

    \I__3818\ : CEMux
    port map (
            O => \N__24805\,
            I => \N__24749\
        );

    \I__3817\ : Span4Mux_v
    port map (
            O => \N__24800\,
            I => \N__24739\
        );

    \I__3816\ : Span4Mux_h
    port map (
            O => \N__24797\,
            I => \N__24739\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__24790\,
            I => \N__24739\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__24787\,
            I => \N__24739\
        );

    \I__3813\ : CEMux
    port map (
            O => \N__24786\,
            I => \N__24736\
        );

    \I__3812\ : CEMux
    port map (
            O => \N__24785\,
            I => \N__24733\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__24782\,
            I => \N__24729\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24726\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__24776\,
            I => \N__24723\
        );

    \I__3808\ : CEMux
    port map (
            O => \N__24775\,
            I => \N__24720\
        );

    \I__3807\ : CEMux
    port map (
            O => \N__24774\,
            I => \N__24717\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__24771\,
            I => \N__24713\
        );

    \I__3805\ : CEMux
    port map (
            O => \N__24770\,
            I => \N__24710\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__24767\,
            I => \N__24707\
        );

    \I__3803\ : CEMux
    port map (
            O => \N__24766\,
            I => \N__24704\
        );

    \I__3802\ : Span4Mux_v
    port map (
            O => \N__24763\,
            I => \N__24700\
        );

    \I__3801\ : Span4Mux_v
    port map (
            O => \N__24760\,
            I => \N__24695\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__24757\,
            I => \N__24695\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__24752\,
            I => \N__24690\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__24749\,
            I => \N__24690\
        );

    \I__3797\ : CEMux
    port map (
            O => \N__24748\,
            I => \N__24687\
        );

    \I__3796\ : Span4Mux_h
    port map (
            O => \N__24739\,
            I => \N__24682\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__24736\,
            I => \N__24682\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__24733\,
            I => \N__24679\
        );

    \I__3793\ : CEMux
    port map (
            O => \N__24732\,
            I => \N__24676\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__24729\,
            I => \N__24673\
        );

    \I__3791\ : Span4Mux_h
    port map (
            O => \N__24726\,
            I => \N__24664\
        );

    \I__3790\ : Span4Mux_v
    port map (
            O => \N__24723\,
            I => \N__24664\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__24720\,
            I => \N__24664\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__24717\,
            I => \N__24664\
        );

    \I__3787\ : CEMux
    port map (
            O => \N__24716\,
            I => \N__24661\
        );

    \I__3786\ : Span4Mux_h
    port map (
            O => \N__24713\,
            I => \N__24652\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__24710\,
            I => \N__24652\
        );

    \I__3784\ : Span4Mux_v
    port map (
            O => \N__24707\,
            I => \N__24652\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__24704\,
            I => \N__24652\
        );

    \I__3782\ : CEMux
    port map (
            O => \N__24703\,
            I => \N__24649\
        );

    \I__3781\ : Span4Mux_v
    port map (
            O => \N__24700\,
            I => \N__24646\
        );

    \I__3780\ : Span4Mux_h
    port map (
            O => \N__24695\,
            I => \N__24643\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__24690\,
            I => \N__24640\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__24687\,
            I => \N__24637\
        );

    \I__3777\ : Span4Mux_v
    port map (
            O => \N__24682\,
            I => \N__24634\
        );

    \I__3776\ : Span4Mux_v
    port map (
            O => \N__24679\,
            I => \N__24629\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__24676\,
            I => \N__24629\
        );

    \I__3774\ : Span4Mux_h
    port map (
            O => \N__24673\,
            I => \N__24622\
        );

    \I__3773\ : Span4Mux_v
    port map (
            O => \N__24664\,
            I => \N__24622\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__24661\,
            I => \N__24622\
        );

    \I__3771\ : Span4Mux_v
    port map (
            O => \N__24652\,
            I => \N__24617\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__24649\,
            I => \N__24617\
        );

    \I__3769\ : Span4Mux_h
    port map (
            O => \N__24646\,
            I => \N__24614\
        );

    \I__3768\ : Span4Mux_v
    port map (
            O => \N__24643\,
            I => \N__24609\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__24640\,
            I => \N__24609\
        );

    \I__3766\ : Span4Mux_h
    port map (
            O => \N__24637\,
            I => \N__24606\
        );

    \I__3765\ : Span4Mux_s2_h
    port map (
            O => \N__24634\,
            I => \N__24601\
        );

    \I__3764\ : Span4Mux_v
    port map (
            O => \N__24629\,
            I => \N__24601\
        );

    \I__3763\ : Span4Mux_v
    port map (
            O => \N__24622\,
            I => \N__24596\
        );

    \I__3762\ : Span4Mux_h
    port map (
            O => \N__24617\,
            I => \N__24596\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__24614\,
            I => \N_748_g\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__24609\,
            I => \N_748_g\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__24606\,
            I => \N_748_g\
        );

    \I__3758\ : Odrv4
    port map (
            O => \N__24601\,
            I => \N_748_g\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__24596\,
            I => \N_748_g\
        );

    \I__3756\ : InMux
    port map (
            O => \N__24585\,
            I => \N__24582\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__24582\,
            I => \N__24579\
        );

    \I__3754\ : Sp12to4
    port map (
            O => \N__24579\,
            I => \N__24576\
        );

    \I__3753\ : Odrv12
    port map (
            O => \N__24576\,
            I => \current_shift_inst.control_input_1_axb_23\
        );

    \I__3752\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24570\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__24570\,
            I => \N__24567\
        );

    \I__3750\ : Odrv12
    port map (
            O => \N__24567\,
            I => il_max_comp1_c
        );

    \I__3749\ : InMux
    port map (
            O => \N__24564\,
            I => \N__24561\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__24561\,
            I => \N__24558\
        );

    \I__3747\ : Span4Mux_h
    port map (
            O => \N__24558\,
            I => \N__24555\
        );

    \I__3746\ : Span4Mux_v
    port map (
            O => \N__24555\,
            I => \N__24552\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__24552\,
            I => il_min_comp2_c
        );

    \I__3744\ : InMux
    port map (
            O => \N__24549\,
            I => \N__24545\
        );

    \I__3743\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24542\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__24545\,
            I => \N__24537\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__24542\,
            I => \N__24537\
        );

    \I__3740\ : Span4Mux_h
    port map (
            O => \N__24537\,
            I => \N__24534\
        );

    \I__3739\ : Odrv4
    port map (
            O => \N__24534\,
            I => \current_shift_inst.control_inputZ0Z_15\
        );

    \I__3738\ : InMux
    port map (
            O => \N__24531\,
            I => \current_shift_inst.control_input_1_cry_14\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__24528\,
            I => \N__24524\
        );

    \I__3736\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24521\
        );

    \I__3735\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24518\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__24521\,
            I => \N__24515\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__24518\,
            I => \N__24512\
        );

    \I__3732\ : Span4Mux_h
    port map (
            O => \N__24515\,
            I => \N__24509\
        );

    \I__3731\ : Span4Mux_h
    port map (
            O => \N__24512\,
            I => \N__24506\
        );

    \I__3730\ : Odrv4
    port map (
            O => \N__24509\,
            I => \current_shift_inst.control_inputZ0Z_16\
        );

    \I__3729\ : Odrv4
    port map (
            O => \N__24506\,
            I => \current_shift_inst.control_inputZ0Z_16\
        );

    \I__3728\ : InMux
    port map (
            O => \N__24501\,
            I => \bfn_7_15_0_\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__24498\,
            I => \N__24494\
        );

    \I__3726\ : InMux
    port map (
            O => \N__24497\,
            I => \N__24491\
        );

    \I__3725\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24488\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24483\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__24488\,
            I => \N__24483\
        );

    \I__3722\ : Odrv12
    port map (
            O => \N__24483\,
            I => \current_shift_inst.control_inputZ0Z_17\
        );

    \I__3721\ : InMux
    port map (
            O => \N__24480\,
            I => \current_shift_inst.control_input_1_cry_16\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__24477\,
            I => \N__24473\
        );

    \I__3719\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24470\
        );

    \I__3718\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24467\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__24470\,
            I => \N__24464\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__24467\,
            I => \N__24461\
        );

    \I__3715\ : Odrv12
    port map (
            O => \N__24464\,
            I => \current_shift_inst.control_inputZ0Z_18\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__24461\,
            I => \current_shift_inst.control_inputZ0Z_18\
        );

    \I__3713\ : InMux
    port map (
            O => \N__24456\,
            I => \current_shift_inst.control_input_1_cry_17\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__24453\,
            I => \N__24449\
        );

    \I__3711\ : InMux
    port map (
            O => \N__24452\,
            I => \N__24446\
        );

    \I__3710\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24443\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__24446\,
            I => \N__24438\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__24443\,
            I => \N__24438\
        );

    \I__3707\ : Odrv12
    port map (
            O => \N__24438\,
            I => \current_shift_inst.control_inputZ0Z_19\
        );

    \I__3706\ : InMux
    port map (
            O => \N__24435\,
            I => \current_shift_inst.control_input_1_cry_18\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__24432\,
            I => \N__24428\
        );

    \I__3704\ : InMux
    port map (
            O => \N__24431\,
            I => \N__24425\
        );

    \I__3703\ : InMux
    port map (
            O => \N__24428\,
            I => \N__24422\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__24425\,
            I => \N__24419\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__24422\,
            I => \N__24416\
        );

    \I__3700\ : Odrv12
    port map (
            O => \N__24419\,
            I => \current_shift_inst.control_inputZ0Z_20\
        );

    \I__3699\ : Odrv4
    port map (
            O => \N__24416\,
            I => \current_shift_inst.control_inputZ0Z_20\
        );

    \I__3698\ : InMux
    port map (
            O => \N__24411\,
            I => \current_shift_inst.control_input_1_cry_19\
        );

    \I__3697\ : InMux
    port map (
            O => \N__24408\,
            I => \N__24404\
        );

    \I__3696\ : CascadeMux
    port map (
            O => \N__24407\,
            I => \N__24401\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__24404\,
            I => \N__24398\
        );

    \I__3694\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24395\
        );

    \I__3693\ : Span4Mux_v
    port map (
            O => \N__24398\,
            I => \N__24390\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__24395\,
            I => \N__24390\
        );

    \I__3691\ : Odrv4
    port map (
            O => \N__24390\,
            I => \current_shift_inst.control_inputZ0Z_21\
        );

    \I__3690\ : InMux
    port map (
            O => \N__24387\,
            I => \current_shift_inst.control_input_1_cry_20\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__24384\,
            I => \N__24380\
        );

    \I__3688\ : InMux
    port map (
            O => \N__24383\,
            I => \N__24377\
        );

    \I__3687\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24374\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__24377\,
            I => \N__24369\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__24374\,
            I => \N__24369\
        );

    \I__3684\ : Odrv12
    port map (
            O => \N__24369\,
            I => \current_shift_inst.control_inputZ0Z_22\
        );

    \I__3683\ : InMux
    port map (
            O => \N__24366\,
            I => \current_shift_inst.control_input_1_cry_21\
        );

    \I__3682\ : CascadeMux
    port map (
            O => \N__24363\,
            I => \N__24359\
        );

    \I__3681\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24356\
        );

    \I__3680\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24353\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__24356\,
            I => \N__24348\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__24353\,
            I => \N__24348\
        );

    \I__3677\ : Span4Mux_h
    port map (
            O => \N__24348\,
            I => \N__24345\
        );

    \I__3676\ : Odrv4
    port map (
            O => \N__24345\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__3675\ : InMux
    port map (
            O => \N__24342\,
            I => \current_shift_inst.control_input_1_cry_5\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__24339\,
            I => \N__24335\
        );

    \I__3673\ : InMux
    port map (
            O => \N__24338\,
            I => \N__24332\
        );

    \I__3672\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24329\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__24332\,
            I => \N__24324\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24324\
        );

    \I__3669\ : Span4Mux_h
    port map (
            O => \N__24324\,
            I => \N__24321\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__24321\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__3667\ : InMux
    port map (
            O => \N__24318\,
            I => \current_shift_inst.control_input_1_cry_6\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__24315\,
            I => \N__24311\
        );

    \I__3665\ : InMux
    port map (
            O => \N__24314\,
            I => \N__24308\
        );

    \I__3664\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24305\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__24308\,
            I => \N__24300\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24300\
        );

    \I__3661\ : Span4Mux_h
    port map (
            O => \N__24300\,
            I => \N__24297\
        );

    \I__3660\ : Odrv4
    port map (
            O => \N__24297\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__3659\ : InMux
    port map (
            O => \N__24294\,
            I => \bfn_7_14_0_\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__24291\,
            I => \N__24287\
        );

    \I__3657\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24284\
        );

    \I__3656\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24281\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__24284\,
            I => \N__24276\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__24281\,
            I => \N__24276\
        );

    \I__3653\ : Span4Mux_h
    port map (
            O => \N__24276\,
            I => \N__24273\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__24273\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__3651\ : InMux
    port map (
            O => \N__24270\,
            I => \current_shift_inst.control_input_1_cry_8\
        );

    \I__3650\ : InMux
    port map (
            O => \N__24267\,
            I => \N__24263\
        );

    \I__3649\ : CascadeMux
    port map (
            O => \N__24266\,
            I => \N__24260\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__24263\,
            I => \N__24257\
        );

    \I__3647\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24254\
        );

    \I__3646\ : Span4Mux_v
    port map (
            O => \N__24257\,
            I => \N__24249\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__24254\,
            I => \N__24249\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__24249\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__3643\ : InMux
    port map (
            O => \N__24246\,
            I => \current_shift_inst.control_input_1_cry_9\
        );

    \I__3642\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24239\
        );

    \I__3641\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24236\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__24239\,
            I => \N__24231\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__24236\,
            I => \N__24231\
        );

    \I__3638\ : Span4Mux_h
    port map (
            O => \N__24231\,
            I => \N__24228\
        );

    \I__3637\ : Odrv4
    port map (
            O => \N__24228\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__3636\ : InMux
    port map (
            O => \N__24225\,
            I => \current_shift_inst.control_input_1_cry_10\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__24222\,
            I => \N__24218\
        );

    \I__3634\ : InMux
    port map (
            O => \N__24221\,
            I => \N__24215\
        );

    \I__3633\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24212\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__24215\,
            I => \N__24209\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__24212\,
            I => \N__24206\
        );

    \I__3630\ : Odrv12
    port map (
            O => \N__24209\,
            I => \current_shift_inst.control_inputZ0Z_12\
        );

    \I__3629\ : Odrv4
    port map (
            O => \N__24206\,
            I => \current_shift_inst.control_inputZ0Z_12\
        );

    \I__3628\ : InMux
    port map (
            O => \N__24201\,
            I => \current_shift_inst.control_input_1_cry_11\
        );

    \I__3627\ : InMux
    port map (
            O => \N__24198\,
            I => \N__24194\
        );

    \I__3626\ : CascadeMux
    port map (
            O => \N__24197\,
            I => \N__24191\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__24194\,
            I => \N__24188\
        );

    \I__3624\ : InMux
    port map (
            O => \N__24191\,
            I => \N__24185\
        );

    \I__3623\ : Span4Mux_v
    port map (
            O => \N__24188\,
            I => \N__24180\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__24185\,
            I => \N__24180\
        );

    \I__3621\ : Odrv4
    port map (
            O => \N__24180\,
            I => \current_shift_inst.control_inputZ0Z_13\
        );

    \I__3620\ : InMux
    port map (
            O => \N__24177\,
            I => \current_shift_inst.control_input_1_cry_12\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__24174\,
            I => \N__24170\
        );

    \I__3618\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24167\
        );

    \I__3617\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24164\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__24167\,
            I => \N__24159\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__24164\,
            I => \N__24159\
        );

    \I__3614\ : Odrv12
    port map (
            O => \N__24159\,
            I => \current_shift_inst.control_inputZ0Z_14\
        );

    \I__3613\ : InMux
    port map (
            O => \N__24156\,
            I => \current_shift_inst.control_input_1_cry_13\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__24153\,
            I => \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa_cascade_\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__24150\,
            I => \N__24147\
        );

    \I__3610\ : InMux
    port map (
            O => \N__24147\,
            I => \N__24144\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__24144\,
            I => \N__24141\
        );

    \I__3608\ : Span4Mux_s3_h
    port map (
            O => \N__24141\,
            I => \N__24138\
        );

    \I__3607\ : Span4Mux_h
    port map (
            O => \N__24138\,
            I => \N__24135\
        );

    \I__3606\ : Odrv4
    port map (
            O => \N__24135\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__3605\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24128\
        );

    \I__3604\ : CascadeMux
    port map (
            O => \N__24131\,
            I => \N__24124\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__24128\,
            I => \N__24121\
        );

    \I__3602\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24118\
        );

    \I__3601\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24115\
        );

    \I__3600\ : Span4Mux_v
    port map (
            O => \N__24121\,
            I => \N__24112\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__24118\,
            I => \N__24107\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__24115\,
            I => \N__24107\
        );

    \I__3597\ : Span4Mux_h
    port map (
            O => \N__24112\,
            I => \N__24104\
        );

    \I__3596\ : Span4Mux_h
    port map (
            O => \N__24107\,
            I => \N__24101\
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__24104\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__24101\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__3593\ : CascadeMux
    port map (
            O => \N__24096\,
            I => \N__24092\
        );

    \I__3592\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24089\
        );

    \I__3591\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24086\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__24089\,
            I => \N__24081\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__24086\,
            I => \N__24081\
        );

    \I__3588\ : Span4Mux_h
    port map (
            O => \N__24081\,
            I => \N__24078\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__24078\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__3586\ : InMux
    port map (
            O => \N__24075\,
            I => \current_shift_inst.control_input_1_cry_0\
        );

    \I__3585\ : CascadeMux
    port map (
            O => \N__24072\,
            I => \N__24069\
        );

    \I__3584\ : InMux
    port map (
            O => \N__24069\,
            I => \N__24065\
        );

    \I__3583\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24062\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__24065\,
            I => \N__24059\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__24062\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__3580\ : Odrv12
    port map (
            O => \N__24059\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__3579\ : InMux
    port map (
            O => \N__24054\,
            I => \current_shift_inst.control_input_1_cry_1\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__24051\,
            I => \N__24047\
        );

    \I__3577\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24044\
        );

    \I__3576\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24041\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__24044\,
            I => \N__24036\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__24041\,
            I => \N__24036\
        );

    \I__3573\ : Odrv12
    port map (
            O => \N__24036\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__3572\ : InMux
    port map (
            O => \N__24033\,
            I => \current_shift_inst.control_input_1_cry_2\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__24030\,
            I => \N__24026\
        );

    \I__3570\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24023\
        );

    \I__3569\ : InMux
    port map (
            O => \N__24026\,
            I => \N__24020\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__24023\,
            I => \N__24015\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__24020\,
            I => \N__24015\
        );

    \I__3566\ : Odrv12
    port map (
            O => \N__24015\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__3565\ : InMux
    port map (
            O => \N__24012\,
            I => \current_shift_inst.control_input_1_cry_3\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__24009\,
            I => \N__24005\
        );

    \I__3563\ : InMux
    port map (
            O => \N__24008\,
            I => \N__24002\
        );

    \I__3562\ : InMux
    port map (
            O => \N__24005\,
            I => \N__23999\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__24002\,
            I => \N__23996\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__23999\,
            I => \N__23993\
        );

    \I__3559\ : Odrv12
    port map (
            O => \N__23996\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__3558\ : Odrv4
    port map (
            O => \N__23993\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__3557\ : InMux
    port map (
            O => \N__23988\,
            I => \current_shift_inst.control_input_1_cry_4\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__23985\,
            I => \N__23982\
        );

    \I__3555\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23979\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__23979\,
            I => \N__23975\
        );

    \I__3553\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23970\
        );

    \I__3552\ : Span4Mux_v
    port map (
            O => \N__23975\,
            I => \N__23967\
        );

    \I__3551\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23964\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__23973\,
            I => \N__23961\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__23970\,
            I => \N__23958\
        );

    \I__3548\ : Span4Mux_h
    port map (
            O => \N__23967\,
            I => \N__23953\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__23964\,
            I => \N__23953\
        );

    \I__3546\ : InMux
    port map (
            O => \N__23961\,
            I => \N__23950\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__23958\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__23953\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__23950\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__23943\,
            I => \N__23940\
        );

    \I__3541\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23937\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__23937\,
            I => \N__23934\
        );

    \I__3539\ : Span4Mux_h
    port map (
            O => \N__23934\,
            I => \N__23931\
        );

    \I__3538\ : Odrv4
    port map (
            O => \N__23931\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__3537\ : InMux
    port map (
            O => \N__23928\,
            I => \N__23925\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__23925\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__23922\,
            I => \N__23911\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__23921\,
            I => \N__23908\
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__23920\,
            I => \N__23902\
        );

    \I__3532\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23892\
        );

    \I__3531\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23892\
        );

    \I__3530\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23889\
        );

    \I__3529\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23882\
        );

    \I__3528\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23882\
        );

    \I__3527\ : InMux
    port map (
            O => \N__23914\,
            I => \N__23882\
        );

    \I__3526\ : InMux
    port map (
            O => \N__23911\,
            I => \N__23871\
        );

    \I__3525\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23871\
        );

    \I__3524\ : InMux
    port map (
            O => \N__23907\,
            I => \N__23871\
        );

    \I__3523\ : InMux
    port map (
            O => \N__23906\,
            I => \N__23871\
        );

    \I__3522\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23871\
        );

    \I__3521\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23855\
        );

    \I__3520\ : InMux
    port map (
            O => \N__23901\,
            I => \N__23855\
        );

    \I__3519\ : InMux
    port map (
            O => \N__23900\,
            I => \N__23855\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__23899\,
            I => \N__23852\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__23898\,
            I => \N__23848\
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__23897\,
            I => \N__23845\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__23892\,
            I => \N__23834\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__23889\,
            I => \N__23834\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__23882\,
            I => \N__23834\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__23871\,
            I => \N__23834\
        );

    \I__3511\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23827\
        );

    \I__3510\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23827\
        );

    \I__3509\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23827\
        );

    \I__3508\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23818\
        );

    \I__3507\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23818\
        );

    \I__3506\ : InMux
    port map (
            O => \N__23865\,
            I => \N__23818\
        );

    \I__3505\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23818\
        );

    \I__3504\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23815\
        );

    \I__3503\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23812\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__23855\,
            I => \N__23809\
        );

    \I__3501\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23796\
        );

    \I__3500\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23796\
        );

    \I__3499\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23796\
        );

    \I__3498\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23796\
        );

    \I__3497\ : InMux
    port map (
            O => \N__23844\,
            I => \N__23796\
        );

    \I__3496\ : InMux
    port map (
            O => \N__23843\,
            I => \N__23796\
        );

    \I__3495\ : Span4Mux_v
    port map (
            O => \N__23834\,
            I => \N__23785\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__23827\,
            I => \N__23785\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__23818\,
            I => \N__23785\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__23815\,
            I => \N__23785\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__23812\,
            I => \N__23782\
        );

    \I__3490\ : Span4Mux_v
    port map (
            O => \N__23809\,
            I => \N__23777\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__23796\,
            I => \N__23777\
        );

    \I__3488\ : InMux
    port map (
            O => \N__23795\,
            I => \N__23774\
        );

    \I__3487\ : InMux
    port map (
            O => \N__23794\,
            I => \N__23771\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__23785\,
            I => \current_shift_inst.PI_CTRL.N_170\
        );

    \I__3485\ : Odrv4
    port map (
            O => \N__23782\,
            I => \current_shift_inst.PI_CTRL.N_170\
        );

    \I__3484\ : Odrv4
    port map (
            O => \N__23777\,
            I => \current_shift_inst.PI_CTRL.N_170\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__23774\,
            I => \current_shift_inst.PI_CTRL.N_170\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__23771\,
            I => \current_shift_inst.PI_CTRL.N_170\
        );

    \I__3481\ : InMux
    port map (
            O => \N__23760\,
            I => \N__23748\
        );

    \I__3480\ : InMux
    port map (
            O => \N__23759\,
            I => \N__23748\
        );

    \I__3479\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23748\
        );

    \I__3478\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23742\
        );

    \I__3477\ : InMux
    port map (
            O => \N__23756\,
            I => \N__23737\
        );

    \I__3476\ : InMux
    port map (
            O => \N__23755\,
            I => \N__23737\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__23748\,
            I => \N__23725\
        );

    \I__3474\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23720\
        );

    \I__3473\ : InMux
    port map (
            O => \N__23746\,
            I => \N__23720\
        );

    \I__3472\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23717\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__23742\,
            I => \N__23714\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__23737\,
            I => \N__23711\
        );

    \I__3469\ : InMux
    port map (
            O => \N__23736\,
            I => \N__23702\
        );

    \I__3468\ : InMux
    port map (
            O => \N__23735\,
            I => \N__23702\
        );

    \I__3467\ : InMux
    port map (
            O => \N__23734\,
            I => \N__23702\
        );

    \I__3466\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23702\
        );

    \I__3465\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23691\
        );

    \I__3464\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23691\
        );

    \I__3463\ : InMux
    port map (
            O => \N__23730\,
            I => \N__23691\
        );

    \I__3462\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23691\
        );

    \I__3461\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23691\
        );

    \I__3460\ : Span4Mux_h
    port map (
            O => \N__23725\,
            I => \N__23675\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__23720\,
            I => \N__23670\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__23717\,
            I => \N__23670\
        );

    \I__3457\ : Span4Mux_v
    port map (
            O => \N__23714\,
            I => \N__23661\
        );

    \I__3456\ : Span4Mux_v
    port map (
            O => \N__23711\,
            I => \N__23661\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__23702\,
            I => \N__23661\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23661\
        );

    \I__3453\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23648\
        );

    \I__3452\ : InMux
    port map (
            O => \N__23689\,
            I => \N__23648\
        );

    \I__3451\ : InMux
    port map (
            O => \N__23688\,
            I => \N__23648\
        );

    \I__3450\ : InMux
    port map (
            O => \N__23687\,
            I => \N__23648\
        );

    \I__3449\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23648\
        );

    \I__3448\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23648\
        );

    \I__3447\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23633\
        );

    \I__3446\ : InMux
    port map (
            O => \N__23683\,
            I => \N__23633\
        );

    \I__3445\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23633\
        );

    \I__3444\ : InMux
    port map (
            O => \N__23681\,
            I => \N__23633\
        );

    \I__3443\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23633\
        );

    \I__3442\ : InMux
    port map (
            O => \N__23679\,
            I => \N__23633\
        );

    \I__3441\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23633\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__23675\,
            I => \current_shift_inst.PI_CTRL.N_171\
        );

    \I__3439\ : Odrv4
    port map (
            O => \N__23670\,
            I => \current_shift_inst.PI_CTRL.N_171\
        );

    \I__3438\ : Odrv4
    port map (
            O => \N__23661\,
            I => \current_shift_inst.PI_CTRL.N_171\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__23648\,
            I => \current_shift_inst.PI_CTRL.N_171\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__23633\,
            I => \current_shift_inst.PI_CTRL.N_171\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__23622\,
            I => \N__23614\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__23621\,
            I => \N__23607\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__23620\,
            I => \N__23604\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__23619\,
            I => \N__23596\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__23618\,
            I => \N__23593\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__23617\,
            I => \N__23590\
        );

    \I__3429\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23585\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__23613\,
            I => \N__23576\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__23612\,
            I => \N__23573\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__23611\,
            I => \N__23570\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__23610\,
            I => \N__23567\
        );

    \I__3424\ : InMux
    port map (
            O => \N__23607\,
            I => \N__23558\
        );

    \I__3423\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23558\
        );

    \I__3422\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23558\
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__23602\,
            I => \N__23554\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__23601\,
            I => \N__23551\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__23600\,
            I => \N__23548\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__23599\,
            I => \N__23545\
        );

    \I__3417\ : InMux
    port map (
            O => \N__23596\,
            I => \N__23539\
        );

    \I__3416\ : InMux
    port map (
            O => \N__23593\,
            I => \N__23532\
        );

    \I__3415\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23532\
        );

    \I__3414\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23532\
        );

    \I__3413\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23529\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__23585\,
            I => \N__23526\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__23584\,
            I => \N__23521\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__23583\,
            I => \N__23518\
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__23582\,
            I => \N__23515\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__23581\,
            I => \N__23512\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__23580\,
            I => \N__23509\
        );

    \I__3406\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23505\
        );

    \I__3405\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23502\
        );

    \I__3404\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23491\
        );

    \I__3403\ : InMux
    port map (
            O => \N__23570\,
            I => \N__23491\
        );

    \I__3402\ : InMux
    port map (
            O => \N__23567\,
            I => \N__23491\
        );

    \I__3401\ : InMux
    port map (
            O => \N__23566\,
            I => \N__23491\
        );

    \I__3400\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23491\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__23558\,
            I => \N__23488\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__23557\,
            I => \N__23485\
        );

    \I__3397\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23472\
        );

    \I__3396\ : InMux
    port map (
            O => \N__23551\,
            I => \N__23472\
        );

    \I__3395\ : InMux
    port map (
            O => \N__23548\,
            I => \N__23472\
        );

    \I__3394\ : InMux
    port map (
            O => \N__23545\,
            I => \N__23472\
        );

    \I__3393\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23472\
        );

    \I__3392\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23472\
        );

    \I__3391\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23469\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__23539\,
            I => \N__23460\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__23532\,
            I => \N__23460\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__23529\,
            I => \N__23460\
        );

    \I__3387\ : Span4Mux_h
    port map (
            O => \N__23526\,
            I => \N__23460\
        );

    \I__3386\ : InMux
    port map (
            O => \N__23525\,
            I => \N__23457\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__23524\,
            I => \N__23454\
        );

    \I__3384\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23449\
        );

    \I__3383\ : InMux
    port map (
            O => \N__23518\,
            I => \N__23449\
        );

    \I__3382\ : InMux
    port map (
            O => \N__23515\,
            I => \N__23440\
        );

    \I__3381\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23440\
        );

    \I__3380\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23440\
        );

    \I__3379\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23440\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__23505\,
            I => \N__23437\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__23502\,
            I => \N__23432\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__23491\,
            I => \N__23432\
        );

    \I__3375\ : Span4Mux_h
    port map (
            O => \N__23488\,
            I => \N__23429\
        );

    \I__3374\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23426\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__23472\,
            I => \N__23417\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__23469\,
            I => \N__23417\
        );

    \I__3371\ : Sp12to4
    port map (
            O => \N__23460\,
            I => \N__23417\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__23457\,
            I => \N__23417\
        );

    \I__3369\ : InMux
    port map (
            O => \N__23454\,
            I => \N__23414\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__23449\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__23440\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__23437\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3365\ : Odrv4
    port map (
            O => \N__23432\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3364\ : Odrv4
    port map (
            O => \N__23429\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__23426\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3362\ : Odrv12
    port map (
            O => \N__23417\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__23414\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3360\ : InMux
    port map (
            O => \N__23397\,
            I => \N__23394\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__23394\,
            I => \N__23391\
        );

    \I__3358\ : Span4Mux_h
    port map (
            O => \N__23391\,
            I => \N__23388\
        );

    \I__3357\ : Odrv4
    port map (
            O => \N__23388\,
            I => il_max_comp2_c
        );

    \I__3356\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__23382\,
            I => \N__23377\
        );

    \I__3354\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23374\
        );

    \I__3353\ : InMux
    port map (
            O => \N__23380\,
            I => \N__23371\
        );

    \I__3352\ : Span4Mux_v
    port map (
            O => \N__23377\,
            I => \N__23368\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__23374\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__23371\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3349\ : Odrv4
    port map (
            O => \N__23368\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3348\ : InMux
    port map (
            O => \N__23361\,
            I => \N__23358\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__23358\,
            I => \N__23353\
        );

    \I__3346\ : InMux
    port map (
            O => \N__23357\,
            I => \N__23350\
        );

    \I__3345\ : InMux
    port map (
            O => \N__23356\,
            I => \N__23347\
        );

    \I__3344\ : Span4Mux_v
    port map (
            O => \N__23353\,
            I => \N__23344\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__23350\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__23347\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3341\ : Odrv4
    port map (
            O => \N__23344\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23337\,
            I => \N__23333\
        );

    \I__3339\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23329\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__23333\,
            I => \N__23326\
        );

    \I__3337\ : InMux
    port map (
            O => \N__23332\,
            I => \N__23323\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__23329\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__23326\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__23323\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3333\ : InMux
    port map (
            O => \N__23316\,
            I => \N__23311\
        );

    \I__3332\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23308\
        );

    \I__3331\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23305\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__23311\,
            I => \N__23302\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__23308\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__23305\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__23302\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3326\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23290\
        );

    \I__3325\ : InMux
    port map (
            O => \N__23294\,
            I => \N__23287\
        );

    \I__3324\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23284\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__23290\,
            I => \N__23281\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__23287\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__23284\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__23281\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3319\ : InMux
    port map (
            O => \N__23274\,
            I => \N__23270\
        );

    \I__3318\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23266\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__23270\,
            I => \N__23263\
        );

    \I__3316\ : InMux
    port map (
            O => \N__23269\,
            I => \N__23260\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__23266\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3314\ : Odrv12
    port map (
            O => \N__23263\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__23260\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3312\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23249\
        );

    \I__3311\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23246\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__23249\,
            I => \N__23240\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__23246\,
            I => \N__23240\
        );

    \I__3308\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23237\
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__23240\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__23237\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__23232\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__3304\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23225\
        );

    \I__3303\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23222\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__23225\,
            I => \N__23216\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__23222\,
            I => \N__23216\
        );

    \I__3300\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23213\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__23216\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__23213\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3297\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23205\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__23205\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__3295\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23198\
        );

    \I__3294\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23194\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__23198\,
            I => \N__23191\
        );

    \I__3292\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23188\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__23194\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3290\ : Odrv12
    port map (
            O => \N__23191\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__23188\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__23181\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__3287\ : InMux
    port map (
            O => \N__23178\,
            I => \N__23175\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__23175\,
            I => \N__23170\
        );

    \I__3285\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23167\
        );

    \I__3284\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23164\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__23170\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__23167\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__23164\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3280\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23145\
        );

    \I__3279\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23142\
        );

    \I__3278\ : InMux
    port map (
            O => \N__23155\,
            I => \N__23133\
        );

    \I__3277\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23133\
        );

    \I__3276\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23133\
        );

    \I__3275\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23133\
        );

    \I__3274\ : InMux
    port map (
            O => \N__23151\,
            I => \N__23124\
        );

    \I__3273\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23124\
        );

    \I__3272\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23124\
        );

    \I__3271\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23124\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__23145\,
            I => \N__23119\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__23142\,
            I => \N__23119\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__23133\,
            I => \N__23116\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__23124\,
            I => \N__23113\
        );

    \I__3266\ : Span4Mux_h
    port map (
            O => \N__23119\,
            I => \N__23110\
        );

    \I__3265\ : Odrv12
    port map (
            O => \N__23116\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__23113\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__3263\ : Odrv4
    port map (
            O => \N__23110\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__3262\ : InMux
    port map (
            O => \N__23103\,
            I => \N__23100\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__23100\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__3260\ : InMux
    port map (
            O => \N__23097\,
            I => \N__23092\
        );

    \I__3259\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23089\
        );

    \I__3258\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23085\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__23092\,
            I => \N__23082\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__23089\,
            I => \N__23079\
        );

    \I__3255\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23076\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__23085\,
            I => \N__23073\
        );

    \I__3253\ : Span4Mux_h
    port map (
            O => \N__23082\,
            I => \N__23068\
        );

    \I__3252\ : Span4Mux_h
    port map (
            O => \N__23079\,
            I => \N__23068\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__23076\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3250\ : Odrv12
    port map (
            O => \N__23073\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3249\ : Odrv4
    port map (
            O => \N__23068\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3248\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23058\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__23058\,
            I => \N__23055\
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__23055\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23052\,
            I => \N__23045\
        );

    \I__3244\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23045\
        );

    \I__3243\ : InMux
    port map (
            O => \N__23050\,
            I => \N__23042\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__23045\,
            I => \N__23038\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__23042\,
            I => \N__23035\
        );

    \I__3240\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23032\
        );

    \I__3239\ : Span4Mux_h
    port map (
            O => \N__23038\,
            I => \N__23029\
        );

    \I__3238\ : Odrv4
    port map (
            O => \N__23035\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__23032\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__23029\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3235\ : InMux
    port map (
            O => \N__23022\,
            I => \N__23019\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__23019\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__3233\ : InMux
    port map (
            O => \N__23016\,
            I => \N__23013\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__23013\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__3231\ : InMux
    port map (
            O => \N__23010\,
            I => \N__23007\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__23007\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__23004\,
            I => \N__23000\
        );

    \I__3228\ : InMux
    port map (
            O => \N__23003\,
            I => \N__22997\
        );

    \I__3227\ : InMux
    port map (
            O => \N__23000\,
            I => \N__22993\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__22997\,
            I => \N__22989\
        );

    \I__3225\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22986\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__22993\,
            I => \N__22983\
        );

    \I__3223\ : InMux
    port map (
            O => \N__22992\,
            I => \N__22980\
        );

    \I__3222\ : Sp12to4
    port map (
            O => \N__22989\,
            I => \N__22975\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__22986\,
            I => \N__22975\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__22983\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__22980\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3218\ : Odrv12
    port map (
            O => \N__22975\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__22968\,
            I => \N__22965\
        );

    \I__3216\ : InMux
    port map (
            O => \N__22965\,
            I => \N__22962\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__22962\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__22959\,
            I => \N__22953\
        );

    \I__3213\ : InMux
    port map (
            O => \N__22958\,
            I => \N__22950\
        );

    \I__3212\ : CascadeMux
    port map (
            O => \N__22957\,
            I => \N__22947\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__22956\,
            I => \N__22944\
        );

    \I__3210\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22941\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22938\
        );

    \I__3208\ : InMux
    port map (
            O => \N__22947\,
            I => \N__22935\
        );

    \I__3207\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22932\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__22941\,
            I => \N__22929\
        );

    \I__3205\ : Span4Mux_h
    port map (
            O => \N__22938\,
            I => \N__22926\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__22935\,
            I => \N__22923\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__22932\,
            I => \N__22918\
        );

    \I__3202\ : Sp12to4
    port map (
            O => \N__22929\,
            I => \N__22918\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__22926\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__22923\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3199\ : Odrv12
    port map (
            O => \N__22918\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3198\ : InMux
    port map (
            O => \N__22911\,
            I => \N__22908\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__22908\,
            I => \N__22905\
        );

    \I__3196\ : Span4Mux_v
    port map (
            O => \N__22905\,
            I => \N__22902\
        );

    \I__3195\ : Odrv4
    port map (
            O => \N__22902\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__3194\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22896\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__22896\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__22893\,
            I => \N__22890\
        );

    \I__3191\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22887\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__22887\,
            I => \N__22881\
        );

    \I__3189\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22878\
        );

    \I__3188\ : InMux
    port map (
            O => \N__22885\,
            I => \N__22875\
        );

    \I__3187\ : InMux
    port map (
            O => \N__22884\,
            I => \N__22872\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__22881\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__22878\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__22875\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__22872\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__22863\,
            I => \N__22860\
        );

    \I__3181\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22857\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__22857\,
            I => \N__22854\
        );

    \I__3179\ : Span4Mux_v
    port map (
            O => \N__22854\,
            I => \N__22848\
        );

    \I__3178\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22843\
        );

    \I__3177\ : InMux
    port map (
            O => \N__22852\,
            I => \N__22843\
        );

    \I__3176\ : InMux
    port map (
            O => \N__22851\,
            I => \N__22840\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__22848\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__22843\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__22840\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__22833\,
            I => \N__22830\
        );

    \I__3171\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22826\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__22829\,
            I => \N__22823\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__22826\,
            I => \N__22818\
        );

    \I__3168\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22813\
        );

    \I__3167\ : InMux
    port map (
            O => \N__22822\,
            I => \N__22813\
        );

    \I__3166\ : InMux
    port map (
            O => \N__22821\,
            I => \N__22810\
        );

    \I__3165\ : Span4Mux_h
    port map (
            O => \N__22818\,
            I => \N__22805\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__22813\,
            I => \N__22805\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__22810\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__22805\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__3161\ : CascadeMux
    port map (
            O => \N__22800\,
            I => \N__22797\
        );

    \I__3160\ : InMux
    port map (
            O => \N__22797\,
            I => \N__22794\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__22794\,
            I => \N__22791\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__22791\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__3157\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22784\
        );

    \I__3156\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22780\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__22784\,
            I => \N__22777\
        );

    \I__3154\ : InMux
    port map (
            O => \N__22783\,
            I => \N__22774\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22770\
        );

    \I__3152\ : Span4Mux_h
    port map (
            O => \N__22777\,
            I => \N__22765\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__22774\,
            I => \N__22765\
        );

    \I__3150\ : InMux
    port map (
            O => \N__22773\,
            I => \N__22762\
        );

    \I__3149\ : Span4Mux_h
    port map (
            O => \N__22770\,
            I => \N__22755\
        );

    \I__3148\ : Span4Mux_h
    port map (
            O => \N__22765\,
            I => \N__22755\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__22762\,
            I => \N__22755\
        );

    \I__3146\ : Odrv4
    port map (
            O => \N__22755\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3145\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22749\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__22749\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__3143\ : InMux
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__22743\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__22740\,
            I => \N__22737\
        );

    \I__3140\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22732\
        );

    \I__3139\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22729\
        );

    \I__3138\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22726\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__22732\,
            I => \N__22723\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__22729\,
            I => \N__22718\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__22726\,
            I => \N__22718\
        );

    \I__3134\ : Span4Mux_s3_h
    port map (
            O => \N__22723\,
            I => \N__22714\
        );

    \I__3133\ : Span4Mux_h
    port map (
            O => \N__22718\,
            I => \N__22711\
        );

    \I__3132\ : InMux
    port map (
            O => \N__22717\,
            I => \N__22708\
        );

    \I__3131\ : Odrv4
    port map (
            O => \N__22714\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3130\ : Odrv4
    port map (
            O => \N__22711\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__22708\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3128\ : InMux
    port map (
            O => \N__22701\,
            I => \N__22698\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__22698\,
            I => \N__22695\
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__22695\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__22692\,
            I => \N__22689\
        );

    \I__3124\ : InMux
    port map (
            O => \N__22689\,
            I => \N__22685\
        );

    \I__3123\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22682\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__22685\,
            I => \N__22677\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__22682\,
            I => \N__22674\
        );

    \I__3120\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22671\
        );

    \I__3119\ : InMux
    port map (
            O => \N__22680\,
            I => \N__22668\
        );

    \I__3118\ : Span4Mux_h
    port map (
            O => \N__22677\,
            I => \N__22665\
        );

    \I__3117\ : Span4Mux_v
    port map (
            O => \N__22674\,
            I => \N__22658\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__22671\,
            I => \N__22658\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__22668\,
            I => \N__22658\
        );

    \I__3114\ : Odrv4
    port map (
            O => \N__22665\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__22658\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__22653\,
            I => \N__22650\
        );

    \I__3111\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22647\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__22647\,
            I => \N__22644\
        );

    \I__3109\ : Odrv12
    port map (
            O => \N__22644\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__22641\,
            I => \N__22638\
        );

    \I__3107\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22635\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__22635\,
            I => \N__22632\
        );

    \I__3105\ : Odrv12
    port map (
            O => \N__22632\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__3104\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22626\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__22626\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__22623\,
            I => \N__22618\
        );

    \I__3101\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22615\
        );

    \I__3100\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22611\
        );

    \I__3099\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22608\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__22615\,
            I => \N__22605\
        );

    \I__3097\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22602\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__22611\,
            I => \N__22599\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__22608\,
            I => \N__22596\
        );

    \I__3094\ : Span4Mux_v
    port map (
            O => \N__22605\,
            I => \N__22591\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__22602\,
            I => \N__22591\
        );

    \I__3092\ : Odrv4
    port map (
            O => \N__22599\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__22596\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3090\ : Odrv4
    port map (
            O => \N__22591\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3089\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22581\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__22581\,
            I => \N__22578\
        );

    \I__3087\ : Span4Mux_v
    port map (
            O => \N__22578\,
            I => \N__22575\
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__22575\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__22572\,
            I => \N__22567\
        );

    \I__3084\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22564\
        );

    \I__3083\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22561\
        );

    \I__3082\ : InMux
    port map (
            O => \N__22567\,
            I => \N__22558\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__22564\,
            I => \N__22554\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__22561\,
            I => \N__22551\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__22558\,
            I => \N__22548\
        );

    \I__3078\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22545\
        );

    \I__3077\ : Span4Mux_v
    port map (
            O => \N__22554\,
            I => \N__22542\
        );

    \I__3076\ : Span4Mux_h
    port map (
            O => \N__22551\,
            I => \N__22539\
        );

    \I__3075\ : Span4Mux_v
    port map (
            O => \N__22548\,
            I => \N__22534\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__22545\,
            I => \N__22534\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__22542\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__22539\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3071\ : Odrv4
    port map (
            O => \N__22534\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3070\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22524\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__22524\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__3068\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22517\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__22520\,
            I => \N__22513\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__22517\,
            I => \N__22510\
        );

    \I__3065\ : InMux
    port map (
            O => \N__22516\,
            I => \N__22506\
        );

    \I__3064\ : InMux
    port map (
            O => \N__22513\,
            I => \N__22503\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__22510\,
            I => \N__22500\
        );

    \I__3062\ : InMux
    port map (
            O => \N__22509\,
            I => \N__22497\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__22506\,
            I => \N__22492\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__22503\,
            I => \N__22492\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__22500\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__22497\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__22492\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3056\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22482\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__22482\,
            I => \N__22477\
        );

    \I__3054\ : InMux
    port map (
            O => \N__22481\,
            I => \N__22474\
        );

    \I__3053\ : InMux
    port map (
            O => \N__22480\,
            I => \N__22470\
        );

    \I__3052\ : Span4Mux_v
    port map (
            O => \N__22477\,
            I => \N__22467\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__22474\,
            I => \N__22464\
        );

    \I__3050\ : InMux
    port map (
            O => \N__22473\,
            I => \N__22461\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__22470\,
            I => \N__22458\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__22467\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__22464\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__22461\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__22458\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__22449\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\
        );

    \I__3043\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22442\
        );

    \I__3042\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22439\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__22442\,
            I => \N__22432\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__22439\,
            I => \N__22432\
        );

    \I__3039\ : InMux
    port map (
            O => \N__22438\,
            I => \N__22429\
        );

    \I__3038\ : InMux
    port map (
            O => \N__22437\,
            I => \N__22426\
        );

    \I__3037\ : Span4Mux_h
    port map (
            O => \N__22432\,
            I => \N__22423\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__22429\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__22426\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__22423\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3033\ : InMux
    port map (
            O => \N__22416\,
            I => \N__22412\
        );

    \I__3032\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22409\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__22412\,
            I => \N__22404\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__22409\,
            I => \N__22401\
        );

    \I__3029\ : InMux
    port map (
            O => \N__22408\,
            I => \N__22398\
        );

    \I__3028\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22395\
        );

    \I__3027\ : Span4Mux_v
    port map (
            O => \N__22404\,
            I => \N__22392\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__22401\,
            I => \N__22385\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__22398\,
            I => \N__22385\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__22395\,
            I => \N__22385\
        );

    \I__3023\ : Span4Mux_v
    port map (
            O => \N__22392\,
            I => \N__22382\
        );

    \I__3022\ : Span4Mux_v
    port map (
            O => \N__22385\,
            I => \N__22379\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__22382\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__22379\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__22374\,
            I => \N__22371\
        );

    \I__3018\ : InMux
    port map (
            O => \N__22371\,
            I => \N__22367\
        );

    \I__3017\ : InMux
    port map (
            O => \N__22370\,
            I => \N__22363\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__22367\,
            I => \N__22360\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__22366\,
            I => \N__22357\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__22363\,
            I => \N__22353\
        );

    \I__3013\ : Span12Mux_s5_h
    port map (
            O => \N__22360\,
            I => \N__22350\
        );

    \I__3012\ : InMux
    port map (
            O => \N__22357\,
            I => \N__22347\
        );

    \I__3011\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22344\
        );

    \I__3010\ : Span4Mux_v
    port map (
            O => \N__22353\,
            I => \N__22341\
        );

    \I__3009\ : Odrv12
    port map (
            O => \N__22350\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__22347\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__22344\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3006\ : Odrv4
    port map (
            O => \N__22341\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__22332\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\
        );

    \I__3004\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22326\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__22326\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\
        );

    \I__3002\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22320\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__22320\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\
        );

    \I__3000\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22314\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__22314\,
            I => \N__22311\
        );

    \I__2998\ : Odrv4
    port map (
            O => \N__22311\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__2997\ : InMux
    port map (
            O => \N__22308\,
            I => \N__22305\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__22305\,
            I => \N__22302\
        );

    \I__2995\ : Odrv4
    port map (
            O => \N__22302\,
            I => \current_shift_inst.PI_CTRL.N_167\
        );

    \I__2994\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22296\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__22296\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__2992\ : InMux
    port map (
            O => \N__22293\,
            I => \N__22290\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__22290\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__22287\,
            I => \current_shift_inst.PI_CTRL.N_171_cascade_\
        );

    \I__2989\ : InMux
    port map (
            O => \N__22284\,
            I => \N__22281\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__22281\,
            I => \N__22275\
        );

    \I__2987\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22270\
        );

    \I__2986\ : InMux
    port map (
            O => \N__22279\,
            I => \N__22270\
        );

    \I__2985\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22267\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__22275\,
            I => \N__22262\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22262\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__22267\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__22262\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__22257\,
            I => \N__22254\
        );

    \I__2979\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22251\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__22251\,
            I => \N__22248\
        );

    \I__2977\ : Span4Mux_h
    port map (
            O => \N__22248\,
            I => \N__22245\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__22245\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__22242\,
            I => \N__22239\
        );

    \I__2974\ : InMux
    port map (
            O => \N__22239\,
            I => \N__22235\
        );

    \I__2973\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22232\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__22235\,
            I => \N__22227\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__22232\,
            I => \N__22224\
        );

    \I__2970\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22221\
        );

    \I__2969\ : InMux
    port map (
            O => \N__22230\,
            I => \N__22218\
        );

    \I__2968\ : Span4Mux_v
    port map (
            O => \N__22227\,
            I => \N__22215\
        );

    \I__2967\ : Span4Mux_v
    port map (
            O => \N__22224\,
            I => \N__22208\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__22221\,
            I => \N__22208\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__22218\,
            I => \N__22208\
        );

    \I__2964\ : Odrv4
    port map (
            O => \N__22215\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2963\ : Odrv4
    port map (
            O => \N__22208\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2962\ : InMux
    port map (
            O => \N__22203\,
            I => \N__22200\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__22200\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__22197\,
            I => \N__22193\
        );

    \I__2959\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22189\
        );

    \I__2958\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22185\
        );

    \I__2957\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22182\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__22189\,
            I => \N__22179\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__22188\,
            I => \N__22176\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__22185\,
            I => \N__22173\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__22182\,
            I => \N__22168\
        );

    \I__2952\ : Span4Mux_h
    port map (
            O => \N__22179\,
            I => \N__22168\
        );

    \I__2951\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22165\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__22173\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__22168\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__22165\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2947\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22155\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__22155\,
            I => \N__22152\
        );

    \I__2945\ : Span4Mux_h
    port map (
            O => \N__22152\,
            I => \N__22149\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__22149\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__22146\,
            I => \N__22142\
        );

    \I__2942\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22139\
        );

    \I__2941\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22135\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__22139\,
            I => \N__22131\
        );

    \I__2939\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22128\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__22135\,
            I => \N__22125\
        );

    \I__2937\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22122\
        );

    \I__2936\ : Span4Mux_h
    port map (
            O => \N__22131\,
            I => \N__22119\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__22128\,
            I => \N__22116\
        );

    \I__2934\ : Span4Mux_v
    port map (
            O => \N__22125\,
            I => \N__22111\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__22122\,
            I => \N__22111\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__22119\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2931\ : Odrv4
    port map (
            O => \N__22116\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2930\ : Odrv4
    port map (
            O => \N__22111\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2929\ : InMux
    port map (
            O => \N__22104\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__2928\ : InMux
    port map (
            O => \N__22101\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__2927\ : InMux
    port map (
            O => \N__22098\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__2926\ : InMux
    port map (
            O => \N__22095\,
            I => \bfn_5_7_0_\
        );

    \I__2925\ : InMux
    port map (
            O => \N__22092\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__2924\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22086\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__22086\,
            I => \N__22083\
        );

    \I__2922\ : Span4Mux_v
    port map (
            O => \N__22083\,
            I => \N__22080\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__22080\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__22077\,
            I => \N__22074\
        );

    \I__2919\ : InMux
    port map (
            O => \N__22074\,
            I => \N__22071\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__22071\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__2917\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22065\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__22065\,
            I => \N__22060\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22057\
        );

    \I__2914\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22053\
        );

    \I__2913\ : Span12Mux_s4_h
    port map (
            O => \N__22060\,
            I => \N__22048\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__22057\,
            I => \N__22048\
        );

    \I__2911\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22045\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__22053\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2909\ : Odrv12
    port map (
            O => \N__22048\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__22045\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__22038\,
            I => \N__22034\
        );

    \I__2906\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22030\
        );

    \I__2905\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22027\
        );

    \I__2904\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22024\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__22030\,
            I => \counterZ0Z_1\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__22027\,
            I => \counterZ0Z_1\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__22024\,
            I => \counterZ0Z_1\
        );

    \I__2900\ : InMux
    port map (
            O => \N__22017\,
            I => \N__22009\
        );

    \I__2899\ : InMux
    port map (
            O => \N__22016\,
            I => \N__22009\
        );

    \I__2898\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22006\
        );

    \I__2897\ : InMux
    port map (
            O => \N__22014\,
            I => \N__22003\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__22009\,
            I => \counterZ0Z_0\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__22006\,
            I => \counterZ0Z_0\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__22003\,
            I => \counterZ0Z_0\
        );

    \I__2893\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21989\
        );

    \I__2892\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21989\
        );

    \I__2891\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21981\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__21989\,
            I => \N__21978\
        );

    \I__2889\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21973\
        );

    \I__2888\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21973\
        );

    \I__2887\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21970\
        );

    \I__2886\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21965\
        );

    \I__2885\ : InMux
    port map (
            O => \N__21984\,
            I => \N__21965\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__21981\,
            I => \current_shift_inst.PI_CTRL.un2_counterZ0\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__21978\,
            I => \current_shift_inst.PI_CTRL.un2_counterZ0\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__21973\,
            I => \current_shift_inst.PI_CTRL.un2_counterZ0\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__21970\,
            I => \current_shift_inst.PI_CTRL.un2_counterZ0\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__21965\,
            I => \current_shift_inst.PI_CTRL.un2_counterZ0\
        );

    \I__2879\ : InMux
    port map (
            O => \N__21954\,
            I => \N__21950\
        );

    \I__2878\ : InMux
    port map (
            O => \N__21953\,
            I => \N__21947\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__21950\,
            I => clk_10khz_i
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__21947\,
            I => clk_10khz_i
        );

    \I__2875\ : InMux
    port map (
            O => \N__21942\,
            I => \bfn_5_6_0_\
        );

    \I__2874\ : InMux
    port map (
            O => \N__21939\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__2873\ : InMux
    port map (
            O => \N__21936\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__2872\ : InMux
    port map (
            O => \N__21933\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__2871\ : InMux
    port map (
            O => \N__21930\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__2870\ : InMux
    port map (
            O => \N__21927\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__2869\ : InMux
    port map (
            O => \N__21924\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__2868\ : InMux
    port map (
            O => \N__21921\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__2867\ : InMux
    port map (
            O => \N__21918\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__2866\ : InMux
    port map (
            O => \N__21915\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__2865\ : InMux
    port map (
            O => \N__21912\,
            I => \N__21908\
        );

    \I__2864\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21905\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__21908\,
            I => \N__21902\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__21905\,
            I => \counterZ0Z_11\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__21902\,
            I => \counterZ0Z_11\
        );

    \I__2860\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21893\
        );

    \I__2859\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21890\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__21893\,
            I => \counterZ0Z_6\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__21890\,
            I => \counterZ0Z_6\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__21885\,
            I => \N__21881\
        );

    \I__2855\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21878\
        );

    \I__2854\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21875\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__21878\,
            I => \counterZ0Z_12\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__21875\,
            I => \counterZ0Z_12\
        );

    \I__2851\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21866\
        );

    \I__2850\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21863\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__21866\,
            I => \counterZ0Z_10\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__21863\,
            I => \counterZ0Z_10\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__21858\,
            I => \current_shift_inst.PI_CTRL.un2_counterZ0Z_1_cascade_\
        );

    \I__2846\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21851\
        );

    \I__2845\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21848\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__21851\,
            I => \counterZ0Z_8\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__21848\,
            I => \counterZ0Z_8\
        );

    \I__2842\ : InMux
    port map (
            O => \N__21843\,
            I => \N__21839\
        );

    \I__2841\ : InMux
    port map (
            O => \N__21842\,
            I => \N__21836\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__21839\,
            I => \counterZ0Z_7\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__21836\,
            I => \counterZ0Z_7\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__21831\,
            I => \N__21828\
        );

    \I__2837\ : InMux
    port map (
            O => \N__21828\,
            I => \N__21824\
        );

    \I__2836\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21821\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__21824\,
            I => \N__21818\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__21821\,
            I => \counterZ0Z_9\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__21818\,
            I => \counterZ0Z_9\
        );

    \I__2832\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21809\
        );

    \I__2831\ : InMux
    port map (
            O => \N__21812\,
            I => \N__21806\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__21809\,
            I => \counterZ0Z_5\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__21806\,
            I => \counterZ0Z_5\
        );

    \I__2828\ : InMux
    port map (
            O => \N__21801\,
            I => \N__21798\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__21798\,
            I => \current_shift_inst.PI_CTRL.un2_counterZ0Z_8\
        );

    \I__2826\ : InMux
    port map (
            O => \N__21795\,
            I => \N__21791\
        );

    \I__2825\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21788\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__21791\,
            I => \counterZ0Z_2\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__21788\,
            I => \counterZ0Z_2\
        );

    \I__2822\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21779\
        );

    \I__2821\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21776\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__21779\,
            I => \counterZ0Z_3\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__21776\,
            I => \counterZ0Z_3\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__21771\,
            I => \N__21767\
        );

    \I__2817\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21764\
        );

    \I__2816\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21761\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__21764\,
            I => \counterZ0Z_4\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__21761\,
            I => \counterZ0Z_4\
        );

    \I__2813\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21753\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__21753\,
            I => \current_shift_inst.PI_CTRL.un2_counterZ0Z_7\
        );

    \I__2811\ : InMux
    port map (
            O => \N__21750\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__2810\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21744\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__21744\,
            I => \N__21741\
        );

    \I__2808\ : Odrv4
    port map (
            O => \N__21741\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__2807\ : InMux
    port map (
            O => \N__21738\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__2806\ : InMux
    port map (
            O => \N__21735\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__2805\ : InMux
    port map (
            O => \N__21732\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__2804\ : InMux
    port map (
            O => \N__21729\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__2803\ : InMux
    port map (
            O => \N__21726\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__2802\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21720\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__21720\,
            I => \N__21717\
        );

    \I__2800\ : Span4Mux_v
    port map (
            O => \N__21717\,
            I => \N__21714\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__21714\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__2798\ : InMux
    port map (
            O => \N__21711\,
            I => \bfn_4_16_0_\
        );

    \I__2797\ : InMux
    port map (
            O => \N__21708\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\
        );

    \I__2796\ : InMux
    port map (
            O => \N__21705\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__2795\ : InMux
    port map (
            O => \N__21702\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__2794\ : InMux
    port map (
            O => \N__21699\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__2793\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21693\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__21693\,
            I => \N__21690\
        );

    \I__2791\ : Odrv4
    port map (
            O => \N__21690\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__2790\ : InMux
    port map (
            O => \N__21687\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__2789\ : InMux
    port map (
            O => \N__21684\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__2788\ : InMux
    port map (
            O => \N__21681\,
            I => \N__21675\
        );

    \I__2787\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21675\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__21675\,
            I => \N__21671\
        );

    \I__2785\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21667\
        );

    \I__2784\ : Span4Mux_h
    port map (
            O => \N__21671\,
            I => \N__21664\
        );

    \I__2783\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21661\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__21667\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__21664\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__21661\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2779\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21651\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__21651\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__2777\ : InMux
    port map (
            O => \N__21648\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__2776\ : InMux
    port map (
            O => \N__21645\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__2775\ : InMux
    port map (
            O => \N__21642\,
            I => \bfn_4_15_0_\
        );

    \I__2774\ : InMux
    port map (
            O => \N__21639\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\
        );

    \I__2773\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21633\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__21633\,
            I => \N__21630\
        );

    \I__2771\ : Odrv12
    port map (
            O => \N__21630\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__2770\ : InMux
    port map (
            O => \N__21627\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\
        );

    \I__2769\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__21621\,
            I => \N__21618\
        );

    \I__2767\ : Span4Mux_h
    port map (
            O => \N__21618\,
            I => \N__21613\
        );

    \I__2766\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21610\
        );

    \I__2765\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21607\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__21613\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__21610\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__21607\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2761\ : InMux
    port map (
            O => \N__21600\,
            I => \N__21597\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__21597\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__2759\ : InMux
    port map (
            O => \N__21594\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__2758\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21586\
        );

    \I__2757\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21580\
        );

    \I__2756\ : InMux
    port map (
            O => \N__21589\,
            I => \N__21580\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__21586\,
            I => \N__21577\
        );

    \I__2754\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21574\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__21580\,
            I => \N__21569\
        );

    \I__2752\ : Span4Mux_h
    port map (
            O => \N__21577\,
            I => \N__21569\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__21574\,
            I => \N__21566\
        );

    \I__2750\ : Odrv4
    port map (
            O => \N__21569\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2749\ : Odrv12
    port map (
            O => \N__21566\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2748\ : InMux
    port map (
            O => \N__21561\,
            I => \N__21558\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__21558\,
            I => \N__21555\
        );

    \I__2746\ : Odrv12
    port map (
            O => \N__21555\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__2745\ : InMux
    port map (
            O => \N__21552\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__2744\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21546\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__21546\,
            I => \N__21543\
        );

    \I__2742\ : Span4Mux_h
    port map (
            O => \N__21543\,
            I => \N__21537\
        );

    \I__2741\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21534\
        );

    \I__2740\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21529\
        );

    \I__2739\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21529\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__21537\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__21534\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__21529\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2735\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21519\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__21519\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__2733\ : InMux
    port map (
            O => \N__21516\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__2732\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21510\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__21510\,
            I => \N__21507\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__21507\,
            I => \N__21501\
        );

    \I__2729\ : InMux
    port map (
            O => \N__21506\,
            I => \N__21498\
        );

    \I__2728\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21493\
        );

    \I__2727\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21493\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__21501\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__21498\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__21493\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2723\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21483\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__21483\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__2721\ : InMux
    port map (
            O => \N__21480\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__2720\ : InMux
    port map (
            O => \N__21477\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__2719\ : InMux
    port map (
            O => \N__21474\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__2718\ : InMux
    port map (
            O => \N__21471\,
            I => \bfn_4_14_0_\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__21468\,
            I => \N__21464\
        );

    \I__2716\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21457\
        );

    \I__2715\ : InMux
    port map (
            O => \N__21464\,
            I => \N__21457\
        );

    \I__2714\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21454\
        );

    \I__2713\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21451\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__21457\,
            I => \N__21448\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__21454\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__21451\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__21448\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2708\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21438\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__21438\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__2706\ : InMux
    port map (
            O => \N__21435\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\
        );

    \I__2705\ : InMux
    port map (
            O => \N__21432\,
            I => \N__21429\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__21429\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\
        );

    \I__2703\ : InMux
    port map (
            O => \N__21426\,
            I => \N__21423\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__21423\,
            I => \N__21418\
        );

    \I__2701\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21414\
        );

    \I__2700\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21411\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__21418\,
            I => \N__21408\
        );

    \I__2698\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21405\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__21414\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__21411\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__21408\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__21405\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__21396\,
            I => \N__21393\
        );

    \I__2692\ : InMux
    port map (
            O => \N__21393\,
            I => \N__21390\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__21390\,
            I => \N__21387\
        );

    \I__2690\ : Odrv4
    port map (
            O => \N__21387\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__2689\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21381\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__21381\,
            I => \N__21378\
        );

    \I__2687\ : Span4Mux_v
    port map (
            O => \N__21378\,
            I => \N__21373\
        );

    \I__2686\ : InMux
    port map (
            O => \N__21377\,
            I => \N__21370\
        );

    \I__2685\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21367\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__21373\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__21370\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__21367\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2681\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21357\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__21357\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\
        );

    \I__2679\ : InMux
    port map (
            O => \N__21354\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2678\ : IoInMux
    port map (
            O => \N__21351\,
            I => \N__21348\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__21348\,
            I => \N__21345\
        );

    \I__2676\ : Span12Mux_s6_v
    port map (
            O => \N__21345\,
            I => \N__21342\
        );

    \I__2675\ : Span12Mux_h
    port map (
            O => \N__21342\,
            I => \N__21339\
        );

    \I__2674\ : Odrv12
    port map (
            O => \N__21339\,
            I => pwm_output_c
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__21336\,
            I => \current_shift_inst.PI_CTRL.N_170_cascade_\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__21333\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\
        );

    \I__2671\ : InMux
    port map (
            O => \N__21330\,
            I => \N__21327\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__21327\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\
        );

    \I__2669\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21321\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__21321\,
            I => \current_shift_inst.PI_CTRL.N_168\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__21318\,
            I => \N__21315\
        );

    \I__2666\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21312\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__21312\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\
        );

    \I__2664\ : InMux
    port map (
            O => \N__21309\,
            I => \N__21306\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__21306\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__21303\,
            I => \N__21300\
        );

    \I__2661\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21297\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N__21294\
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__21294\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__2658\ : InMux
    port map (
            O => \N__21291\,
            I => \N__21288\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__21288\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__21285\,
            I => \N__21282\
        );

    \I__2655\ : InMux
    port map (
            O => \N__21282\,
            I => \N__21279\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__21279\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__2653\ : InMux
    port map (
            O => \N__21276\,
            I => \N__21273\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__21273\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__21270\,
            I => \N__21267\
        );

    \I__2650\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21264\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__21264\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__2648\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21258\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__21258\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2646\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21252\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__21252\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__21249\,
            I => \N__21246\
        );

    \I__2643\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21243\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__21243\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__21240\,
            I => \N__21237\
        );

    \I__2640\ : InMux
    port map (
            O => \N__21237\,
            I => \N__21234\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__21234\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__2638\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21228\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__21228\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__21225\,
            I => \N__21222\
        );

    \I__2635\ : InMux
    port map (
            O => \N__21222\,
            I => \N__21219\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__21219\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__2633\ : InMux
    port map (
            O => \N__21216\,
            I => \N__21213\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__21213\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__21210\,
            I => \N__21207\
        );

    \I__2630\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21204\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__21204\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__2628\ : InMux
    port map (
            O => \N__21201\,
            I => \N__21198\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__21198\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__21195\,
            I => \N__21192\
        );

    \I__2625\ : InMux
    port map (
            O => \N__21192\,
            I => \N__21189\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__21189\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__2623\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21183\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__21183\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2621\ : InMux
    port map (
            O => \N__21180\,
            I => un5_counter_cry_6
        );

    \I__2620\ : InMux
    port map (
            O => \N__21177\,
            I => un5_counter_cry_7
        );

    \I__2619\ : InMux
    port map (
            O => \N__21174\,
            I => \bfn_3_19_0_\
        );

    \I__2618\ : InMux
    port map (
            O => \N__21171\,
            I => un5_counter_cry_9
        );

    \I__2617\ : InMux
    port map (
            O => \N__21168\,
            I => un5_counter_cry_10
        );

    \I__2616\ : InMux
    port map (
            O => \N__21165\,
            I => un5_counter_cry_11
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__21162\,
            I => \N__21159\
        );

    \I__2614\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__21156\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__2612\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21150\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__21150\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__2609\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21141\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__21141\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__2607\ : InMux
    port map (
            O => \N__21138\,
            I => \N__21135\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__21135\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__21132\,
            I => \N__21126\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__21131\,
            I => \N__21122\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__21130\,
            I => \N__21118\
        );

    \I__2602\ : InMux
    port map (
            O => \N__21129\,
            I => \N__21102\
        );

    \I__2601\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21102\
        );

    \I__2600\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21102\
        );

    \I__2599\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21102\
        );

    \I__2598\ : InMux
    port map (
            O => \N__21121\,
            I => \N__21102\
        );

    \I__2597\ : InMux
    port map (
            O => \N__21118\,
            I => \N__21102\
        );

    \I__2596\ : InMux
    port map (
            O => \N__21117\,
            I => \N__21102\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__21102\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__2594\ : InMux
    port map (
            O => \N__21099\,
            I => \N__21096\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__21096\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__21093\,
            I => \N__21090\
        );

    \I__2591\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21087\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__21087\,
            I => \N__21084\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__21084\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__2588\ : InMux
    port map (
            O => \N__21081\,
            I => un5_counter_cry_1
        );

    \I__2587\ : InMux
    port map (
            O => \N__21078\,
            I => un5_counter_cry_2
        );

    \I__2586\ : InMux
    port map (
            O => \N__21075\,
            I => un5_counter_cry_3
        );

    \I__2585\ : InMux
    port map (
            O => \N__21072\,
            I => un5_counter_cry_4
        );

    \I__2584\ : InMux
    port map (
            O => \N__21069\,
            I => un5_counter_cry_5
        );

    \I__2583\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21063\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__21063\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__2581\ : InMux
    port map (
            O => \N__21060\,
            I => \N__21057\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__21057\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__21054\,
            I => \N__21051\
        );

    \I__2578\ : InMux
    port map (
            O => \N__21051\,
            I => \N__21048\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__21048\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__21045\,
            I => \N__21042\
        );

    \I__2575\ : InMux
    port map (
            O => \N__21042\,
            I => \N__21039\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__21039\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__21036\,
            I => \N__21033\
        );

    \I__2572\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21030\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__21030\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__21027\,
            I => \N__21024\
        );

    \I__2569\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21021\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__21021\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__21018\,
            I => \N__21015\
        );

    \I__2566\ : InMux
    port map (
            O => \N__21015\,
            I => \N__21012\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__21012\,
            I => \N__21009\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__21009\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__2563\ : InMux
    port map (
            O => \N__21006\,
            I => \N__21003\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__21003\,
            I => \N__21000\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__21000\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__20997\,
            I => \N__20994\
        );

    \I__2559\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20991\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__20991\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__20988\,
            I => \N__20985\
        );

    \I__2556\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20982\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__20982\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2554\ : InMux
    port map (
            O => \N__20979\,
            I => \N__20976\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__20976\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__20973\,
            I => \N__20970\
        );

    \I__2551\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20967\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__20967\,
            I => \N__20964\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__20964\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__20961\,
            I => \N__20958\
        );

    \I__2547\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20955\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__20955\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__2545\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20949\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__20949\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__20946\,
            I => \N__20943\
        );

    \I__2542\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20940\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__20940\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__20937\,
            I => \N__20934\
        );

    \I__2539\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20931\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__20931\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__20928\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__20925\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__20922\,
            I => \N__20919\
        );

    \I__2534\ : InMux
    port map (
            O => \N__20919\,
            I => \N__20916\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__20916\,
            I => \current_shift_inst.PI_CTRL.un1_enablelt3_0\
        );

    \I__2532\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20910\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__20910\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__2529\ : InMux
    port map (
            O => \N__20904\,
            I => \N__20901\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__20901\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__2526\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20892\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__20892\,
            I => \N__20889\
        );

    \I__2524\ : Odrv4
    port map (
            O => \N__20889\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__20886\,
            I => \N__20883\
        );

    \I__2522\ : InMux
    port map (
            O => \N__20883\,
            I => \N__20880\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__20880\,
            I => \N__20877\
        );

    \I__2520\ : Odrv4
    port map (
            O => \N__20877\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2519\ : InMux
    port map (
            O => \N__20874\,
            I => \N__20870\
        );

    \I__2518\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20866\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__20870\,
            I => \N__20863\
        );

    \I__2516\ : InMux
    port map (
            O => \N__20869\,
            I => \N__20860\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__20866\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2514\ : Odrv12
    port map (
            O => \N__20863\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__20860\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__20853\,
            I => \N__20850\
        );

    \I__2511\ : InMux
    port map (
            O => \N__20850\,
            I => \N__20847\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__20847\,
            I => \N__20844\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__20844\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__2508\ : InMux
    port map (
            O => \N__20841\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__20838\,
            I => \N__20833\
        );

    \I__2506\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20830\
        );

    \I__2505\ : InMux
    port map (
            O => \N__20836\,
            I => \N__20827\
        );

    \I__2504\ : InMux
    port map (
            O => \N__20833\,
            I => \N__20824\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__20830\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__20827\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__20824\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2500\ : InMux
    port map (
            O => \N__20817\,
            I => \N__20814\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__20814\,
            I => \N__20811\
        );

    \I__2498\ : Span4Mux_s3_h
    port map (
            O => \N__20811\,
            I => \N__20808\
        );

    \I__2497\ : Odrv4
    port map (
            O => \N__20808\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__2496\ : InMux
    port map (
            O => \N__20805\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__2495\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20797\
        );

    \I__2494\ : InMux
    port map (
            O => \N__20801\,
            I => \N__20794\
        );

    \I__2493\ : InMux
    port map (
            O => \N__20800\,
            I => \N__20791\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__20797\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__20794\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__20791\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__20784\,
            I => \N__20781\
        );

    \I__2488\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20778\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__20778\,
            I => \N__20775\
        );

    \I__2486\ : Odrv4
    port map (
            O => \N__20775\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__2485\ : InMux
    port map (
            O => \N__20772\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__2484\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20765\
        );

    \I__2483\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20762\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__20765\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__20762\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2480\ : InMux
    port map (
            O => \N__20757\,
            I => \N__20754\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__20754\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__2478\ : InMux
    port map (
            O => \N__20751\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__2477\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20743\
        );

    \I__2476\ : InMux
    port map (
            O => \N__20747\,
            I => \N__20740\
        );

    \I__2475\ : InMux
    port map (
            O => \N__20746\,
            I => \N__20737\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__20743\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__20740\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__20737\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2471\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20727\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__20727\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__2469\ : InMux
    port map (
            O => \N__20724\,
            I => \bfn_3_11_0_\
        );

    \I__2468\ : InMux
    port map (
            O => \N__20721\,
            I => \N__20717\
        );

    \I__2467\ : InMux
    port map (
            O => \N__20720\,
            I => \N__20714\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__20717\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__20714\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2464\ : InMux
    port map (
            O => \N__20709\,
            I => \N__20706\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__20706\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__2462\ : InMux
    port map (
            O => \N__20703\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__2461\ : InMux
    port map (
            O => \N__20700\,
            I => \N__20696\
        );

    \I__2460\ : InMux
    port map (
            O => \N__20699\,
            I => \N__20693\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__20696\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__20693\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2457\ : InMux
    port map (
            O => \N__20688\,
            I => \N__20685\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__20685\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__2455\ : InMux
    port map (
            O => \N__20682\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__2454\ : InMux
    port map (
            O => \N__20679\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__2453\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20673\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__20673\,
            I => \N__20670\
        );

    \I__2451\ : Span4Mux_s3_h
    port map (
            O => \N__20670\,
            I => \N__20667\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__20667\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__2449\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20661\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__20661\,
            I => \N__20658\
        );

    \I__2447\ : Span4Mux_h
    port map (
            O => \N__20658\,
            I => \N__20655\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__20655\,
            I => \pwm_generator_inst.O_5\
        );

    \I__2445\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20649\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__20649\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__2443\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20643\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__20643\,
            I => \N__20640\
        );

    \I__2441\ : Span4Mux_h
    port map (
            O => \N__20640\,
            I => \N__20637\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__20637\,
            I => \pwm_generator_inst.O_6\
        );

    \I__2439\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20631\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__20631\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__2437\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20625\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__20625\,
            I => \N__20622\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__20622\,
            I => \N__20619\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__20619\,
            I => \pwm_generator_inst.O_7\
        );

    \I__2433\ : InMux
    port map (
            O => \N__20616\,
            I => \N__20613\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__20613\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \I__2431\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20607\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__20607\,
            I => \N__20604\
        );

    \I__2429\ : Span4Mux_v
    port map (
            O => \N__20604\,
            I => \N__20601\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__20601\,
            I => \pwm_generator_inst.O_8\
        );

    \I__2427\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20595\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__20595\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__2425\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20589\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__20589\,
            I => \N__20586\
        );

    \I__2423\ : Span4Mux_v
    port map (
            O => \N__20586\,
            I => \N__20583\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__20583\,
            I => \pwm_generator_inst.O_9\
        );

    \I__2421\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__20577\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__2419\ : InMux
    port map (
            O => \N__20574\,
            I => \N__20569\
        );

    \I__2418\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20566\
        );

    \I__2417\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20563\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__20569\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__20566\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__20563\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2413\ : CascadeMux
    port map (
            O => \N__20556\,
            I => \N__20553\
        );

    \I__2412\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20550\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__20550\,
            I => \N__20547\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__20547\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__2409\ : InMux
    port map (
            O => \N__20544\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__20541\,
            I => \N__20537\
        );

    \I__2407\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20530\
        );

    \I__2406\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20527\
        );

    \I__2405\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20522\
        );

    \I__2404\ : InMux
    port map (
            O => \N__20535\,
            I => \N__20522\
        );

    \I__2403\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20519\
        );

    \I__2402\ : InMux
    port map (
            O => \N__20533\,
            I => \N__20510\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__20530\,
            I => \N__20503\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__20527\,
            I => \N__20503\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__20522\,
            I => \N__20503\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__20519\,
            I => \N__20500\
        );

    \I__2397\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20487\
        );

    \I__2396\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20487\
        );

    \I__2395\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20487\
        );

    \I__2394\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20487\
        );

    \I__2393\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20487\
        );

    \I__2392\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20487\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__20510\,
            I => \N__20480\
        );

    \I__2390\ : Span4Mux_v
    port map (
            O => \N__20503\,
            I => \N__20480\
        );

    \I__2389\ : Span4Mux_h
    port map (
            O => \N__20500\,
            I => \N__20480\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__20487\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2387\ : Odrv4
    port map (
            O => \N__20480\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2386\ : InMux
    port map (
            O => \N__20475\,
            I => \N__20472\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__20472\,
            I => \N__20468\
        );

    \I__2384\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20465\
        );

    \I__2383\ : Span4Mux_h
    port map (
            O => \N__20468\,
            I => \N__20460\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__20465\,
            I => \N__20460\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__20460\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__2380\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20454\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__20454\,
            I => \N__20451\
        );

    \I__2378\ : Odrv4
    port map (
            O => \N__20451\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__2377\ : InMux
    port map (
            O => \N__20448\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__2376\ : InMux
    port map (
            O => \N__20445\,
            I => \N__20442\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__20442\,
            I => \N__20439\
        );

    \I__2374\ : Odrv12
    port map (
            O => \N__20439\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__2373\ : InMux
    port map (
            O => \N__20436\,
            I => \N__20433\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__20433\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__2371\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20427\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__20427\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__20424\,
            I => \N__20418\
        );

    \I__2368\ : CascadeMux
    port map (
            O => \N__20423\,
            I => \N__20415\
        );

    \I__2367\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20411\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__20421\,
            I => \N__20403\
        );

    \I__2365\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20398\
        );

    \I__2364\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20398\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__20414\,
            I => \N__20395\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__20411\,
            I => \N__20392\
        );

    \I__2361\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20389\
        );

    \I__2360\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20378\
        );

    \I__2359\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20378\
        );

    \I__2358\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20378\
        );

    \I__2357\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20378\
        );

    \I__2356\ : InMux
    port map (
            O => \N__20403\,
            I => \N__20378\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__20398\,
            I => \N__20375\
        );

    \I__2354\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20372\
        );

    \I__2353\ : Span4Mux_h
    port map (
            O => \N__20392\,
            I => \N__20369\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__20389\,
            I => \N__20366\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__20378\,
            I => \N__20363\
        );

    \I__2350\ : Span4Mux_h
    port map (
            O => \N__20375\,
            I => \N__20358\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__20372\,
            I => \N__20358\
        );

    \I__2348\ : Span4Mux_v
    port map (
            O => \N__20369\,
            I => \N__20355\
        );

    \I__2347\ : Span4Mux_h
    port map (
            O => \N__20366\,
            I => \N__20352\
        );

    \I__2346\ : Span4Mux_v
    port map (
            O => \N__20363\,
            I => \N__20347\
        );

    \I__2345\ : Span4Mux_s2_h
    port map (
            O => \N__20358\,
            I => \N__20347\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__20355\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__20352\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__20347\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__20340\,
            I => \N__20331\
        );

    \I__2340\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20324\
        );

    \I__2339\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20324\
        );

    \I__2338\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20321\
        );

    \I__2337\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20318\
        );

    \I__2336\ : InMux
    port map (
            O => \N__20335\,
            I => \N__20307\
        );

    \I__2335\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20307\
        );

    \I__2334\ : InMux
    port map (
            O => \N__20331\,
            I => \N__20307\
        );

    \I__2333\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20307\
        );

    \I__2332\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20307\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__20324\,
            I => \N__20301\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__20321\,
            I => \N__20301\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__20318\,
            I => \N__20296\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__20307\,
            I => \N__20296\
        );

    \I__2327\ : InMux
    port map (
            O => \N__20306\,
            I => \N__20293\
        );

    \I__2326\ : Span4Mux_v
    port map (
            O => \N__20301\,
            I => \N__20290\
        );

    \I__2325\ : Span4Mux_h
    port map (
            O => \N__20296\,
            I => \N__20285\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__20293\,
            I => \N__20285\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__20290\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__20285\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__20280\,
            I => \N__20271\
        );

    \I__2320\ : InMux
    port map (
            O => \N__20279\,
            I => \N__20264\
        );

    \I__2319\ : InMux
    port map (
            O => \N__20278\,
            I => \N__20264\
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__20277\,
            I => \N__20258\
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__20276\,
            I => \N__20255\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__20275\,
            I => \N__20252\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__20274\,
            I => \N__20247\
        );

    \I__2314\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20244\
        );

    \I__2313\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20239\
        );

    \I__2312\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20239\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__20264\,
            I => \N__20229\
        );

    \I__2310\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20222\
        );

    \I__2309\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20222\
        );

    \I__2308\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20222\
        );

    \I__2307\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20215\
        );

    \I__2306\ : InMux
    port map (
            O => \N__20255\,
            I => \N__20215\
        );

    \I__2305\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20215\
        );

    \I__2304\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20210\
        );

    \I__2303\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20210\
        );

    \I__2302\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20207\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__20244\,
            I => \N__20202\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__20239\,
            I => \N__20202\
        );

    \I__2299\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20176\
        );

    \I__2298\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20176\
        );

    \I__2297\ : InMux
    port map (
            O => \N__20236\,
            I => \N__20176\
        );

    \I__2296\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20176\
        );

    \I__2295\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20176\
        );

    \I__2294\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20176\
        );

    \I__2293\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20176\
        );

    \I__2292\ : Span4Mux_s1_h
    port map (
            O => \N__20229\,
            I => \N__20171\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__20222\,
            I => \N__20171\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__20215\,
            I => \N__20162\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__20210\,
            I => \N__20162\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__20207\,
            I => \N__20162\
        );

    \I__2287\ : Span4Mux_v
    port map (
            O => \N__20202\,
            I => \N__20162\
        );

    \I__2286\ : InMux
    port map (
            O => \N__20201\,
            I => \N__20157\
        );

    \I__2285\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20157\
        );

    \I__2284\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20154\
        );

    \I__2283\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20137\
        );

    \I__2282\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20137\
        );

    \I__2281\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20137\
        );

    \I__2280\ : InMux
    port map (
            O => \N__20195\,
            I => \N__20137\
        );

    \I__2279\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20137\
        );

    \I__2278\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20137\
        );

    \I__2277\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20137\
        );

    \I__2276\ : InMux
    port map (
            O => \N__20191\,
            I => \N__20137\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__20176\,
            I => \N__20132\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__20171\,
            I => \N__20132\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__20162\,
            I => \N_19_1\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__20157\,
            I => \N_19_1\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__20154\,
            I => \N_19_1\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__20137\,
            I => \N_19_1\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__20132\,
            I => \N_19_1\
        );

    \I__2268\ : InMux
    port map (
            O => \N__20121\,
            I => \N__20118\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__20118\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__2266\ : InMux
    port map (
            O => \N__20115\,
            I => \N__20112\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__20112\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__2264\ : InMux
    port map (
            O => \N__20109\,
            I => \N__20106\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__20106\,
            I => \N__20103\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__20103\,
            I => \N__20100\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__20100\,
            I => \pwm_generator_inst.O_0\
        );

    \I__2260\ : InMux
    port map (
            O => \N__20097\,
            I => \N__20094\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__20094\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__2258\ : InMux
    port map (
            O => \N__20091\,
            I => \N__20088\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__20088\,
            I => \N__20085\
        );

    \I__2256\ : Span4Mux_v
    port map (
            O => \N__20085\,
            I => \N__20082\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__20082\,
            I => \pwm_generator_inst.O_1\
        );

    \I__2254\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20076\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__20076\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__2252\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20070\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__20070\,
            I => \N__20067\
        );

    \I__2250\ : Span4Mux_v
    port map (
            O => \N__20067\,
            I => \N__20064\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__20064\,
            I => \pwm_generator_inst.O_2\
        );

    \I__2248\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20058\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__20058\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__2246\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20052\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__20052\,
            I => \N__20049\
        );

    \I__2244\ : Span4Mux_h
    port map (
            O => \N__20049\,
            I => \N__20046\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__20046\,
            I => \pwm_generator_inst.O_3\
        );

    \I__2242\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20040\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__20040\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__2240\ : InMux
    port map (
            O => \N__20037\,
            I => \N__20034\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__20034\,
            I => \N__20031\
        );

    \I__2238\ : Span4Mux_h
    port map (
            O => \N__20031\,
            I => \N__20028\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__20028\,
            I => \pwm_generator_inst.O_4\
        );

    \I__2236\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20022\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__20022\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__2234\ : InMux
    port map (
            O => \N__20019\,
            I => \N__20016\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__20016\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__2232\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20010\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__20010\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__2230\ : InMux
    port map (
            O => \N__20007\,
            I => \N__20004\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__20004\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__2228\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19998\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__19998\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__2226\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19992\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__19992\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__2224\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19986\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__19986\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__2222\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19980\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__19980\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__2220\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19974\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__19974\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__2218\ : InMux
    port map (
            O => \N__19971\,
            I => \N__19967\
        );

    \I__2217\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19964\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__19967\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__19964\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__19959\,
            I => \N__19955\
        );

    \I__2213\ : InMux
    port map (
            O => \N__19958\,
            I => \N__19952\
        );

    \I__2212\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19949\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19946\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__19949\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__19946\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__19941\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\
        );

    \I__2207\ : InMux
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__19935\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2205\ : InMux
    port map (
            O => \N__19932\,
            I => \N__19928\
        );

    \I__2204\ : InMux
    port map (
            O => \N__19931\,
            I => \N__19925\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__19928\,
            I => \N__19920\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__19925\,
            I => \N__19920\
        );

    \I__2201\ : Span4Mux_s3_h
    port map (
            O => \N__19920\,
            I => \N__19917\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__19917\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2199\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19910\
        );

    \I__2198\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19907\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__19910\,
            I => \N__19902\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__19907\,
            I => \N__19902\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__19902\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__19899\,
            I => \N__19896\
        );

    \I__2193\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19893\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__19893\,
            I => \N__19889\
        );

    \I__2191\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19886\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__19889\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__19886\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2188\ : InMux
    port map (
            O => \N__19881\,
            I => \N__19878\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__19878\,
            I => \N__19874\
        );

    \I__2186\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19871\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__19874\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__19871\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2183\ : InMux
    port map (
            O => \N__19866\,
            I => \N__19863\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__19863\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2181\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19857\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19854\
        );

    \I__2179\ : Span12Mux_s11_v
    port map (
            O => \N__19854\,
            I => \N__19851\
        );

    \I__2178\ : Odrv12
    port map (
            O => \N__19851\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2177\ : InMux
    port map (
            O => \N__19848\,
            I => \N__19844\
        );

    \I__2176\ : InMux
    port map (
            O => \N__19847\,
            I => \N__19841\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__19844\,
            I => \N__19838\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__19841\,
            I => \N__19835\
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__19838\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__19835\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__19830\,
            I => \N__19827\
        );

    \I__2170\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19823\
        );

    \I__2169\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19820\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__19823\,
            I => \N__19815\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__19820\,
            I => \N__19815\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__19815\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2165\ : InMux
    port map (
            O => \N__19812\,
            I => \N__19808\
        );

    \I__2164\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19805\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19802\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__19805\,
            I => \N__19799\
        );

    \I__2161\ : Span4Mux_v
    port map (
            O => \N__19802\,
            I => \N__19796\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__19799\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__19796\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2158\ : InMux
    port map (
            O => \N__19791\,
            I => \N__19788\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__19788\,
            I => \N__19785\
        );

    \I__2156\ : Span12Mux_v
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__2155\ : Odrv12
    port map (
            O => \N__19782\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2154\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19775\
        );

    \I__2153\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19772\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__19775\,
            I => \N__19769\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__19772\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__19769\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2149\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19760\
        );

    \I__2148\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19757\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__19760\,
            I => \N__19754\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__19757\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__19754\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2144\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19743\
        );

    \I__2143\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19743\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__19743\,
            I => \N__19740\
        );

    \I__2141\ : Odrv12
    port map (
            O => \N__19740\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2140\ : InMux
    port map (
            O => \N__19737\,
            I => \N__19733\
        );

    \I__2139\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19730\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__19733\,
            I => \N__19725\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19725\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__19725\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__19722\,
            I => \N__19718\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__19721\,
            I => \N__19715\
        );

    \I__2133\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19712\
        );

    \I__2132\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19709\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__19712\,
            I => \N__19704\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__19709\,
            I => \N__19704\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__19704\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2128\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19697\
        );

    \I__2127\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19694\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__19697\,
            I => \N__19691\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__19694\,
            I => \N__19688\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__19691\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__19688\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2122\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19679\
        );

    \I__2121\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19676\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__19679\,
            I => \N__19673\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__19676\,
            I => \N__19670\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__19673\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2117\ : Odrv12
    port map (
            O => \N__19670\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2116\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19661\
        );

    \I__2115\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19658\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__19661\,
            I => \N__19655\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__19658\,
            I => \N__19652\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__19655\,
            I => \N__19649\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__19652\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__19649\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__19644\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\
        );

    \I__2108\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19638\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__19638\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__2106\ : InMux
    port map (
            O => \N__19635\,
            I => \N__19632\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__19632\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2104\ : InMux
    port map (
            O => \N__19629\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2103\ : InMux
    port map (
            O => \N__19626\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2102\ : InMux
    port map (
            O => \N__19623\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2101\ : InMux
    port map (
            O => \N__19620\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2100\ : InMux
    port map (
            O => \N__19617\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2099\ : InMux
    port map (
            O => \N__19614\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2098\ : InMux
    port map (
            O => \N__19611\,
            I => \N__19607\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__19610\,
            I => \N__19601\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__19607\,
            I => \N__19597\
        );

    \I__2095\ : InMux
    port map (
            O => \N__19606\,
            I => \N__19594\
        );

    \I__2094\ : InMux
    port map (
            O => \N__19605\,
            I => \N__19587\
        );

    \I__2093\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19587\
        );

    \I__2092\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19587\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__19600\,
            I => \N__19583\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__19597\,
            I => \N__19573\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__19594\,
            I => \N__19573\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__19587\,
            I => \N__19573\
        );

    \I__2087\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19570\
        );

    \I__2086\ : InMux
    port map (
            O => \N__19583\,
            I => \N__19561\
        );

    \I__2085\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19561\
        );

    \I__2084\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19561\
        );

    \I__2083\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19561\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__19573\,
            I => \N__19558\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__19570\,
            I => \N__19553\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__19561\,
            I => \N__19553\
        );

    \I__2079\ : Sp12to4
    port map (
            O => \N__19558\,
            I => \N__19548\
        );

    \I__2078\ : Span12Mux_s10_v
    port map (
            O => \N__19553\,
            I => \N__19548\
        );

    \I__2077\ : Odrv12
    port map (
            O => \N__19548\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2076\ : InMux
    port map (
            O => \N__19545\,
            I => \N__19542\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__19542\,
            I => \N__19538\
        );

    \I__2074\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19535\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__19538\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__19535\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__19530\,
            I => \N__19527\
        );

    \I__2070\ : InMux
    port map (
            O => \N__19527\,
            I => \N__19523\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__19526\,
            I => \N__19520\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__19523\,
            I => \N__19517\
        );

    \I__2067\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19514\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__19517\,
            I => \N__19509\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__19514\,
            I => \N__19509\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__19509\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__19506\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_\
        );

    \I__2062\ : InMux
    port map (
            O => \N__19503\,
            I => \N__19498\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__19502\,
            I => \N__19495\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__19501\,
            I => \N__19492\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__19498\,
            I => \N__19488\
        );

    \I__2058\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19481\
        );

    \I__2057\ : InMux
    port map (
            O => \N__19492\,
            I => \N__19481\
        );

    \I__2056\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19481\
        );

    \I__2055\ : Span4Mux_s2_h
    port map (
            O => \N__19488\,
            I => \N__19472\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__19481\,
            I => \N__19472\
        );

    \I__2053\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19469\
        );

    \I__2052\ : InMux
    port map (
            O => \N__19479\,
            I => \N__19462\
        );

    \I__2051\ : InMux
    port map (
            O => \N__19478\,
            I => \N__19462\
        );

    \I__2050\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19462\
        );

    \I__2049\ : Span4Mux_v
    port map (
            O => \N__19472\,
            I => \N__19459\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__19469\,
            I => \N__19454\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__19462\,
            I => \N__19454\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__19459\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2045\ : Odrv12
    port map (
            O => \N__19454\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2044\ : InMux
    port map (
            O => \N__19449\,
            I => \N__19446\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__19446\,
            I => \N__19442\
        );

    \I__2042\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19439\
        );

    \I__2041\ : Span4Mux_v
    port map (
            O => \N__19442\,
            I => \N__19434\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__19439\,
            I => \N__19434\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__19434\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2038\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19428\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__19428\,
            I => \N__19424\
        );

    \I__2036\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19421\
        );

    \I__2035\ : Odrv12
    port map (
            O => \N__19424\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__19421\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2033\ : InMux
    port map (
            O => \N__19416\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2032\ : InMux
    port map (
            O => \N__19413\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2031\ : InMux
    port map (
            O => \N__19410\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2030\ : InMux
    port map (
            O => \N__19407\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2029\ : InMux
    port map (
            O => \N__19404\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2028\ : InMux
    port map (
            O => \N__19401\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2027\ : InMux
    port map (
            O => \N__19398\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2026\ : InMux
    port map (
            O => \N__19395\,
            I => \bfn_2_16_0_\
        );

    \I__2025\ : InMux
    port map (
            O => \N__19392\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2024\ : InMux
    port map (
            O => \N__19389\,
            I => \N__19385\
        );

    \I__2023\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19382\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__19385\,
            I => \N__19378\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__19382\,
            I => \N__19375\
        );

    \I__2020\ : InMux
    port map (
            O => \N__19381\,
            I => \N__19372\
        );

    \I__2019\ : Span4Mux_v
    port map (
            O => \N__19378\,
            I => \N__19369\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__19375\,
            I => \N__19364\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__19372\,
            I => \N__19364\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__19369\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__19364\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2014\ : InMux
    port map (
            O => \N__19359\,
            I => \bfn_2_14_0_\
        );

    \I__2013\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19351\
        );

    \I__2012\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19348\
        );

    \I__2011\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19345\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__19351\,
            I => \N__19342\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__19348\,
            I => \N__19339\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__19345\,
            I => \N__19336\
        );

    \I__2007\ : Span4Mux_v
    port map (
            O => \N__19342\,
            I => \N__19331\
        );

    \I__2006\ : Span4Mux_s2_h
    port map (
            O => \N__19339\,
            I => \N__19331\
        );

    \I__2005\ : Odrv12
    port map (
            O => \N__19336\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__19331\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2003\ : InMux
    port map (
            O => \N__19326\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2002\ : InMux
    port map (
            O => \N__19323\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2001\ : InMux
    port map (
            O => \N__19320\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2000\ : InMux
    port map (
            O => \N__19317\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__1999\ : InMux
    port map (
            O => \N__19314\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__1998\ : InMux
    port map (
            O => \N__19311\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__1997\ : InMux
    port map (
            O => \N__19308\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__1996\ : InMux
    port map (
            O => \N__19305\,
            I => \bfn_2_15_0_\
        );

    \I__1995\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19299\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__19299\,
            I => \N__19296\
        );

    \I__1993\ : Span4Mux_v
    port map (
            O => \N__19296\,
            I => \N__19292\
        );

    \I__1992\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19289\
        );

    \I__1991\ : Span4Mux_s2_h
    port map (
            O => \N__19292\,
            I => \N__19286\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__19289\,
            I => \N__19283\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__19286\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__19283\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1987\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19275\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__19275\,
            I => \N__19272\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__19272\,
            I => \N__19269\
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__19269\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__1983\ : InMux
    port map (
            O => \N__19266\,
            I => \N__19263\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__19263\,
            I => \N__19260\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__19260\,
            I => \N__19257\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__19257\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__1979\ : InMux
    port map (
            O => \N__19254\,
            I => \N__19251\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__19251\,
            I => \N__19248\
        );

    \I__1977\ : Span4Mux_s3_h
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__1976\ : Odrv4
    port map (
            O => \N__19245\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__1975\ : InMux
    port map (
            O => \N__19242\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__1974\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19236\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__19236\,
            I => \N__19233\
        );

    \I__1972\ : Span4Mux_s3_h
    port map (
            O => \N__19233\,
            I => \N__19230\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__19230\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__1970\ : InMux
    port map (
            O => \N__19227\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__1969\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19219\
        );

    \I__1968\ : InMux
    port map (
            O => \N__19223\,
            I => \N__19216\
        );

    \I__1967\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19213\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__19219\,
            I => \N__19210\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__19216\,
            I => \N__19205\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__19213\,
            I => \N__19205\
        );

    \I__1963\ : Span4Mux_s3_h
    port map (
            O => \N__19210\,
            I => \N__19200\
        );

    \I__1962\ : Span4Mux_s3_h
    port map (
            O => \N__19205\,
            I => \N__19200\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__19200\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__1960\ : InMux
    port map (
            O => \N__19197\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__1959\ : InMux
    port map (
            O => \N__19194\,
            I => \N__19188\
        );

    \I__1958\ : InMux
    port map (
            O => \N__19193\,
            I => \N__19183\
        );

    \I__1957\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19183\
        );

    \I__1956\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19180\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__19188\,
            I => \N__19177\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__19183\,
            I => \N__19172\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__19180\,
            I => \N__19172\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__19177\,
            I => \N__19167\
        );

    \I__1951\ : Span4Mux_v
    port map (
            O => \N__19172\,
            I => \N__19167\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__19167\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__1949\ : InMux
    port map (
            O => \N__19164\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__19161\,
            I => \N__19158\
        );

    \I__1947\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19153\
        );

    \I__1946\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19150\
        );

    \I__1945\ : InMux
    port map (
            O => \N__19156\,
            I => \N__19147\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__19153\,
            I => \N__19144\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__19150\,
            I => \N__19141\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__19147\,
            I => \N__19138\
        );

    \I__1941\ : Span4Mux_s2_h
    port map (
            O => \N__19144\,
            I => \N__19133\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__19141\,
            I => \N__19133\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__19138\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__19133\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__1937\ : InMux
    port map (
            O => \N__19128\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__1936\ : InMux
    port map (
            O => \N__19125\,
            I => \N__19120\
        );

    \I__1935\ : InMux
    port map (
            O => \N__19124\,
            I => \N__19117\
        );

    \I__1934\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19114\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__19120\,
            I => \N__19111\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__19117\,
            I => \N__19106\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__19114\,
            I => \N__19106\
        );

    \I__1930\ : Span4Mux_v
    port map (
            O => \N__19111\,
            I => \N__19101\
        );

    \I__1929\ : Span4Mux_v
    port map (
            O => \N__19106\,
            I => \N__19101\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__19101\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__1927\ : InMux
    port map (
            O => \N__19098\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__1926\ : InMux
    port map (
            O => \N__19095\,
            I => \N__19090\
        );

    \I__1925\ : InMux
    port map (
            O => \N__19094\,
            I => \N__19087\
        );

    \I__1924\ : InMux
    port map (
            O => \N__19093\,
            I => \N__19084\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__19090\,
            I => \N__19081\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__19087\,
            I => \N__19076\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__19084\,
            I => \N__19076\
        );

    \I__1920\ : Span4Mux_v
    port map (
            O => \N__19081\,
            I => \N__19071\
        );

    \I__1919\ : Span4Mux_v
    port map (
            O => \N__19076\,
            I => \N__19071\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__19071\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__1917\ : InMux
    port map (
            O => \N__19068\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__19065\,
            I => \N__19062\
        );

    \I__1915\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19058\
        );

    \I__1914\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19055\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__19058\,
            I => \N__19050\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__19055\,
            I => \N__19050\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__19050\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1910\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19044\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__19044\,
            I => \N__19041\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__19041\,
            I => \N__19038\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__19038\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__1906\ : InMux
    port map (
            O => \N__19035\,
            I => \N__19029\
        );

    \I__1905\ : InMux
    port map (
            O => \N__19034\,
            I => \N__19029\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__19029\,
            I => \N__19026\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__19026\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__19023\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\
        );

    \I__1901\ : InMux
    port map (
            O => \N__19020\,
            I => \N__19017\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__19017\,
            I => \N__19014\
        );

    \I__1899\ : Span4Mux_v
    port map (
            O => \N__19014\,
            I => \N__19011\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__19011\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__1897\ : InMux
    port map (
            O => \N__19008\,
            I => \N__19004\
        );

    \I__1896\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19001\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__19004\,
            I => \N__18996\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__19001\,
            I => \N__18996\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__18996\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__18993\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\
        );

    \I__1891\ : CascadeMux
    port map (
            O => \N__18990\,
            I => \N__18987\
        );

    \I__1890\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18984\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__18984\,
            I => \N__18981\
        );

    \I__1888\ : Span4Mux_h
    port map (
            O => \N__18981\,
            I => \N__18978\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__18978\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__18975\,
            I => \N__18972\
        );

    \I__1885\ : InMux
    port map (
            O => \N__18972\,
            I => \N__18968\
        );

    \I__1884\ : InMux
    port map (
            O => \N__18971\,
            I => \N__18965\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__18968\,
            I => \N__18960\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__18965\,
            I => \N__18960\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__18960\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__1880\ : InMux
    port map (
            O => \N__18957\,
            I => \N__18954\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__18954\,
            I => \N__18951\
        );

    \I__1878\ : Odrv12
    port map (
            O => \N__18951\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__1877\ : InMux
    port map (
            O => \N__18948\,
            I => \N__18945\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__18945\,
            I => \N__18941\
        );

    \I__1875\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18938\
        );

    \I__1874\ : Span4Mux_h
    port map (
            O => \N__18941\,
            I => \N__18935\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__18938\,
            I => \N__18932\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__18935\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1871\ : Odrv4
    port map (
            O => \N__18932\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1870\ : InMux
    port map (
            O => \N__18927\,
            I => \N__18924\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__18924\,
            I => \N__18921\
        );

    \I__1868\ : Odrv12
    port map (
            O => \N__18921\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__18918\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__1866\ : InMux
    port map (
            O => \N__18915\,
            I => \N__18912\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__18912\,
            I => \N__18909\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__18909\,
            I => \N__18906\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__18906\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__18903\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\
        );

    \I__1861\ : InMux
    port map (
            O => \N__18900\,
            I => \N__18897\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__18897\,
            I => \N__18894\
        );

    \I__1859\ : Span4Mux_h
    port map (
            O => \N__18894\,
            I => \N__18891\
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__18891\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__18888\,
            I => \N__18885\
        );

    \I__1856\ : InMux
    port map (
            O => \N__18885\,
            I => \N__18877\
        );

    \I__1855\ : InMux
    port map (
            O => \N__18884\,
            I => \N__18874\
        );

    \I__1854\ : InMux
    port map (
            O => \N__18883\,
            I => \N__18867\
        );

    \I__1853\ : InMux
    port map (
            O => \N__18882\,
            I => \N__18867\
        );

    \I__1852\ : InMux
    port map (
            O => \N__18881\,
            I => \N__18867\
        );

    \I__1851\ : InMux
    port map (
            O => \N__18880\,
            I => \N__18864\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__18877\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__18874\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__18867\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__18864\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__18855\,
            I => \current_shift_inst.PI_CTRL.N_118_cascade_\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__18852\,
            I => \N__18848\
        );

    \I__1844\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18844\
        );

    \I__1843\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18839\
        );

    \I__1842\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18839\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__18844\,
            I => \N__18836\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__18839\,
            I => \N__18831\
        );

    \I__1839\ : Span4Mux_v
    port map (
            O => \N__18836\,
            I => \N__18831\
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__18831\,
            I => pwm_duty_input_9
        );

    \I__1837\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18822\
        );

    \I__1836\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18822\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__18822\,
            I => \N__18819\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__18819\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__18816\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\
        );

    \I__1832\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18810\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__18810\,
            I => \N__18807\
        );

    \I__1830\ : Odrv12
    port map (
            O => \N__18807\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__1829\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18800\
        );

    \I__1828\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18797\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__18800\,
            I => \N__18794\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__18797\,
            I => \N__18791\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__18794\,
            I => \N__18788\
        );

    \I__1824\ : Span4Mux_h
    port map (
            O => \N__18791\,
            I => \N__18785\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__18788\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__18785\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__18780\,
            I => \N__18777\
        );

    \I__1820\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18774\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__18774\,
            I => \N__18771\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__18771\,
            I => \N__18768\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__18768\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__1816\ : InMux
    port map (
            O => \N__18765\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__1815\ : InMux
    port map (
            O => \N__18762\,
            I => \N__18759\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__18759\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__1813\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18753\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__18753\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__1811\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18747\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__18747\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__18744\,
            I => \current_shift_inst.PI_CTRL.N_94_cascade_\
        );

    \I__1808\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18736\
        );

    \I__1807\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18731\
        );

    \I__1806\ : InMux
    port map (
            O => \N__18739\,
            I => \N__18731\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__18736\,
            I => \current_shift_inst.PI_CTRL.N_120\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__18731\,
            I => \current_shift_inst.PI_CTRL.N_120\
        );

    \I__1803\ : InMux
    port map (
            O => \N__18726\,
            I => \N__18723\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__18723\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__18720\,
            I => \N__18717\
        );

    \I__1800\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18713\
        );

    \I__1799\ : InMux
    port map (
            O => \N__18716\,
            I => \N__18710\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__18713\,
            I => \N__18705\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__18710\,
            I => \N__18705\
        );

    \I__1796\ : Span4Mux_h
    port map (
            O => \N__18705\,
            I => \N__18702\
        );

    \I__1795\ : Span4Mux_v
    port map (
            O => \N__18702\,
            I => \N__18699\
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__18699\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__18696\,
            I => \current_shift_inst.PI_CTRL.N_98_cascade_\
        );

    \I__1792\ : InMux
    port map (
            O => \N__18693\,
            I => \N__18689\
        );

    \I__1791\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18686\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__18689\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__18686\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__18681\,
            I => \N__18677\
        );

    \I__1787\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18669\
        );

    \I__1786\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18669\
        );

    \I__1785\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18669\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__18669\,
            I => \N__18666\
        );

    \I__1783\ : Span12Mux_h
    port map (
            O => \N__18666\,
            I => \N__18663\
        );

    \I__1782\ : Odrv12
    port map (
            O => \N__18663\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1781\ : InMux
    port map (
            O => \N__18660\,
            I => \N__18657\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__18657\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__1779\ : InMux
    port map (
            O => \N__18654\,
            I => \N__18651\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__18651\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__1777\ : InMux
    port map (
            O => \N__18648\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__1776\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18642\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__18642\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__1774\ : InMux
    port map (
            O => \N__18639\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__1773\ : InMux
    port map (
            O => \N__18636\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__1772\ : InMux
    port map (
            O => \N__18633\,
            I => \N__18630\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__18630\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__1770\ : InMux
    port map (
            O => \N__18627\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__1769\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18621\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__18621\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__1767\ : InMux
    port map (
            O => \N__18618\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__1766\ : InMux
    port map (
            O => \N__18615\,
            I => \N__18612\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__18612\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__1764\ : InMux
    port map (
            O => \N__18609\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__1763\ : InMux
    port map (
            O => \N__18606\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__1762\ : InMux
    port map (
            O => \N__18603\,
            I => \bfn_2_8_0_\
        );

    \I__1761\ : InMux
    port map (
            O => \N__18600\,
            I => \N__18597\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__18597\,
            I => un7_start_stop_0_a3
        );

    \I__1759\ : InMux
    port map (
            O => \N__18594\,
            I => \N__18591\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__18591\,
            I => \N_34_i_i\
        );

    \I__1757\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18585\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__18585\,
            I => \N__18582\
        );

    \I__1755\ : Glb2LocalMux
    port map (
            O => \N__18582\,
            I => \N__18579\
        );

    \I__1754\ : GlobalMux
    port map (
            O => \N__18579\,
            I => clk_12mhz
        );

    \I__1753\ : IoInMux
    port map (
            O => \N__18576\,
            I => \N__18573\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__18573\,
            I => \N__18570\
        );

    \I__1751\ : IoSpan4Mux
    port map (
            O => \N__18570\,
            I => \N__18567\
        );

    \I__1750\ : Span4Mux_s0_v
    port map (
            O => \N__18567\,
            I => \N__18564\
        );

    \I__1749\ : Span4Mux_h
    port map (
            O => \N__18564\,
            I => \N__18561\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__18561\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__1747\ : InMux
    port map (
            O => \N__18558\,
            I => \N__18555\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__18555\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__1745\ : InMux
    port map (
            O => \N__18552\,
            I => \N__18549\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__18549\,
            I => \N__18546\
        );

    \I__1743\ : Odrv12
    port map (
            O => \N__18546\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__1742\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18540\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__18540\,
            I => \N__18537\
        );

    \I__1740\ : Odrv12
    port map (
            O => \N__18537\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__1739\ : InMux
    port map (
            O => \N__18534\,
            I => \N__18531\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__18531\,
            I => \N__18528\
        );

    \I__1737\ : Odrv12
    port map (
            O => \N__18528\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__1736\ : InMux
    port map (
            O => \N__18525\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__1735\ : InMux
    port map (
            O => \N__18522\,
            I => \N__18519\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__18519\,
            I => \N__18516\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__18516\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__1732\ : InMux
    port map (
            O => \N__18513\,
            I => \N__18510\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__18510\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__18507\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__1729\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18501\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__18501\,
            I => \N__18498\
        );

    \I__1727\ : Odrv12
    port map (
            O => \N__18498\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__1726\ : InMux
    port map (
            O => \N__18495\,
            I => \bfn_1_15_0_\
        );

    \I__1725\ : InMux
    port map (
            O => \N__18492\,
            I => \N__18489\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__18489\,
            I => \N__18486\
        );

    \I__1723\ : Odrv12
    port map (
            O => \N__18486\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__1722\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18480\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__18480\,
            I => \N__18477\
        );

    \I__1720\ : Odrv12
    port map (
            O => \N__18477\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__1719\ : InMux
    port map (
            O => \N__18474\,
            I => \N__18471\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__18471\,
            I => \N__18468\
        );

    \I__1717\ : Odrv12
    port map (
            O => \N__18468\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__1716\ : InMux
    port map (
            O => \N__18465\,
            I => \N__18462\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__18462\,
            I => \N__18459\
        );

    \I__1714\ : Odrv12
    port map (
            O => \N__18459\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__1713\ : InMux
    port map (
            O => \N__18456\,
            I => \N__18453\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__18453\,
            I => \N__18450\
        );

    \I__1711\ : Odrv12
    port map (
            O => \N__18450\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__1710\ : InMux
    port map (
            O => \N__18447\,
            I => \N__18444\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__18444\,
            I => \N__18441\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__18441\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__1707\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18435\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__18435\,
            I => \N__18432\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__18432\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__1704\ : InMux
    port map (
            O => \N__18429\,
            I => \N__18426\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__18426\,
            I => \N__18423\
        );

    \I__1702\ : Odrv12
    port map (
            O => \N__18423\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__1701\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18417\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__18417\,
            I => \N__18414\
        );

    \I__1699\ : Span4Mux_h
    port map (
            O => \N__18414\,
            I => \N__18411\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__18411\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1697\ : InMux
    port map (
            O => \N__18408\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__1696\ : InMux
    port map (
            O => \N__18405\,
            I => \N__18402\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__18402\,
            I => \N__18399\
        );

    \I__1694\ : Span4Mux_h
    port map (
            O => \N__18399\,
            I => \N__18396\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__18396\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1692\ : InMux
    port map (
            O => \N__18393\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__1691\ : InMux
    port map (
            O => \N__18390\,
            I => \N__18387\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__18387\,
            I => \N__18384\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__18384\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1688\ : InMux
    port map (
            O => \N__18381\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__1687\ : InMux
    port map (
            O => \N__18378\,
            I => \N__18375\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__18375\,
            I => \N__18372\
        );

    \I__1685\ : Odrv12
    port map (
            O => \N__18372\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__1684\ : InMux
    port map (
            O => \N__18369\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__18366\,
            I => \N__18363\
        );

    \I__1682\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18360\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__18360\,
            I => \N__18357\
        );

    \I__1680\ : Odrv12
    port map (
            O => \N__18357\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__1679\ : InMux
    port map (
            O => \N__18354\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__1678\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18348\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__18348\,
            I => \N__18345\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__18345\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__1675\ : InMux
    port map (
            O => \N__18342\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__1674\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18336\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__18336\,
            I => \N__18333\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__18333\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__1671\ : InMux
    port map (
            O => \N__18330\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__18327\,
            I => \N__18324\
        );

    \I__1669\ : InMux
    port map (
            O => \N__18324\,
            I => \N__18321\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__18321\,
            I => \N__18318\
        );

    \I__1667\ : Span4Mux_v
    port map (
            O => \N__18318\,
            I => \N__18315\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__18315\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1665\ : InMux
    port map (
            O => \N__18312\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1664\ : InMux
    port map (
            O => \N__18309\,
            I => \N__18306\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__18306\,
            I => \N__18303\
        );

    \I__1662\ : Span4Mux_v
    port map (
            O => \N__18303\,
            I => \N__18300\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__18300\,
            I => \N__18297\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__18297\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1659\ : InMux
    port map (
            O => \N__18294\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__18291\,
            I => \N__18288\
        );

    \I__1657\ : InMux
    port map (
            O => \N__18288\,
            I => \N__18285\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__18285\,
            I => \N__18282\
        );

    \I__1655\ : Span4Mux_v
    port map (
            O => \N__18282\,
            I => \N__18279\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__18279\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1653\ : InMux
    port map (
            O => \N__18276\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__1652\ : InMux
    port map (
            O => \N__18273\,
            I => \N__18270\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__18270\,
            I => \N__18267\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__18267\,
            I => \N__18264\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__18264\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__1648\ : InMux
    port map (
            O => \N__18261\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__18258\,
            I => \N__18255\
        );

    \I__1646\ : InMux
    port map (
            O => \N__18255\,
            I => \N__18252\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__18252\,
            I => \N__18249\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__18249\,
            I => \N__18246\
        );

    \I__1643\ : Span4Mux_s1_h
    port map (
            O => \N__18246\,
            I => \N__18243\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__18243\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__1641\ : InMux
    port map (
            O => \N__18240\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__1640\ : InMux
    port map (
            O => \N__18237\,
            I => \N__18234\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__18234\,
            I => \N__18231\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__18231\,
            I => \N__18228\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__18228\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__1636\ : InMux
    port map (
            O => \N__18225\,
            I => \N__18222\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__18222\,
            I => \N__18218\
        );

    \I__1634\ : InMux
    port map (
            O => \N__18221\,
            I => \N__18215\
        );

    \I__1633\ : Span4Mux_v
    port map (
            O => \N__18218\,
            I => \N__18207\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__18215\,
            I => \N__18207\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__18214\,
            I => \N__18204\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__18213\,
            I => \N__18200\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__18212\,
            I => \N__18196\
        );

    \I__1628\ : Span4Mux_v
    port map (
            O => \N__18207\,
            I => \N__18192\
        );

    \I__1627\ : InMux
    port map (
            O => \N__18204\,
            I => \N__18179\
        );

    \I__1626\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18179\
        );

    \I__1625\ : InMux
    port map (
            O => \N__18200\,
            I => \N__18179\
        );

    \I__1624\ : InMux
    port map (
            O => \N__18199\,
            I => \N__18179\
        );

    \I__1623\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18179\
        );

    \I__1622\ : InMux
    port map (
            O => \N__18195\,
            I => \N__18179\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__18192\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__18179\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1619\ : InMux
    port map (
            O => \N__18174\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__1618\ : InMux
    port map (
            O => \N__18171\,
            I => \N__18168\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__18168\,
            I => \N__18165\
        );

    \I__1616\ : Odrv12
    port map (
            O => \N__18165\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__1615\ : InMux
    port map (
            O => \N__18162\,
            I => \bfn_1_13_0_\
        );

    \I__1614\ : InMux
    port map (
            O => \N__18159\,
            I => \N__18156\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__18156\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\
        );

    \I__1612\ : InMux
    port map (
            O => \N__18153\,
            I => \N__18150\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__18150\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__18147\,
            I => \N__18144\
        );

    \I__1609\ : InMux
    port map (
            O => \N__18144\,
            I => \N__18141\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__18141\,
            I => \N__18138\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__18138\,
            I => \N__18135\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__18135\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1605\ : InMux
    port map (
            O => \N__18132\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1604\ : InMux
    port map (
            O => \N__18129\,
            I => \N__18126\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__18126\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__18123\,
            I => \N__18120\
        );

    \I__1601\ : InMux
    port map (
            O => \N__18120\,
            I => \N__18117\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__18117\,
            I => \N__18114\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__18114\,
            I => \N__18111\
        );

    \I__1598\ : Span4Mux_s1_h
    port map (
            O => \N__18111\,
            I => \N__18108\
        );

    \I__1597\ : Odrv4
    port map (
            O => \N__18108\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1596\ : InMux
    port map (
            O => \N__18105\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1595\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18099\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__18099\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__18096\,
            I => \N__18093\
        );

    \I__1592\ : InMux
    port map (
            O => \N__18093\,
            I => \N__18090\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__18090\,
            I => \N__18087\
        );

    \I__1590\ : Span4Mux_v
    port map (
            O => \N__18087\,
            I => \N__18084\
        );

    \I__1589\ : Odrv4
    port map (
            O => \N__18084\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1588\ : InMux
    port map (
            O => \N__18081\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1587\ : InMux
    port map (
            O => \N__18078\,
            I => \N__18075\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__18075\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__18072\,
            I => \N__18069\
        );

    \I__1584\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18066\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__18066\,
            I => \N__18063\
        );

    \I__1582\ : Span4Mux_v
    port map (
            O => \N__18063\,
            I => \N__18060\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__18060\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__1580\ : InMux
    port map (
            O => \N__18057\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__1579\ : InMux
    port map (
            O => \N__18054\,
            I => \N__18051\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__18051\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__18048\,
            I => \N__18045\
        );

    \I__1576\ : InMux
    port map (
            O => \N__18045\,
            I => \N__18042\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__18042\,
            I => \N__18039\
        );

    \I__1574\ : Span4Mux_v
    port map (
            O => \N__18039\,
            I => \N__18036\
        );

    \I__1573\ : Odrv4
    port map (
            O => \N__18036\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__1572\ : InMux
    port map (
            O => \N__18033\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__1571\ : InMux
    port map (
            O => \N__18030\,
            I => \N__18027\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__18027\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__18024\,
            I => \N__18021\
        );

    \I__1568\ : InMux
    port map (
            O => \N__18021\,
            I => \N__18018\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__18018\,
            I => \N__18015\
        );

    \I__1566\ : Span4Mux_v
    port map (
            O => \N__18015\,
            I => \N__18012\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__18012\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__1564\ : InMux
    port map (
            O => \N__18009\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__1563\ : InMux
    port map (
            O => \N__18006\,
            I => \N__18003\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__18003\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__18000\,
            I => \N__17997\
        );

    \I__1560\ : InMux
    port map (
            O => \N__17997\,
            I => \N__17994\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__17994\,
            I => \N__17991\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__17991\,
            I => \N__17988\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__17988\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__1556\ : InMux
    port map (
            O => \N__17985\,
            I => \bfn_1_12_0_\
        );

    \I__1555\ : InMux
    port map (
            O => \N__17982\,
            I => \N__17979\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__17979\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__1553\ : CascadeMux
    port map (
            O => \N__17976\,
            I => \N__17973\
        );

    \I__1552\ : InMux
    port map (
            O => \N__17973\,
            I => \N__17970\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__17970\,
            I => \N__17967\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__17967\,
            I => \N__17964\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__17964\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1548\ : InMux
    port map (
            O => \N__17961\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__17958\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__17955\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\
        );

    \I__1545\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17947\
        );

    \I__1544\ : InMux
    port map (
            O => \N__17951\,
            I => \N__17942\
        );

    \I__1543\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17942\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__17947\,
            I => \N__17939\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__17942\,
            I => pwm_duty_input_6
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__17939\,
            I => pwm_duty_input_6
        );

    \I__1539\ : InMux
    port map (
            O => \N__17934\,
            I => \N__17929\
        );

    \I__1538\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17924\
        );

    \I__1537\ : InMux
    port map (
            O => \N__17932\,
            I => \N__17924\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__17929\,
            I => \N__17921\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__17924\,
            I => pwm_duty_input_7
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__17921\,
            I => pwm_duty_input_7
        );

    \I__1533\ : InMux
    port map (
            O => \N__17916\,
            I => \N__17911\
        );

    \I__1532\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17906\
        );

    \I__1531\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17906\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__17911\,
            I => \N__17903\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__17906\,
            I => pwm_duty_input_5
        );

    \I__1528\ : Odrv4
    port map (
            O => \N__17903\,
            I => pwm_duty_input_5
        );

    \I__1527\ : InMux
    port map (
            O => \N__17898\,
            I => \N__17895\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__17895\,
            I => \N__17890\
        );

    \I__1525\ : InMux
    port map (
            O => \N__17894\,
            I => \N__17885\
        );

    \I__1524\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17885\
        );

    \I__1523\ : Span4Mux_v
    port map (
            O => \N__17890\,
            I => \N__17882\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__17885\,
            I => pwm_duty_input_4
        );

    \I__1521\ : Odrv4
    port map (
            O => \N__17882\,
            I => pwm_duty_input_4
        );

    \I__1520\ : InMux
    port map (
            O => \N__17877\,
            I => \N__17872\
        );

    \I__1519\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17869\
        );

    \I__1518\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17866\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__17872\,
            I => \N__17863\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__17869\,
            I => pwm_duty_input_8
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__17866\,
            I => pwm_duty_input_8
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__17863\,
            I => pwm_duty_input_8
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__17856\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\
        );

    \I__1512\ : InMux
    port map (
            O => \N__17853\,
            I => \N__17848\
        );

    \I__1511\ : InMux
    port map (
            O => \N__17852\,
            I => \N__17843\
        );

    \I__1510\ : InMux
    port map (
            O => \N__17851\,
            I => \N__17843\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__17848\,
            I => \N__17840\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__17843\,
            I => pwm_duty_input_3
        );

    \I__1507\ : Odrv4
    port map (
            O => \N__17840\,
            I => pwm_duty_input_3
        );

    \I__1506\ : InMux
    port map (
            O => \N__17835\,
            I => \N__17832\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__17832\,
            I => \N__17829\
        );

    \I__1504\ : Span4Mux_v
    port map (
            O => \N__17829\,
            I => \N__17826\
        );

    \I__1503\ : Odrv4
    port map (
            O => \N__17826\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__17823\,
            I => \N__17820\
        );

    \I__1501\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17817\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__17817\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1499\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17811\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__17811\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__17808\,
            I => \N__17805\
        );

    \I__1496\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17802\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__17802\,
            I => \N__17799\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__17799\,
            I => \N__17796\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__17796\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1492\ : InMux
    port map (
            O => \N__17793\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1491\ : InMux
    port map (
            O => \N__17790\,
            I => \N__17786\
        );

    \I__1490\ : InMux
    port map (
            O => \N__17789\,
            I => \N__17783\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__17786\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__17783\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__17778\,
            I => \N__17775\
        );

    \I__1486\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17772\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__17772\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_counter_cry_8,
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_3_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_3_10_0_\
        );

    \IN_MUX_bfv_3_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_3_11_0_\
        );

    \IN_MUX_bfv_4_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_6_0_\
        );

    \IN_MUX_bfv_4_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_4_7_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_10_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_11_0_\
        );

    \IN_MUX_bfv_10_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_10_12_0_\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_16_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_16_14_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_15_25_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_14_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_14_27_0_\
        );

    \IN_MUX_bfv_14_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_14_28_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_7\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_15\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_23\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_2_16_0_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__39831\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_461_i_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__31110\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_185_i_g\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__28527\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_463_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__34290\,
            CLKHFEN => \N__34292\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__34291\,
            RGB2PWM => \N__18594\,
            RGB1 => rgb_g_wire,
            CURREN => \N__34566\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__18600\,
            RGB0PWM => \N__45622\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__18225\,
            in1 => \N__17789\,
            in2 => \_gnd_net_\,
            in3 => \N__20199\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19611\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46077\,
            ce => \N__24873\,
            sr => \N__45526\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__20201\,
            in1 => \N__20306\,
            in2 => \N__20414\,
            in3 => \N__18762\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46075\,
            ce => 'H',
            sr => \N__45534\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__17790\,
            in1 => \N__20200\,
            in2 => \N__17778\,
            in3 => \N__18221\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19266\,
            in2 => \_gnd_net_\,
            in3 => \N__18741\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46073\,
            ce => \N__24867\,
            sr => \N__45541\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18740\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19239\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46071\,
            ce => \N__24824\,
            sr => \N__45548\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__18884\,
            in1 => \N__18726\,
            in2 => \N__18720\,
            in3 => \N__19194\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46071\,
            ce => \N__24824\,
            sr => \N__45548\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__19224\,
            in1 => \N__18750\,
            in2 => \_gnd_net_\,
            in3 => \N__18693\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46071\,
            ce => \N__24824\,
            sr => \N__45548\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101110"
        )
    port map (
            in0 => \N__19389\,
            in1 => \N__19503\,
            in2 => \N__18888\,
            in3 => \N__19606\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46071\,
            ce => \N__24824\,
            sr => \N__45548\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19254\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18739\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46071\,
            ce => \N__24824\,
            sr => \N__45548\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__19156\,
            in1 => \N__19491\,
            in2 => \N__19610\,
            in3 => \N__18883\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46066\,
            ce => \N__24866\,
            sr => \N__45555\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__18882\,
            in1 => \N__19605\,
            in2 => \N__19502\,
            in3 => \N__19095\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46066\,
            ce => \N__24866\,
            sr => \N__45555\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17932\,
            in2 => \_gnd_net_\,
            in3 => \N__17914\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__17875\,
            in1 => \N__18847\,
            in2 => \N__17958\,
            in3 => \N__17950\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110001"
        )
    port map (
            in0 => \N__17852\,
            in1 => \N__17893\,
            in2 => \N__17955\,
            in3 => \N__33147\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__18881\,
            in1 => \N__19604\,
            in2 => \N__19501\,
            in3 => \N__19125\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46066\,
            ce => \N__24866\,
            sr => \N__45555\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17951\,
            in1 => \N__17933\,
            in2 => \N__18852\,
            in3 => \N__17915\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__17894\,
            in1 => \N__17876\,
            in2 => \N__17856\,
            in3 => \N__17851\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17835\,
            in2 => \N__17823\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17814\,
            in2 => \N__17808\,
            in3 => \N__17793\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18153\,
            in2 => \N__18147\,
            in3 => \N__18132\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18129\,
            in2 => \N__18123\,
            in3 => \N__18105\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18102\,
            in2 => \N__18096\,
            in3 => \N__18081\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18078\,
            in2 => \N__18072\,
            in3 => \N__18057\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18054\,
            in2 => \N__18048\,
            in3 => \N__18033\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18030\,
            in2 => \N__18024\,
            in3 => \N__18009\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18006\,
            in2 => \N__18000\,
            in3 => \N__17985\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17982\,
            in2 => \N__17976\,
            in3 => \N__17961\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18195\,
            in2 => \N__18327\,
            in3 => \N__18312\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18309\,
            in2 => \N__18212\,
            in3 => \N__18294\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18199\,
            in2 => \N__18291\,
            in3 => \N__18276\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18273\,
            in2 => \N__18213\,
            in3 => \N__18261\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18203\,
            in2 => \N__18258\,
            in3 => \N__18240\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18237\,
            in2 => \N__18214\,
            in3 => \N__18174\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18171\,
            in1 => \N__18522\,
            in2 => \_gnd_net_\,
            in3 => \N__18162\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIKH62_13_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19700\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIR3F5_14_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19541\,
            in1 => \N__19892\,
            in2 => \N__19530\,
            in3 => \N__18159\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20471\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18420\,
            in2 => \_gnd_net_\,
            in3 => \N__18408\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18405\,
            in2 => \_gnd_net_\,
            in3 => \N__18393\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18390\,
            in2 => \_gnd_net_\,
            in3 => \N__18381\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18378\,
            in2 => \_gnd_net_\,
            in3 => \N__18369\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34449\,
            in2 => \N__18366\,
            in3 => \N__18354\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18351\,
            in2 => \N__34556\,
            in3 => \N__18342\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18339\,
            in2 => \N__34557\,
            in3 => \N__18330\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18504\,
            in2 => \_gnd_net_\,
            in3 => \N__18495\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18492\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18483\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18474\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18465\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18456\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18447\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18438\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18429\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18552\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18543\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18534\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18525\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIV2LD_8_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19355\,
            in2 => \_gnd_net_\,
            in3 => \N__19381\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19094\,
            in1 => \N__19124\,
            in2 => \N__19161\,
            in3 => \N__18513\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_11_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19914\,
            in1 => \N__19971\,
            in2 => \N__19959\,
            in3 => \N__19932\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19093\,
            in2 => \_gnd_net_\,
            in3 => \N__19157\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__19356\,
            in1 => \N__19123\,
            in2 => \N__18507\,
            in3 => \N__19388\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_start_stop_0_a3_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29399\,
            in2 => \_gnd_net_\,
            in3 => \N__45620\,
            lcout => un7_start_stop_0_a3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.N_34_i_i_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__45621\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29403\,
            lcout => \N_34_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18588\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_2_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18558\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46076\,
            ce => 'H',
            sr => \N__45518\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__20409\,
            in1 => \N__20335\,
            in2 => \N__20277\,
            in3 => \N__18615\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46076\,
            ce => 'H',
            sr => \N__45518\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__20250\,
            in1 => \N__20407\,
            in2 => \N__20340\,
            in3 => \N__18633\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46076\,
            ce => 'H',
            sr => \N__45518\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__20406\,
            in1 => \N__20330\,
            in2 => \N__20275\,
            in3 => \N__18645\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46076\,
            ce => 'H',
            sr => \N__45518\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__18654\,
            in1 => \N__20251\,
            in2 => \N__20421\,
            in3 => \N__20329\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46076\,
            ce => 'H',
            sr => \N__45518\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__20408\,
            in1 => \N__20334\,
            in2 => \N__20276\,
            in3 => \N__18624\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46076\,
            ce => 'H',
            sr => \N__45518\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18927\,
            in2 => \N__20541\,
            in3 => \N__20540\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20457\,
            in2 => \_gnd_net_\,
            in3 => \N__18648\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18756\,
            in2 => \_gnd_net_\,
            in3 => \N__18639\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18957\,
            in2 => \_gnd_net_\,
            in3 => \N__18636\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19278\,
            in2 => \_gnd_net_\,
            in3 => \N__18627\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18813\,
            in2 => \_gnd_net_\,
            in3 => \N__18618\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19047\,
            in2 => \_gnd_net_\,
            in3 => \N__18609\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19020\,
            in2 => \_gnd_net_\,
            in3 => \N__18606\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18990\,
            in3 => \N__18603\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__20676\,
            in1 => \N__20536\,
            in2 => \N__18780\,
            in3 => \N__18765\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__18804\,
            in1 => \N__20874\,
            in2 => \N__20853\,
            in3 => \N__20535\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__19478\,
            in1 => \N__19582\,
            in2 => \N__18681\,
            in3 => \N__19192\,
            lcout => \current_shift_inst.PI_CTRL.N_94\,
            ltout => \current_shift_inst.PI_CTRL.N_94_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__19223\,
            in1 => \N__18660\,
            in2 => \N__18744\,
            in3 => \N__18692\,
            lcout => \current_shift_inst.PI_CTRL.N_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__19193\,
            in1 => \N__18680\,
            in2 => \N__19600\,
            in3 => \N__19479\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19191\,
            in2 => \_gnd_net_\,
            in3 => \N__19222\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__18716\,
            in1 => \N__19581\,
            in2 => \N__18696\,
            in3 => \N__18880\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__19580\,
            in1 => \N__18676\,
            in2 => \_gnd_net_\,
            in3 => \N__19477\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPN72_23_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19682\,
            in2 => \_gnd_net_\,
            in3 => \N__19665\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_10_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19860\,
            in1 => \N__19431\,
            in2 => \N__18918\,
            in3 => \N__19449\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18915\,
            in1 => \N__19791\,
            in2 => \N__18903\,
            in3 => \N__18900\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => \current_shift_inst.PI_CTRL.N_118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__19586\,
            in1 => \N__19354\,
            in2 => \N__18855\,
            in3 => \N__19480\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46063\,
            ce => \N__24872\,
            sr => \N__45549\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20748\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19061\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20574\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18944\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18827\,
            in2 => \_gnd_net_\,
            in3 => \N__20769\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__18828\,
            in1 => \N__20757\,
            in2 => \N__18816\,
            in3 => \N__20533\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18971\,
            in2 => \_gnd_net_\,
            in3 => \N__20837\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20873\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18803\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19295\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__20730\,
            in1 => \N__20747\,
            in2 => \N__19065\,
            in3 => \N__20516\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20721\,
            in2 => \_gnd_net_\,
            in3 => \N__19034\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__19035\,
            in1 => \N__20709\,
            in2 => \N__19023\,
            in3 => \N__20517\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20700\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__19008\,
            in1 => \N__20518\,
            in2 => \N__18993\,
            in3 => \N__20688\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__20514\,
            in1 => \N__20817\,
            in2 => \N__18975\,
            in3 => \N__20836\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__20573\,
            in1 => \N__18948\,
            in2 => \N__20556\,
            in3 => \N__20513\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__20515\,
            in1 => \N__20801\,
            in2 => \N__20784\,
            in3 => \N__19302\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21426\,
            in2 => \N__21396\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__46055\,
            ce => \N__24862\,
            sr => \N__45565\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21384\,
            in2 => \N__20973\,
            in3 => \N__19242\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__46055\,
            ce => \N__24862\,
            sr => \N__45565\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21624\,
            in2 => \N__24150\,
            in3 => \N__19227\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__46055\,
            ce => \N__24862\,
            sr => \N__45565\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21591\,
            in2 => \N__20886\,
            in3 => \N__19197\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__46055\,
            ce => \N__24862\,
            sr => \N__45565\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21549\,
            in2 => \N__20907\,
            in3 => \N__19164\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__46055\,
            ce => \N__24862\,
            sr => \N__45565\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21513\,
            in2 => \N__20898\,
            in3 => \N__19128\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__46055\,
            ce => \N__24862\,
            sr => \N__45565\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22284\,
            in2 => \N__20988\,
            in3 => \N__19098\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__46055\,
            ce => \N__24862\,
            sr => \N__45565\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20979\,
            in2 => \N__22740\,
            in3 => \N__19068\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__46055\,
            ce => \N__24862\,
            sr => \N__45565\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23050\,
            in2 => \N__20937\,
            in3 => \N__19359\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__46047\,
            ce => \N__24812\,
            sr => \N__45569\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21463\,
            in2 => \N__20946\,
            in3 => \N__19326\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__46047\,
            ce => \N__24812\,
            sr => \N__45569\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21006\,
            in2 => \N__22863\,
            in3 => \N__19323\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__46047\,
            ce => \N__24812\,
            sr => \N__45569\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22196\,
            in2 => \N__22641\,
            in3 => \N__19320\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__46047\,
            ce => \N__24812\,
            sr => \N__45569\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22485\,
            in2 => \N__20961\,
            in3 => \N__19317\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__46047\,
            ce => \N__24812\,
            sr => \N__45569\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22621\,
            in2 => \N__21045\,
            in3 => \N__19314\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__46047\,
            ce => \N__24812\,
            sr => \N__45569\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21674\,
            in2 => \N__22653\,
            in3 => \N__19311\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__46047\,
            ce => \N__24812\,
            sr => \N__45569\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20952\,
            in2 => \N__23985\,
            in3 => \N__19308\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__46047\,
            ce => \N__24812\,
            sr => \N__45569\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22787\,
            in2 => \N__21093\,
            in3 => \N__19305\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__46039\,
            ce => \N__24748\,
            sr => \N__45572\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21066\,
            in2 => \N__22374\,
            in3 => \N__19416\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__46039\,
            ce => \N__24748\,
            sr => \N__45572\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22416\,
            in2 => \N__21054\,
            in3 => \N__19413\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__46039\,
            ce => \N__24748\,
            sr => \N__45572\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22438\,
            in2 => \N__21027\,
            in3 => \N__19410\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__46039\,
            ce => \N__24748\,
            sr => \N__45572\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21060\,
            in2 => \N__23004\,
            in3 => \N__19407\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__46039\,
            ce => \N__24748\,
            sr => \N__45572\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23097\,
            in2 => \N__21018\,
            in3 => \N__19404\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__46039\,
            ce => \N__24748\,
            sr => \N__45572\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22521\,
            in2 => \N__21036\,
            in3 => \N__19401\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__46039\,
            ce => \N__24748\,
            sr => \N__45572\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21099\,
            in2 => \N__22893\,
            in3 => \N__19398\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__46039\,
            ce => \N__24748\,
            sr => \N__45572\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22068\,
            in2 => \N__20997\,
            in3 => \N__19395\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__46028\,
            ce => \N__24786\,
            sr => \N__45575\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21117\,
            in2 => \N__22242\,
            in3 => \N__19392\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__46028\,
            ce => \N__24786\,
            sr => \N__45575\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22571\,
            in2 => \N__21130\,
            in3 => \N__19629\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__46028\,
            ce => \N__24786\,
            sr => \N__45575\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21121\,
            in2 => \N__22692\,
            in3 => \N__19626\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__46028\,
            ce => \N__24786\,
            sr => \N__45575\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22958\,
            in2 => \N__21131\,
            in3 => \N__19623\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__46028\,
            ce => \N__24786\,
            sr => \N__45575\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21125\,
            in2 => \N__22833\,
            in3 => \N__19620\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__46028\,
            ce => \N__24786\,
            sr => \N__45575\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22145\,
            in2 => \N__21132\,
            in3 => \N__19617\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__46028\,
            ce => \N__24786\,
            sr => \N__45575\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23579\,
            in1 => \N__21129\,
            in2 => \_gnd_net_\,
            in3 => \N__19614\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46028\,
            ce => \N__24786\,
            sr => \N__45575\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19545\,
            in1 => \N__19848\,
            in2 => \N__19526\,
            in3 => \N__19811\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19866\,
            in1 => \N__19938\,
            in2 => \N__19506\,
            in3 => \N__19635\,
            lcout => \current_shift_inst.PI_CTRL.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__19445\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19427\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19970\,
            in1 => \N__19958\,
            in2 => \N__19941\,
            in3 => \N__19826\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19931\,
            in1 => \N__19913\,
            in2 => \N__19899\,
            in3 => \N__19881\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIFF4_21_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19736\,
            in1 => \N__19778\,
            in2 => \N__19721\,
            in3 => \N__19763\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1SC4_17_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19749\,
            in1 => \N__19847\,
            in2 => \N__19830\,
            in3 => \N__19812\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19779\,
            in2 => \_gnd_net_\,
            in3 => \N__19764\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19748\,
            in1 => \N__19737\,
            in2 => \N__19722\,
            in3 => \N__19701\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19683\,
            in1 => \N__19664\,
            in2 => \N__19644\,
            in3 => \N__19641\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_6_LC_3_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20019\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46074\,
            ce => 'H',
            sr => \N__45511\
        );

    \pwm_generator_inst.threshold_5_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20013\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46074\,
            ce => 'H',
            sr => \N__45511\
        );

    \pwm_generator_inst.threshold_7_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19995\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46074\,
            ce => 'H',
            sr => \N__45511\
        );

    \pwm_generator_inst.threshold_4_LC_3_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20007\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46074\,
            ce => 'H',
            sr => \N__45511\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_3_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__20422\,
            in1 => \N__20336\,
            in2 => \N__20274\,
            in3 => \N__20001\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46074\,
            ce => 'H',
            sr => \N__45511\
        );

    \pwm_generator_inst.threshold_0_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19989\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46074\,
            ce => 'H',
            sr => \N__45511\
        );

    \pwm_generator_inst.threshold_3_LC_3_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20430\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46074\,
            ce => 'H',
            sr => \N__45511\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__20338\,
            in1 => \N__19983\,
            in2 => \N__20423\,
            in3 => \N__20269\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46072\,
            ce => 'H',
            sr => \N__45519\
        );

    \pwm_generator_inst.threshold_1_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19977\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46072\,
            ce => 'H',
            sr => \N__45519\
        );

    \pwm_generator_inst.threshold_9_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20445\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46072\,
            ce => 'H',
            sr => \N__45519\
        );

    \pwm_generator_inst.threshold_8_LC_3_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20115\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46072\,
            ce => 'H',
            sr => \N__45519\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__20339\,
            in1 => \N__20270\,
            in2 => \N__20424\,
            in3 => \N__20436\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46072\,
            ce => 'H',
            sr => \N__45519\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__20410\,
            in1 => \N__20337\,
            in2 => \N__20280\,
            in3 => \N__20121\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46067\,
            ce => 'H',
            sr => \N__45527\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20097\,
            in2 => \_gnd_net_\,
            in3 => \N__20109\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20079\,
            in2 => \_gnd_net_\,
            in3 => \N__20091\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20061\,
            in2 => \_gnd_net_\,
            in3 => \N__20073\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20043\,
            in2 => \_gnd_net_\,
            in3 => \N__20055\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20025\,
            in2 => \_gnd_net_\,
            in3 => \N__20037\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20652\,
            in2 => \_gnd_net_\,
            in3 => \N__20664\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20634\,
            in2 => \_gnd_net_\,
            in3 => \N__20646\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20616\,
            in2 => \_gnd_net_\,
            in3 => \N__20628\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20598\,
            in2 => \_gnd_net_\,
            in3 => \N__20610\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_3_10_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20580\,
            in2 => \_gnd_net_\,
            in3 => \N__20592\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20572\,
            in2 => \_gnd_net_\,
            in3 => \N__20544\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__20534\,
            in1 => \N__20475\,
            in2 => \_gnd_net_\,
            in3 => \N__20448\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20869\,
            in2 => \_gnd_net_\,
            in3 => \N__20841\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20838\,
            in3 => \N__20805\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20800\,
            in2 => \_gnd_net_\,
            in3 => \N__20772\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20768\,
            in2 => \_gnd_net_\,
            in3 => \N__20751\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20746\,
            in2 => \_gnd_net_\,
            in3 => \N__20724\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_3_11_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20720\,
            in2 => \_gnd_net_\,
            in3 => \N__20703\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20699\,
            in2 => \_gnd_net_\,
            in3 => \N__20682\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20679\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22735\,
            in2 => \_gnd_net_\,
            in3 => \N__21505\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__22280\,
            in1 => \N__23052\,
            in2 => \N__20928\,
            in3 => \N__21467\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22736\,
            in1 => \N__22279\,
            in2 => \N__21468\,
            in3 => \N__21504\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__21589\,
            in1 => \N__23051\,
            in2 => \N__20925\,
            in3 => \N__21540\,
            lcout => \current_shift_inst.PI_CTRL.N_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__21376\,
            in1 => \N__21616\,
            in2 => \_gnd_net_\,
            in3 => \N__21421\,
            lcout => \current_shift_inst.PI_CTRL.un1_enablelt3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010001"
        )
    port map (
            in0 => \N__21541\,
            in1 => \N__21590\,
            in2 => \N__20922\,
            in3 => \N__20913\,
            lcout => \current_shift_inst.PI_CTRL.N_167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24029\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46048\,
            ce => \N__24822\,
            sr => \N__45561\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24008\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46048\,
            ce => \N__24822\,
            sr => \N__45561\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24050\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46048\,
            ce => \N__24822\,
            sr => \N__45561\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24362\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46048\,
            ce => \N__24822\,
            sr => \N__45561\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24338\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46048\,
            ce => \N__24822\,
            sr => \N__45561\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24095\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46048\,
            ce => \N__24822\,
            sr => \N__45561\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24221\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46040\,
            ce => \N__24770\,
            sr => \N__45566\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__21654\,
            in1 => \N__23900\,
            in2 => \N__23620\,
            in3 => \N__23758\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46040\,
            ce => \N__24770\,
            sr => \N__45566\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100000001"
        )
    port map (
            in0 => \N__23760\,
            in1 => \N__23603\,
            in2 => \N__23920\,
            in3 => \N__21441\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46040\,
            ce => \N__24770\,
            sr => \N__45566\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24549\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46040\,
            ce => \N__24770\,
            sr => \N__45566\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24290\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46040\,
            ce => \N__24770\,
            sr => \N__45566\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__21747\,
            in1 => \N__23901\,
            in2 => \N__23621\,
            in3 => \N__23759\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46040\,
            ce => \N__24770\,
            sr => \N__45566\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24314\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46040\,
            ce => \N__24770\,
            sr => \N__45566\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24497\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => \N__24716\,
            sr => \N__45570\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24431\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => \N__24716\,
            sr => \N__45570\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24476\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => \N__24716\,
            sr => \N__45570\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24198\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => \N__24716\,
            sr => \N__45570\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24383\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => \N__24716\,
            sr => \N__45570\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24452\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46029\,
            ce => \N__24716\,
            sr => \N__45570\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24408\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46018\,
            ce => \N__24766\,
            sr => \N__45573\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24267\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46018\,
            ce => \N__24766\,
            sr => \N__45573\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24941\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46018\,
            ce => \N__24766\,
            sr => \N__45573\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24915\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46018\,
            ce => \N__24766\,
            sr => \N__45573\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24971\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46018\,
            ce => \N__24766\,
            sr => \N__45573\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24527\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46010\,
            ce => \N__24703\,
            sr => \N__45576\
        );

    \un5_counter_cry_1_c_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22015\,
            in2 => \N__22038\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => un5_counter_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21795\,
            in2 => \_gnd_net_\,
            in3 => \N__21081\,
            lcout => \counterZ0Z_2\,
            ltout => OPEN,
            carryin => un5_counter_cry_1,
            carryout => un5_counter_cry_2,
            clk => \N__46001\,
            ce => 'H',
            sr => \N__45577\
        );

    \counter_3_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21783\,
            in2 => \_gnd_net_\,
            in3 => \N__21078\,
            lcout => \counterZ0Z_3\,
            ltout => OPEN,
            carryin => un5_counter_cry_2,
            carryout => un5_counter_cry_3,
            clk => \N__46001\,
            ce => 'H',
            sr => \N__45577\
        );

    \counter_4_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21770\,
            in2 => \_gnd_net_\,
            in3 => \N__21075\,
            lcout => \counterZ0Z_4\,
            ltout => OPEN,
            carryin => un5_counter_cry_3,
            carryout => un5_counter_cry_4,
            clk => \N__46001\,
            ce => 'H',
            sr => \N__45577\
        );

    \counter_5_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21995\,
            in1 => \N__21813\,
            in2 => \_gnd_net_\,
            in3 => \N__21072\,
            lcout => \counterZ0Z_5\,
            ltout => OPEN,
            carryin => un5_counter_cry_4,
            carryout => un5_counter_cry_5,
            clk => \N__46001\,
            ce => 'H',
            sr => \N__45577\
        );

    \counter_6_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21897\,
            in2 => \_gnd_net_\,
            in3 => \N__21069\,
            lcout => \counterZ0Z_6\,
            ltout => OPEN,
            carryin => un5_counter_cry_5,
            carryout => un5_counter_cry_6,
            clk => \N__46001\,
            ce => 'H',
            sr => \N__45577\
        );

    \counter_7_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21996\,
            in1 => \N__21843\,
            in2 => \_gnd_net_\,
            in3 => \N__21180\,
            lcout => \counterZ0Z_7\,
            ltout => OPEN,
            carryin => un5_counter_cry_6,
            carryout => un5_counter_cry_7,
            clk => \N__46001\,
            ce => 'H',
            sr => \N__45577\
        );

    \counter_8_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21986\,
            in1 => \N__21855\,
            in2 => \_gnd_net_\,
            in3 => \N__21177\,
            lcout => \counterZ0Z_8\,
            ltout => OPEN,
            carryin => un5_counter_cry_7,
            carryout => un5_counter_cry_8,
            clk => \N__46001\,
            ce => 'H',
            sr => \N__45577\
        );

    \counter_9_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21987\,
            in1 => \N__21827\,
            in2 => \_gnd_net_\,
            in3 => \N__21174\,
            lcout => \counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => un5_counter_cry_9,
            clk => \N__45993\,
            ce => 'H',
            sr => \N__45579\
        );

    \counter_10_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21870\,
            in2 => \_gnd_net_\,
            in3 => \N__21171\,
            lcout => \counterZ0Z_10\,
            ltout => OPEN,
            carryin => un5_counter_cry_9,
            carryout => un5_counter_cry_10,
            clk => \N__45993\,
            ce => 'H',
            sr => \N__45579\
        );

    \counter_11_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21911\,
            in2 => \_gnd_net_\,
            in3 => \N__21168\,
            lcout => \counterZ0Z_11\,
            ltout => OPEN,
            carryin => un5_counter_cry_10,
            carryout => un5_counter_cry_11,
            clk => \N__45993\,
            ce => 'H',
            sr => \N__45579\
        );

    \counter_12_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21994\,
            in1 => \N__21884\,
            in2 => \_gnd_net_\,
            in3 => \N__21165\,
            lcout => \counterZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45993\,
            ce => 'H',
            sr => \N__45579\
        );

    \clk_10khz_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21954\,
            in2 => \_gnd_net_\,
            in3 => \N__21988\,
            lcout => clk_10khz_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45993\,
            ce => 'H',
            sr => \N__45579\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21153\,
            in2 => \N__21162\,
            in3 => \N__23293\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_4_6_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21138\,
            in2 => \N__21147\,
            in3 => \N__23314\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21291\,
            in2 => \N__21303\,
            in3 => \N__23221\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21276\,
            in2 => \N__21285\,
            in3 => \N__23245\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23269\,
            in1 => \N__21261\,
            in2 => \N__21270\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21255\,
            in2 => \N__21249\,
            in3 => \N__23332\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21231\,
            in2 => \N__21240\,
            in3 => \N__23173\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23197\,
            in1 => \N__21216\,
            in2 => \N__21225\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21201\,
            in2 => \N__21210\,
            in3 => \N__23356\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_4_7_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21186\,
            in2 => \N__21195\,
            in3 => \N__23380\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21354\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46068\,
            ce => 'H',
            sr => \N__45512\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__21636\,
            in1 => \N__23862\,
            in2 => \N__23622\,
            in3 => \N__23757\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46064\,
            ce => \N__24823\,
            sr => \N__45520\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__21561\,
            in1 => \N__23794\,
            in2 => \_gnd_net_\,
            in3 => \N__23747\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46059\,
            ce => \N__24775\,
            sr => \N__45535\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22911\,
            in1 => \N__21330\,
            in2 => \N__22077\,
            in3 => \N__21309\,
            lcout => \current_shift_inst.PI_CTRL.N_170\,
            ltout => \current_shift_inst.PI_CTRL.N_170_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111011001010"
        )
    port map (
            in0 => \N__23588\,
            in1 => \N__21723\,
            in2 => \N__21336\,
            in3 => \N__23746\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46059\,
            ce => \N__24775\,
            sr => \N__45535\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22408\,
            in1 => \N__22446\,
            in2 => \N__22366\,
            in3 => \N__22516\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGGAM_21_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22570\,
            in1 => \N__22230\,
            in2 => \N__22959\,
            in3 => \N__23096\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIONJC1_12_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21680\,
            in1 => \N__22473\,
            in2 => \N__21333\,
            in3 => \N__21432\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIQV7U3_20_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21324\,
            in1 => \N__22063\,
            in2 => \N__21318\,
            in3 => \N__23003\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22788\,
            in1 => \N__22622\,
            in2 => \N__22197\,
            in3 => \N__21681\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI676B_27_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22680\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23688\,
            in1 => \N__23589\,
            in2 => \N__23898\,
            in3 => \N__21522\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46049\,
            ce => \N__24774\,
            sr => \N__45550\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__21360\,
            in1 => \N__23844\,
            in2 => \_gnd_net_\,
            in3 => \N__23686\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46049\,
            ce => \N__24774\,
            sr => \N__45550\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__23687\,
            in1 => \_gnd_net_\,
            in2 => \N__23897\,
            in3 => \N__21600\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46049\,
            ce => \N__24774\,
            sr => \N__45550\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__21696\,
            in1 => \N__23843\,
            in2 => \N__23617\,
            in3 => \N__23685\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46049\,
            ce => \N__24774\,
            sr => \N__45550\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001011001000"
        )
    port map (
            in0 => \N__23690\,
            in1 => \N__24132\,
            in2 => \N__23899\,
            in3 => \N__21422\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46049\,
            ce => \N__24774\,
            sr => \N__45550\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101010001011"
        )
    port map (
            in0 => \N__21486\,
            in1 => \N__23851\,
            in2 => \N__23618\,
            in3 => \N__23689\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46049\,
            ce => \N__24774\,
            sr => \N__45550\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21417\,
            in2 => \N__24131\,
            in3 => \N__24127\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\,
            clk => \N__46041\,
            ce => \N__24821\,
            sr => \N__45556\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21377\,
            in2 => \N__24096\,
            in3 => \N__21627\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21617\,
            in2 => \N__24072\,
            in3 => \N__21594\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21585\,
            in2 => \N__24051\,
            in3 => \N__21552\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21542\,
            in2 => \N__24030\,
            in3 => \N__21516\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21506\,
            in2 => \N__24009\,
            in3 => \N__21480\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22278\,
            in2 => \N__24363\,
            in3 => \N__21477\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22717\,
            in2 => \N__24339\,
            in3 => \N__21474\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23041\,
            in2 => \N__24315\,
            in3 => \N__21471\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21462\,
            in2 => \N__24291\,
            in3 => \N__21435\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22851\,
            in2 => \N__24266\,
            in3 => \N__21702\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24242\,
            in2 => \N__22188\,
            in3 => \N__21699\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22480\,
            in2 => \N__24222\,
            in3 => \N__21687\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22614\,
            in2 => \N__24197\,
            in3 => \N__21684\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21670\,
            in2 => \N__24174\,
            in3 => \N__21648\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24548\,
            in2 => \N__23973\,
            in3 => \N__21645\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22773\,
            in2 => \N__24528\,
            in3 => \N__21642\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22370\,
            in2 => \N__24498\,
            in3 => \N__21639\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22415\,
            in2 => \N__24477\,
            in3 => \N__21750\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22437\,
            in2 => \N__24453\,
            in3 => \N__21738\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22992\,
            in2 => \N__24432\,
            in3 => \N__21735\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23088\,
            in2 => \N__24407\,
            in3 => \N__21732\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22509\,
            in2 => \N__24384\,
            in3 => \N__21729\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22886\,
            in2 => \N__24972\,
            in3 => \N__21726\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22064\,
            in2 => \N__24942\,
            in3 => \N__21711\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22238\,
            in2 => \N__24916\,
            in3 => \N__21708\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24905\,
            in2 => \N__22572\,
            in3 => \N__21705\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22688\,
            in2 => \N__24917\,
            in3 => \N__21927\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24909\,
            in2 => \N__22957\,
            in3 => \N__21924\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22821\,
            in2 => \N__24918\,
            in3 => \N__21921\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24913\,
            in2 => \N__22146\,
            in3 => \N__21918\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__24914\,
            in1 => \_gnd_net_\,
            in2 => \N__23557\,
            in3 => \N__21915\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un2_counter_1_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21912\,
            in1 => \N__21896\,
            in2 => \N__21885\,
            in3 => \N__22014\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un2_counterZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un2_counter_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21869\,
            in1 => \N__21801\,
            in2 => \N__21858\,
            in3 => \N__21756\,
            lcout => \current_shift_inst.PI_CTRL.un2_counterZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un2_counter_8_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21854\,
            in1 => \N__21842\,
            in2 => \N__21831\,
            in3 => \N__21812\,
            lcout => \current_shift_inst.PI_CTRL.un2_counterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un2_counter_7_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21794\,
            in1 => \N__21782\,
            in2 => \N__21771\,
            in3 => \N__22033\,
            lcout => \current_shift_inst.PI_CTRL.un2_counterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22017\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22037\,
            lcout => \counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45982\,
            ce => 'H',
            sr => \N__45578\
        );

    \counter_0_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21985\,
            in2 => \_gnd_net_\,
            in3 => \N__22016\,
            lcout => \counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45982\,
            ce => 'H',
            sr => \N__45578\
        );

    \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__29392\,
            in1 => \N__21984\,
            in2 => \_gnd_net_\,
            in3 => \N__21953\,
            lcout => \N_748_g\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23152\,
            in1 => \N__23294\,
            in2 => \_gnd_net_\,
            in3 => \N__21942\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__46069\,
            ce => 'H',
            sr => \N__45494\
        );

    \pwm_generator_inst.counter_1_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23148\,
            in1 => \N__23315\,
            in2 => \_gnd_net_\,
            in3 => \N__21939\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__46069\,
            ce => 'H',
            sr => \N__45494\
        );

    \pwm_generator_inst.counter_2_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23153\,
            in1 => \N__23229\,
            in2 => \_gnd_net_\,
            in3 => \N__21936\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__46069\,
            ce => 'H',
            sr => \N__45494\
        );

    \pwm_generator_inst.counter_3_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23149\,
            in1 => \N__23253\,
            in2 => \_gnd_net_\,
            in3 => \N__21933\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__46069\,
            ce => 'H',
            sr => \N__45494\
        );

    \pwm_generator_inst.counter_4_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23154\,
            in1 => \N__23273\,
            in2 => \_gnd_net_\,
            in3 => \N__21930\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__46069\,
            ce => 'H',
            sr => \N__45494\
        );

    \pwm_generator_inst.counter_5_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23150\,
            in1 => \N__23336\,
            in2 => \_gnd_net_\,
            in3 => \N__22104\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__46069\,
            ce => 'H',
            sr => \N__45494\
        );

    \pwm_generator_inst.counter_6_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23155\,
            in1 => \N__23174\,
            in2 => \_gnd_net_\,
            in3 => \N__22101\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__46069\,
            ce => 'H',
            sr => \N__45494\
        );

    \pwm_generator_inst.counter_7_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23151\,
            in1 => \N__23201\,
            in2 => \_gnd_net_\,
            in3 => \N__22098\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__46069\,
            ce => 'H',
            sr => \N__45494\
        );

    \pwm_generator_inst.counter_8_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23157\,
            in1 => \N__23357\,
            in2 => \_gnd_net_\,
            in3 => \N__22095\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__46065\,
            ce => 'H',
            sr => \N__45502\
        );

    \pwm_generator_inst.counter_9_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23156\,
            in1 => \N__23381\,
            in2 => \_gnd_net_\,
            in3 => \N__22092\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46065\,
            ce => 'H',
            sr => \N__45502\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__22089\,
            in1 => \N__23795\,
            in2 => \N__23619\,
            in3 => \N__23745\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46056\,
            ce => \N__24871\,
            sr => \N__45528\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI736M_11_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22192\,
            in1 => \N__23978\,
            in2 => \N__22623\,
            in3 => \N__22783\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI225B_20_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22056\,
            in2 => \_gnd_net_\,
            in3 => \N__22996\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22231\,
            in1 => \N__22138\,
            in2 => \N__22956\,
            in3 => \N__22681\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICB2E2_12_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__23525\,
            in1 => \N__22481\,
            in2 => \N__22449\,
            in3 => \N__22323\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22445\,
            in1 => \N__22407\,
            in2 => \N__22520\,
            in3 => \N__22356\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIQNHC1_21_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__22557\,
            in1 => \N__23095\,
            in2 => \N__22332\,
            in3 => \N__22329\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIC35V7_10_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22317\,
            in1 => \N__22308\,
            in2 => \N__23943\,
            in3 => \N__22299\,
            lcout => \current_shift_inst.PI_CTRL.N_171\,
            ltout => \current_shift_inst.PI_CTRL.N_171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001000101"
        )
    port map (
            in0 => \N__23542\,
            in1 => \N__22293\,
            in2 => \N__22287\,
            in3 => \N__23863\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46042\,
            ce => \N__24857\,
            sr => \N__45542\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23681\,
            in1 => \N__23544\,
            in2 => \N__22257\,
            in3 => \N__23869\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46030\,
            ce => \N__24785\,
            sr => \N__45551\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__22203\,
            in1 => \N__23864\,
            in2 => \N__23599\,
            in3 => \N__23678\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46030\,
            ce => \N__24785\,
            sr => \N__45551\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__22158\,
            in1 => \N__23867\,
            in2 => \N__23602\,
            in3 => \N__23683\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46030\,
            ce => \N__24785\,
            sr => \N__45551\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23680\,
            in1 => \N__23543\,
            in2 => \N__22800\,
            in3 => \N__23868\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46030\,
            ce => \N__24785\,
            sr => \N__45551\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__22752\,
            in1 => \N__23865\,
            in2 => \N__23600\,
            in3 => \N__23679\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46030\,
            ce => \N__24785\,
            sr => \N__45551\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000001101"
        )
    port map (
            in0 => \N__23684\,
            in1 => \N__22746\,
            in2 => \N__23613\,
            in3 => \N__23870\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46030\,
            ce => \N__24785\,
            sr => \N__45551\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__22701\,
            in1 => \N__23866\,
            in2 => \N__23601\,
            in3 => \N__23682\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46030\,
            ce => \N__24785\,
            sr => \N__45551\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24173\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46019\,
            ce => \N__24856\,
            sr => \N__45557\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24243\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46019\,
            ce => \N__24856\,
            sr => \N__45557\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__22629\,
            in1 => \N__23905\,
            in2 => \N__23610\,
            in3 => \N__23728\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46019\,
            ce => \N__24856\,
            sr => \N__45557\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23731\,
            in1 => \N__23565\,
            in2 => \N__23921\,
            in3 => \N__22584\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46019\,
            ce => \N__24856\,
            sr => \N__45557\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__22527\,
            in1 => \N__23907\,
            in2 => \N__23612\,
            in3 => \N__23730\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46019\,
            ce => \N__24856\,
            sr => \N__45557\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__23103\,
            in1 => \N__23906\,
            in2 => \N__23611\,
            in3 => \N__23729\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46019\,
            ce => \N__24856\,
            sr => \N__45557\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100000001"
        )
    port map (
            in0 => \N__23732\,
            in1 => \N__23566\,
            in2 => \N__23922\,
            in3 => \N__23061\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46019\,
            ce => \N__24856\,
            sr => \N__45557\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__23022\,
            in1 => \N__23914\,
            in2 => \N__23580\,
            in3 => \N__23733\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46011\,
            ce => \N__24826\,
            sr => \N__45562\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__23016\,
            in1 => \N__23916\,
            in2 => \N__23582\,
            in3 => \N__23735\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46011\,
            ce => \N__24826\,
            sr => \N__45562\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__23010\,
            in1 => \N__23915\,
            in2 => \N__23581\,
            in3 => \N__23734\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46011\,
            ce => \N__24826\,
            sr => \N__45562\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23736\,
            in1 => \N__23508\,
            in2 => \N__22968\,
            in3 => \N__23917\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46011\,
            ce => \N__24826\,
            sr => \N__45562\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI99AM_10_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22822\,
            in1 => \N__22852\,
            in2 => \N__23524\,
            in3 => \N__22885\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__22899\,
            in1 => \N__23918\,
            in2 => \N__23583\,
            in3 => \N__23755\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46002\,
            ce => \N__24732\,
            sr => \N__45567\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22884\,
            in1 => \N__22853\,
            in2 => \N__22829\,
            in3 => \N__23974\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__23928\,
            in1 => \N__23919\,
            in2 => \N__23584\,
            in3 => \N__23756\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46002\,
            ce => \N__24732\,
            sr => \N__45567\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23397\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNITBL3_9_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23385\,
            in1 => \N__23361\,
            in2 => \_gnd_net_\,
            in3 => \N__23337\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIRPD2_0_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23316\,
            in2 => \_gnd_net_\,
            in3 => \N__23295\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__23274\,
            in1 => \N__23252\,
            in2 => \N__23232\,
            in3 => \N__23228\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_6_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23208\,
            in1 => \N__23202\,
            in2 => \N__23181\,
            in3 => \N__23178\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__29038\,
            in1 => \N__28822\,
            in2 => \N__25104\,
            in3 => \N__28964\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46031\,
            ce => 'H',
            sr => \N__45521\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__29037\,
            in1 => \N__28821\,
            in2 => \_gnd_net_\,
            in3 => \N__28963\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__25016\,
            in1 => \N__29193\,
            in2 => \N__24153\,
            in3 => \N__29158\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46031\,
            ce => 'H',
            sr => \N__45521\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24068\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46020\,
            ce => \N__24846\,
            sr => \N__45529\
        );

    \current_shift_inst.control_input_0_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25185\,
            in2 => \N__26970\,
            in3 => \N__26969\,
            lcout => \current_shift_inst.control_inputZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \current_shift_inst.control_input_1_cry_0\,
            clk => \N__46012\,
            ce => \N__24825\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25260\,
            in2 => \_gnd_net_\,
            in3 => \N__24075\,
            lcout => \current_shift_inst.control_inputZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_0\,
            carryout => \current_shift_inst.control_input_1_cry_1\,
            clk => \N__46012\,
            ce => \N__24825\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25155\,
            in2 => \_gnd_net_\,
            in3 => \N__24054\,
            lcout => \current_shift_inst.control_inputZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_1\,
            carryout => \current_shift_inst.control_input_1_cry_2\,
            clk => \N__46012\,
            ce => \N__24825\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25173\,
            in2 => \_gnd_net_\,
            in3 => \N__24033\,
            lcout => \current_shift_inst.control_inputZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_2\,
            carryout => \current_shift_inst.control_input_1_cry_3\,
            clk => \N__46012\,
            ce => \N__24825\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_4_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25239\,
            in2 => \_gnd_net_\,
            in3 => \N__24012\,
            lcout => \current_shift_inst.control_inputZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_3\,
            carryout => \current_shift_inst.control_input_1_cry_4\,
            clk => \N__46012\,
            ce => \N__24825\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_5_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25143\,
            in2 => \_gnd_net_\,
            in3 => \N__23988\,
            lcout => \current_shift_inst.control_inputZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_4\,
            carryout => \current_shift_inst.control_input_1_cry_5\,
            clk => \N__46012\,
            ce => \N__24825\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_6_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25149\,
            in2 => \_gnd_net_\,
            in3 => \N__24342\,
            lcout => \current_shift_inst.control_inputZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_5\,
            carryout => \current_shift_inst.control_input_1_cry_6\,
            clk => \N__46012\,
            ce => \N__24825\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_7_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25227\,
            in2 => \_gnd_net_\,
            in3 => \N__24318\,
            lcout => \current_shift_inst.control_inputZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_6\,
            carryout => \current_shift_inst.control_input_1_cry_7\,
            clk => \N__46012\,
            ce => \N__24825\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_8_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25200\,
            in2 => \_gnd_net_\,
            in3 => \N__24294\,
            lcout => \current_shift_inst.control_inputZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \current_shift_inst.control_input_1_cry_8\,
            clk => \N__46003\,
            ce => \N__24845\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_9_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25272\,
            in2 => \_gnd_net_\,
            in3 => \N__24270\,
            lcout => \current_shift_inst.control_inputZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_8\,
            carryout => \current_shift_inst.control_input_1_cry_9\,
            clk => \N__46003\,
            ce => \N__24845\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_10_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25113\,
            in2 => \_gnd_net_\,
            in3 => \N__24246\,
            lcout => \current_shift_inst.control_inputZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_9\,
            carryout => \current_shift_inst.control_input_1_cry_10\,
            clk => \N__46003\,
            ce => \N__24845\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_11_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25209\,
            in3 => \N__24225\,
            lcout => \current_shift_inst.control_inputZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_10\,
            carryout => \current_shift_inst.control_input_1_cry_11\,
            clk => \N__46003\,
            ce => \N__24845\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_12_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25125\,
            in2 => \_gnd_net_\,
            in3 => \N__24201\,
            lcout => \current_shift_inst.control_inputZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_11\,
            carryout => \current_shift_inst.control_input_1_cry_12\,
            clk => \N__46003\,
            ce => \N__24845\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_13_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25131\,
            in2 => \_gnd_net_\,
            in3 => \N__24177\,
            lcout => \current_shift_inst.control_inputZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_12\,
            carryout => \current_shift_inst.control_input_1_cry_13\,
            clk => \N__46003\,
            ce => \N__24845\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_14_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25137\,
            in2 => \_gnd_net_\,
            in3 => \N__24156\,
            lcout => \current_shift_inst.control_inputZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_13\,
            carryout => \current_shift_inst.control_input_1_cry_14\,
            clk => \N__46003\,
            ce => \N__24845\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_15_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25119\,
            in2 => \_gnd_net_\,
            in3 => \N__24531\,
            lcout => \current_shift_inst.control_inputZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_14\,
            carryout => \current_shift_inst.control_input_1_cry_15\,
            clk => \N__46003\,
            ce => \N__24845\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_16_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25215\,
            in2 => \_gnd_net_\,
            in3 => \N__24501\,
            lcout => \current_shift_inst.control_inputZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \current_shift_inst.control_input_1_cry_16\,
            clk => \N__45994\,
            ce => \N__24861\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_17_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25248\,
            in2 => \_gnd_net_\,
            in3 => \N__24480\,
            lcout => \current_shift_inst.control_inputZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_16\,
            carryout => \current_shift_inst.control_input_1_cry_17\,
            clk => \N__45994\,
            ce => \N__24861\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_18_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25296\,
            in2 => \_gnd_net_\,
            in3 => \N__24456\,
            lcout => \current_shift_inst.control_inputZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_17\,
            carryout => \current_shift_inst.control_input_1_cry_18\,
            clk => \N__45994\,
            ce => \N__24861\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_19_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25287\,
            in2 => \_gnd_net_\,
            in3 => \N__24435\,
            lcout => \current_shift_inst.control_inputZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_18\,
            carryout => \current_shift_inst.control_input_1_cry_19\,
            clk => \N__45994\,
            ce => \N__24861\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_20_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25194\,
            in2 => \_gnd_net_\,
            in3 => \N__24411\,
            lcout => \current_shift_inst.control_inputZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_19\,
            carryout => \current_shift_inst.control_input_1_cry_20\,
            clk => \N__45994\,
            ce => \N__24861\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_21_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25059\,
            in2 => \_gnd_net_\,
            in3 => \N__24387\,
            lcout => \current_shift_inst.control_inputZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_20\,
            carryout => \current_shift_inst.control_input_1_cry_21\,
            clk => \N__45994\,
            ce => \N__24861\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_22_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25065\,
            in2 => \_gnd_net_\,
            in3 => \N__24366\,
            lcout => \current_shift_inst.control_inputZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_21\,
            carryout => \current_shift_inst.control_input_1_cry_22\,
            clk => \N__45994\,
            ce => \N__24861\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_23_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24585\,
            in2 => \_gnd_net_\,
            in3 => \N__24945\,
            lcout => \current_shift_inst.control_inputZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_22\,
            carryout => \current_shift_inst.control_input_1_cry_23\,
            clk => \N__45994\,
            ce => \N__24861\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_24_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25278\,
            in2 => \_gnd_net_\,
            in3 => \N__24924\,
            lcout => \current_shift_inst.control_inputZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \current_shift_inst.control_input_1_cry_24\,
            clk => \N__45983\,
            ce => \N__24805\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_25_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25626\,
            in2 => \_gnd_net_\,
            in3 => \N__24921\,
            lcout => \current_shift_inst.control_inputZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45983\,
            ce => \N__24805\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_4_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29383\,
            in2 => \_gnd_net_\,
            in3 => \N__38186\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45976\,
            ce => 'H',
            sr => \N__45563\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29814\,
            in1 => \N__32292\,
            in2 => \N__30333\,
            in3 => \N__27807\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29802\,
            in1 => \N__32526\,
            in2 => \N__30334\,
            in3 => \N__27897\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__25650\,
            in1 => \N__26187\,
            in2 => \_gnd_net_\,
            in3 => \N__27092\,
            lcout => \current_shift_inst.control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24573\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24564\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46057\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25026\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46043\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25017\,
            in2 => \_gnd_net_\,
            in3 => \N__24995\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__27497\,
            in1 => \N__29059\,
            in2 => \N__25167\,
            in3 => \N__38213\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46032\,
            ce => 'H',
            sr => \N__45503\
        );

    \phase_controller_inst2.state_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__31792\,
            in1 => \N__25015\,
            in2 => \N__31739\,
            in3 => \N__24996\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46032\,
            ce => 'H',
            sr => \N__45503\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25074\,
            in2 => \N__26316\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26289\,
            in2 => \_gnd_net_\,
            in3 => \N__24984\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25083\,
            in2 => \N__26271\,
            in3 => \N__24981\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26250\,
            in2 => \_gnd_net_\,
            in3 => \N__24978\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26499\,
            in3 => \N__24975\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26478\,
            in2 => \_gnd_net_\,
            in3 => \N__25053\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26460\,
            in2 => \_gnd_net_\,
            in3 => \N__25050\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26433\,
            in2 => \_gnd_net_\,
            in3 => \N__25047\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26403\,
            in2 => \_gnd_net_\,
            in3 => \N__25044\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26385\,
            in2 => \_gnd_net_\,
            in3 => \N__25041\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26352\,
            in2 => \_gnd_net_\,
            in3 => \N__25038\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26334\,
            in2 => \_gnd_net_\,
            in3 => \N__25035\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26655\,
            in2 => \_gnd_net_\,
            in3 => \N__25032\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26637\,
            in2 => \_gnd_net_\,
            in3 => \N__25029\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26619\,
            in2 => \_gnd_net_\,
            in3 => \N__25107\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26585\,
            in2 => \_gnd_net_\,
            in3 => \N__25095\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26565\,
            in2 => \_gnd_net_\,
            in3 => \N__25092\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26547\,
            in2 => \_gnd_net_\,
            in3 => \N__25089\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26529\,
            in2 => \_gnd_net_\,
            in3 => \N__25086\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29148\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29181\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29147\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__27083\,
            in1 => \N__26202\,
            in2 => \_gnd_net_\,
            in3 => \N__25668\,
            lcout => \current_shift_inst.control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__25680\,
            in1 => \N__26217\,
            in2 => \_gnd_net_\,
            in3 => \N__27082\,
            lcout => \current_shift_inst.control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__25992\,
            in1 => \N__25455\,
            in2 => \_gnd_net_\,
            in3 => \N__27079\,
            lcout => \current_shift_inst.control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31722\,
            in2 => \_gnd_net_\,
            in3 => \N__31793\,
            lcout => \phase_controller_inst2.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__25311\,
            in1 => \N__25851\,
            in2 => \_gnd_net_\,
            in3 => \N__27078\,
            lcout => \current_shift_inst.control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__27081\,
            in1 => \N__25950\,
            in2 => \_gnd_net_\,
            in3 => \N__25419\,
            lcout => \current_shift_inst.control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__25965\,
            in1 => \N__25431\,
            in2 => \_gnd_net_\,
            in3 => \N__27080\,
            lcout => \current_shift_inst.control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__27089\,
            in1 => \N__25539\,
            in2 => \_gnd_net_\,
            in3 => \N__26091\,
            lcout => \current_shift_inst.control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__26109\,
            in1 => \N__25551\,
            in2 => \_gnd_net_\,
            in3 => \N__27088\,
            lcout => \current_shift_inst.control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__27087\,
            in1 => \N__26124\,
            in2 => \_gnd_net_\,
            in3 => \N__25566\,
            lcout => \current_shift_inst.control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__25527\,
            in1 => \N__26076\,
            in2 => \_gnd_net_\,
            in3 => \N__27090\,
            lcout => \current_shift_inst.control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__27085\,
            in1 => \N__25368\,
            in2 => \_gnd_net_\,
            in3 => \N__25890\,
            lcout => \current_shift_inst.control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__25512\,
            in1 => \N__26061\,
            in2 => \_gnd_net_\,
            in3 => \N__27091\,
            lcout => \current_shift_inst.control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__27086\,
            in1 => \N__26139\,
            in2 => \_gnd_net_\,
            in3 => \N__25587\,
            lcout => \current_shift_inst.control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__25395\,
            in1 => \N__25923\,
            in2 => \_gnd_net_\,
            in3 => \N__27084\,
            lcout => \current_shift_inst.control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32511\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29591\,
            in1 => \N__31566\,
            in2 => \N__30493\,
            in3 => \N__30729\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__26232\,
            in1 => \N__25704\,
            in2 => \_gnd_net_\,
            in3 => \N__27077\,
            lcout => \current_shift_inst.control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__32484\,
            in1 => \N__30332\,
            in2 => \N__29696\,
            in3 => \N__27867\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__25875\,
            in1 => \N__25338\,
            in2 => \_gnd_net_\,
            in3 => \N__27018\,
            lcout => \current_shift_inst.control_input_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29801\,
            in1 => \N__32757\,
            in2 => \N__30492\,
            in3 => \N__27978\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__27020\,
            in1 => \N__26031\,
            in2 => \_gnd_net_\,
            in3 => \N__25482\,
            lcout => \current_shift_inst.control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__26016\,
            in1 => \N__25467\,
            in2 => \_gnd_net_\,
            in3 => \N__27021\,
            lcout => \current_shift_inst.control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__27022\,
            in1 => \N__25641\,
            in2 => \_gnd_net_\,
            in3 => \N__26175\,
            lcout => \current_shift_inst.control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__25380\,
            in1 => \N__25905\,
            in2 => \_gnd_net_\,
            in3 => \N__27019\,
            lcout => \current_shift_inst.control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__25860\,
            in1 => \N__25320\,
            in2 => \_gnd_net_\,
            in3 => \N__27023\,
            lcout => \current_shift_inst.control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__27026\,
            in1 => \N__25494\,
            in2 => \_gnd_net_\,
            in3 => \N__26046\,
            lcout => \current_shift_inst.control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__25443\,
            in1 => \N__25977\,
            in2 => \_gnd_net_\,
            in3 => \N__27024\,
            lcout => \current_shift_inst.control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__27025\,
            in1 => \N__25935\,
            in2 => \_gnd_net_\,
            in3 => \N__25407\,
            lcout => \current_shift_inst.control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__29692\,
            in1 => \N__27633\,
            in2 => \N__26762\,
            in3 => \N__26703\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27528\,
            in2 => \N__34179\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25353\,
            in2 => \N__26755\,
            in3 => \N__34618\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34619\,
            in1 => \N__29235\,
            in2 => \N__30348\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30145\,
            in2 => \N__26943\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28413\,
            in2 => \N__30349\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25347\,
            in2 => \N__30272\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26835\,
            in2 => \N__30350\,
            in3 => \N__25329\,
            lcout => \current_shift_inst.un38_control_input_0_s0_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25326\,
            in2 => \N__30273\,
            in3 => \N__25314\,
            lcout => \current_shift_inst.un38_control_input_0_s0_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27249\,
            in2 => \N__30278\,
            in3 => \N__25299\,
            lcout => \current_shift_inst.un38_control_input_0_s0_8\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26871\,
            in2 => \N__30282\,
            in3 => \N__25446\,
            lcout => \current_shift_inst.un38_control_input_0_s0_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28350\,
            in2 => \N__30279\,
            in3 => \N__25434\,
            lcout => \current_shift_inst.un38_control_input_0_s0_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28317\,
            in2 => \N__30283\,
            in3 => \N__25422\,
            lcout => \current_shift_inst.un38_control_input_0_s0_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26910\,
            in2 => \N__30280\,
            in3 => \N__25410\,
            lcout => \current_shift_inst.un38_control_input_0_s0_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27240\,
            in2 => \N__30284\,
            in3 => \N__25398\,
            lcout => \current_shift_inst.un38_control_input_0_s0_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28281\,
            in2 => \N__30281\,
            in3 => \N__25383\,
            lcout => \current_shift_inst.un38_control_input_0_s0_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28245\,
            in2 => \N__30285\,
            in3 => \N__25371\,
            lcout => \current_shift_inst.un38_control_input_0_s0_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28566\,
            in2 => \N__30464\,
            in3 => \N__25356\,
            lcout => \current_shift_inst.un38_control_input_0_s0_16\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25593\,
            in2 => \N__30438\,
            in3 => \N__25578\,
            lcout => \current_shift_inst.un38_control_input_0_s0_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25575\,
            in2 => \N__30465\,
            in3 => \N__25554\,
            lcout => \current_shift_inst.un38_control_input_0_s0_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28062\,
            in2 => \N__30439\,
            in3 => \N__25542\,
            lcout => \current_shift_inst.un38_control_input_0_s0_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28098\,
            in2 => \N__30466\,
            in3 => \N__25530\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28449\,
            in2 => \N__30440\,
            in3 => \N__25515\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27306\,
            in2 => \N__30467\,
            in3 => \N__25497\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28026\,
            in2 => \N__30441\,
            in3 => \N__25485\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28188\,
            in2 => \N__30595\,
            in3 => \N__25470\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30448\,
            in2 => \N__27213\,
            in3 => \N__25707\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28158\,
            in2 => \N__30596\,
            in3 => \N__25692\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25689\,
            in2 => \N__30468\,
            in3 => \N__25671\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28386\,
            in2 => \N__30597\,
            in3 => \N__25653\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27297\,
            in2 => \N__30469\,
            in3 => \N__25644\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28545\,
            in2 => \N__30598\,
            in3 => \N__25632\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_0_25_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101101000111"
        )
    port map (
            in0 => \N__27681\,
            in1 => \N__27093\,
            in2 => \N__26157\,
            in3 => \N__25629\,
            lcout => \current_shift_inst.control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_8_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31743\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45930\,
            ce => 'H',
            sr => \N__45581\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25602\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25761\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__28824\,
            in1 => \N__28944\,
            in2 => \N__29084\,
            in3 => \N__25749\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46021\,
            ce => 'H',
            sr => \N__45495\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__28942\,
            in1 => \N__29039\,
            in2 => \N__25743\,
            in3 => \N__28825\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46021\,
            ce => 'H',
            sr => \N__45495\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__28823\,
            in1 => \N__28943\,
            in2 => \N__29083\,
            in3 => \N__25734\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46021\,
            ce => 'H',
            sr => \N__45495\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__28814\,
            in1 => \N__28935\,
            in2 => \N__29085\,
            in3 => \N__25728\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46013\,
            ce => 'H',
            sr => \N__45504\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29189\,
            in1 => \N__26315\,
            in2 => \_gnd_net_\,
            in3 => \N__29152\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__28817\,
            in1 => \N__29058\,
            in2 => \N__25722\,
            in3 => \N__28941\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46013\,
            ce => 'H',
            sr => \N__45504\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__25719\,
            in1 => \N__29046\,
            in2 => \N__28965\,
            in3 => \N__28820\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46013\,
            ce => 'H',
            sr => \N__45504\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__28815\,
            in1 => \N__28936\,
            in2 => \N__29086\,
            in3 => \N__25713\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46013\,
            ce => 'H',
            sr => \N__45504\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__28933\,
            in1 => \N__29047\,
            in2 => \N__25821\,
            in3 => \N__28818\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46013\,
            ce => 'H',
            sr => \N__45504\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__28816\,
            in1 => \N__28937\,
            in2 => \N__29087\,
            in3 => \N__25812\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46013\,
            ce => 'H',
            sr => \N__45504\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__28934\,
            in1 => \N__29048\,
            in2 => \N__25806\,
            in3 => \N__28819\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46013\,
            ce => 'H',
            sr => \N__45504\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__28826\,
            in1 => \N__29099\,
            in2 => \N__28978\,
            in3 => \N__25797\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46004\,
            ce => 'H',
            sr => \N__45513\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__28945\,
            in1 => \N__28830\,
            in2 => \N__29110\,
            in3 => \N__25791\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46004\,
            ce => 'H',
            sr => \N__45513\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__28827\,
            in1 => \N__29100\,
            in2 => \N__28979\,
            in3 => \N__25785\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46004\,
            ce => 'H',
            sr => \N__45513\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__25779\,
            in1 => \N__28831\,
            in2 => \N__28967\,
            in3 => \N__29094\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46004\,
            ce => 'H',
            sr => \N__45513\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010001010"
        )
    port map (
            in0 => \N__25773\,
            in1 => \N__28946\,
            in2 => \N__28836\,
            in3 => \N__29101\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46004\,
            ce => 'H',
            sr => \N__45513\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011000100"
        )
    port map (
            in0 => \N__29103\,
            in1 => \N__25767\,
            in2 => \N__28968\,
            in3 => \N__28832\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46004\,
            ce => 'H',
            sr => \N__45513\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__28828\,
            in1 => \N__29102\,
            in2 => \N__28980\,
            in3 => \N__25833\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46004\,
            ce => 'H',
            sr => \N__45513\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__29098\,
            in1 => \N__28829\,
            in2 => \N__28966\,
            in3 => \N__25827\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46004\,
            ce => 'H',
            sr => \N__45513\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29579\,
            in1 => \N__32204\,
            in2 => \N__30672\,
            in3 => \N__27771\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32994\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45995\,
            ce => \N__32967\,
            sr => \N__45522\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33666\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45984\,
            ce => \N__32966\,
            sr => \N__45530\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34652\,
            in2 => \N__34623\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26679\,
            in2 => \N__34580\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26673\,
            in2 => \N__34588\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26847\,
            in2 => \N__34581\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26811\,
            in2 => \N__34589\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26859\,
            in2 => \N__34582\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26775\,
            in2 => \N__34590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26709\,
            in2 => \N__34583\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26841\,
            in2 => \N__34579\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26817\,
            in2 => \N__34587\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26928\,
            in2 => \N__34576\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26853\,
            in2 => \N__34584\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26823\,
            in2 => \N__34577\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26922\,
            in2 => \N__34585\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26898\,
            in2 => \N__34578\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26916\,
            in2 => \N__34586\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26877\,
            in2 => \N__34567\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26892\,
            in2 => \N__34571\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27135\,
            in2 => \N__34568\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34490\,
            in2 => \N__26886\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27129\,
            in2 => \N__34569\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30807\,
            in2 => \N__34572\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27123\,
            in2 => \N__34570\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27117\,
            in2 => \N__34573\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34375\,
            in2 => \N__27144\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27111\,
            in2 => \N__34478\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28131\,
            in2 => \N__34481\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26949\,
            in2 => \N__34479\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27219\,
            in2 => \N__34482\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27174\,
            in2 => \N__34480\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28224\,
            in2 => \N__34483\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29767\,
            in2 => \_gnd_net_\,
            in3 => \N__25836\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34206\,
            in2 => \N__34178\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26721\,
            in2 => \N__26754\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27159\,
            in2 => \N__30346\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27279\,
            in2 => \N__30424\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30186\,
            in2 => \N__27168\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30705\,
            in2 => \N__30425\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29448\,
            in2 => \N__30347\,
            in3 => \N__25863\,
            lcout => \current_shift_inst.un38_control_input_0_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30141\,
            in2 => \N__27153\,
            in3 => \N__25854\,
            lcout => \current_shift_inst.un38_control_input_0_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28461\,
            in2 => \N__30274\,
            in3 => \N__25839\,
            lcout => \current_shift_inst.un38_control_input_0_s1_8\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26001\,
            in2 => \N__30426\,
            in3 => \N__25980\,
            lcout => \current_shift_inst.un38_control_input_0_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27273\,
            in2 => \N__30275\,
            in3 => \N__25968\,
            lcout => \current_shift_inst.un38_control_input_0_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27336\,
            in2 => \N__30427\,
            in3 => \N__25953\,
            lcout => \current_shift_inst.un38_control_input_0_s1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27348\,
            in2 => \N__30276\,
            in3 => \N__25938\,
            lcout => \current_shift_inst.un38_control_input_0_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27267\,
            in2 => \N__30428\,
            in3 => \N__25926\,
            lcout => \current_shift_inst.un38_control_input_0_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27285\,
            in2 => \N__30277\,
            in3 => \N__25908\,
            lcout => \current_shift_inst.un38_control_input_0_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27354\,
            in2 => \N__30429\,
            in3 => \N__25893\,
            lcout => \current_shift_inst.un38_control_input_0_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28236\,
            in2 => \N__30430\,
            in3 => \N__25878\,
            lcout => \current_shift_inst.un38_control_input_0_s1_16\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27255\,
            in2 => \N__30434\,
            in3 => \N__26127\,
            lcout => \current_shift_inst.un38_control_input_0_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27105\,
            in2 => \N__30431\,
            in3 => \N__26112\,
            lcout => \current_shift_inst.un38_control_input_0_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27318\,
            in2 => \N__30435\,
            in3 => \N__26094\,
            lcout => \current_shift_inst.un38_control_input_0_s1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27342\,
            in2 => \N__30432\,
            in3 => \N__26079\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27330\,
            in2 => \N__30436\,
            in3 => \N__26064\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27312\,
            in2 => \N__30433\,
            in3 => \N__26049\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27261\,
            in2 => \N__30437\,
            in3 => \N__26034\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30238\,
            in2 => \N__27513\,
            in3 => \N__26019\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27198\,
            in2 => \N__30442\,
            in3 => \N__26004\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28176\,
            in2 => \N__30458\,
            in3 => \N__26220\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27186\,
            in2 => \N__30443\,
            in3 => \N__26205\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27231\,
            in2 => \N__30459\,
            in3 => \N__26190\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27324\,
            in2 => \N__30444\,
            in3 => \N__26178\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28544\,
            in2 => \N__30460\,
            in3 => \N__26163\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_2_25_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__29809\,
            in1 => \N__30268\,
            in2 => \_gnd_net_\,
            in3 => \N__26160\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S1_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27486\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45932\,
            ce => 'H',
            sr => \N__45580\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31464\,
            in2 => \_gnd_net_\,
            in3 => \N__33258\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46014\,
            ce => \N__29322\,
            sr => \N__45480\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31463\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33327\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46006\,
            ce => \N__29321\,
            sr => \N__45485\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31886\,
            in2 => \_gnd_net_\,
            in3 => \N__35841\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46006\,
            ce => \N__29321\,
            sr => \N__45485\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011001000"
        )
    port map (
            in0 => \N__28704\,
            in1 => \N__35949\,
            in2 => \N__31895\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46006\,
            ce => \N__29321\,
            sr => \N__45485\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__31890\,
            in1 => \N__35907\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46006\,
            ce => \N__29321\,
            sr => \N__45485\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38076\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46006\,
            ce => \N__29321\,
            sr => \N__45485\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26295\,
            in2 => \N__27384\,
            in3 => \N__26311\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_10_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26277\,
            in2 => \N__27393\,
            in3 => \N__26288\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26256\,
            in2 => \N__27552\,
            in3 => \N__26267\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26238\,
            in2 => \N__27366\,
            in3 => \N__26249\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26484\,
            in2 => \N__26511\,
            in3 => \N__26495\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26466\,
            in2 => \N__27582\,
            in3 => \N__26477\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26459\,
            in1 => \N__26439\,
            in2 => \N__26448\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26432\,
            in1 => \N__26409\,
            in2 => \N__26421\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26391\,
            in2 => \N__27375\,
            in3 => \N__26402\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_10_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26373\,
            in2 => \N__27564\,
            in3 => \N__26384\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26340\,
            in2 => \N__26367\,
            in3 => \N__26351\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26322\,
            in2 => \N__27573\,
            in3 => \N__26333\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26643\,
            in2 => \N__26667\,
            in3 => \N__26654\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26625\,
            in2 => \N__27408\,
            in3 => \N__26636\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26607\,
            in2 => \N__27543\,
            in3 => \N__26618\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26571\,
            in2 => \N__26601\,
            in3 => \N__26589\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26564\,
            in1 => \N__26553\,
            in2 => \N__26802\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26546\,
            in1 => \N__26535\,
            in2 => \N__26793\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26517\,
            in2 => \N__26784\,
            in3 => \N__26528\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26805\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43775\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45977\,
            ce => \N__29316\,
            sr => \N__45505\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43557\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45977\,
            ce => \N__29316\,
            sr => \N__45505\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38043\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45977\,
            ce => \N__29316\,
            sr => \N__45505\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26694\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30910\,
            in1 => \N__32332\,
            in2 => \_gnd_net_\,
            in3 => \N__29464\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__27626\,
            in1 => \N__26696\,
            in2 => \N__26769\,
            in3 => \N__29534\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30911\,
            in1 => \N__32287\,
            in2 => \_gnd_net_\,
            in3 => \N__27793\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__27625\,
            in1 => \N__26695\,
            in2 => \_gnd_net_\,
            in3 => \N__30907\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30908\,
            in1 => \N__31679\,
            in2 => \_gnd_net_\,
            in3 => \N__29251\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__30673\,
            in1 => \N__29535\,
            in2 => \N__32208\,
            in3 => \N__27764\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30909\,
            in1 => \N__31562\,
            in2 => \_gnd_net_\,
            in3 => \N__30721\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32119\,
            in1 => \N__30918\,
            in2 => \_gnd_net_\,
            in3 => \N__28330\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__31633\,
            in1 => \_gnd_net_\,
            in2 => \N__30942\,
            in3 => \N__27601\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32236\,
            in1 => \N__30916\,
            in2 => \_gnd_net_\,
            in3 => \N__28474\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__30494\,
            in1 => \N__29732\,
            in2 => \N__32337\,
            in3 => \N__29465\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32084\,
            in1 => \N__30919\,
            in2 => \_gnd_net_\,
            in3 => \N__27730\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30917\,
            in1 => \N__32197\,
            in2 => \_gnd_net_\,
            in3 => \N__27763\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__31600\,
            in1 => \N__30915\,
            in2 => \_gnd_net_\,
            in3 => \N__28426\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__31634\,
            in1 => \N__29731\,
            in2 => \N__30610\,
            in3 => \N__27602\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__32167\,
            in1 => \N__28363\,
            in2 => \_gnd_net_\,
            in3 => \N__30920\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30921\,
            in1 => \N__32041\,
            in2 => \_gnd_net_\,
            in3 => \N__27695\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32605\,
            in1 => \N__30923\,
            in2 => \_gnd_net_\,
            in3 => \N__28261\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29630\,
            in1 => \N__32080\,
            in2 => \N__30692\,
            in3 => \N__27731\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32644\,
            in1 => \N__30922\,
            in2 => \_gnd_net_\,
            in3 => \N__28297\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30925\,
            in1 => \N__32521\,
            in2 => \_gnd_net_\,
            in3 => \N__27881\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32446\,
            in1 => \N__30926\,
            in2 => \_gnd_net_\,
            in3 => \N__28075\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30924\,
            in1 => \N__32568\,
            in2 => \_gnd_net_\,
            in3 => \N__28577\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30947\,
            in1 => \N__32867\,
            in2 => \_gnd_net_\,
            in3 => \N__28204\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30943\,
            in1 => \N__32473\,
            in2 => \_gnd_net_\,
            in3 => \N__27862\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30945\,
            in1 => \N__32404\,
            in2 => \_gnd_net_\,
            in3 => \N__28111\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32932\,
            in1 => \N__30946\,
            in2 => \_gnd_net_\,
            in3 => \N__27827\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32899\,
            in1 => \N__30944\,
            in2 => \_gnd_net_\,
            in3 => \N__28039\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29697\,
            in1 => \N__32818\,
            in2 => \_gnd_net_\,
            in3 => \N__27997\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__27863\,
            in1 => \N__29698\,
            in2 => \N__32480\,
            in3 => \N__30679\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27017\,
            lcout => \current_shift_inst.N_1819_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29733\,
            in1 => \N__32749\,
            in2 => \_gnd_net_\,
            in3 => \N__27973\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__28400\,
            in1 => \N__29736\,
            in2 => \N__32723\,
            in3 => \N__30471\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29734\,
            in1 => \N__32716\,
            in2 => \_gnd_net_\,
            in3 => \N__28399\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__29705\,
            in1 => \N__27998\,
            in2 => \N__30602\,
            in3 => \N__32819\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__27999\,
            in1 => \N__29706\,
            in2 => \N__32823\,
            in3 => \N__30475\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__27974\,
            in1 => \N__29735\,
            in2 => \N__32756\,
            in3 => \N__30470\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32680\,
            in1 => \N__29704\,
            in2 => \_gnd_net_\,
            in3 => \N__27943\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29703\,
            in1 => \N__31608\,
            in2 => \N__30603\,
            in3 => \N__28437\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29699\,
            in1 => \N__31680\,
            in2 => \N__30624\,
            in3 => \N__29259\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29707\,
            in1 => \N__32291\,
            in2 => \N__30620\,
            in3 => \N__27806\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__27950\,
            in1 => \N__29709\,
            in2 => \N__30623\,
            in3 => \N__32688\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32646\,
            in1 => \N__29702\,
            in2 => \N__30621\,
            in3 => \N__28308\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29700\,
            in1 => \N__31641\,
            in2 => \N__30625\,
            in3 => \N__27609\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29708\,
            in1 => \N__32169\,
            in2 => \N__30619\,
            in3 => \N__28374\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29701\,
            in1 => \N__32045\,
            in2 => \N__30622\,
            in3 => \N__27707\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29821\,
            in1 => \N__32906\,
            in2 => \N__30678\,
            in3 => \N__28050\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32522\,
            in1 => \N__29820\,
            in2 => \N__30667\,
            in3 => \N__27893\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29815\,
            in1 => \N__32247\,
            in2 => \N__30664\,
            in3 => \N__28485\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29819\,
            in1 => \N__32046\,
            in2 => \N__30677\,
            in3 => \N__27711\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29816\,
            in1 => \N__32607\,
            in2 => \N__30666\,
            in3 => \N__28272\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29818\,
            in1 => \N__32085\,
            in2 => \N__30676\,
            in3 => \N__27738\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29817\,
            in1 => \N__32411\,
            in2 => \N__30665\,
            in3 => \N__28122\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29803\,
            in1 => \N__32126\,
            in2 => \N__30688\,
            in3 => \N__28341\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29822\,
            in1 => \N__32373\,
            in2 => \N__30668\,
            in3 => \N__30834\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29823\,
            in1 => \N__32687\,
            in2 => \N__30670\,
            in3 => \N__27954\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__32448\,
            in1 => \N__30588\,
            in2 => \N__29844\,
            in3 => \N__28086\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__27837\,
            in1 => \N__29808\,
            in2 => \N__30669\,
            in3 => \N__32940\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29807\,
            in1 => \N__32939\,
            in2 => \N__30689\,
            in3 => \N__27836\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__28212\,
            in1 => \N__29824\,
            in2 => \N__30671\,
            in3 => \N__32868\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_2_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__27439\,
            in1 => \N__31760\,
            in2 => \N__27472\,
            in3 => \N__40794\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46023\,
            ce => 'H',
            sr => \N__45458\
        );

    \phase_controller_inst2.state_3_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__27441\,
            in1 => \N__27504\,
            in2 => \N__27473\,
            in3 => \N__30969\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46015\,
            ce => 'H',
            sr => \N__45465\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__33434\,
            in1 => \N__31996\,
            in2 => \_gnd_net_\,
            in3 => \N__31936\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27462\,
            in2 => \_gnd_net_\,
            in3 => \N__27440\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__33440\,
            in1 => \N__32001\,
            in2 => \_gnd_net_\,
            in3 => \N__31938\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45997\,
            ce => \N__29320\,
            sr => \N__45481\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__28598\,
            in1 => \N__36368\,
            in2 => \N__31896\,
            in3 => \N__28687\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45997\,
            ce => \N__29320\,
            sr => \N__45481\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__28686\,
            in1 => \N__31891\,
            in2 => \N__36488\,
            in3 => \N__28597\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45997\,
            ce => \N__29320\,
            sr => \N__45481\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011101111"
        )
    port map (
            in0 => \N__33384\,
            in1 => \N__31998\,
            in2 => \N__33132\,
            in3 => \N__31482\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45986\,
            ce => \N__29280\,
            sr => \N__45486\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__35989\,
            in1 => \_gnd_net_\,
            in2 => \N__28691\,
            in3 => \N__31885\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45986\,
            ce => \N__29280\,
            sr => \N__45486\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__31883\,
            in1 => \N__28671\,
            in2 => \_gnd_net_\,
            in3 => \N__35729\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45986\,
            ce => \N__29280\,
            sr => \N__45486\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31480\,
            in2 => \_gnd_net_\,
            in3 => \N__33302\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45986\,
            ce => \N__29280\,
            sr => \N__45486\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31481\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33357\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45986\,
            ce => \N__29280\,
            sr => \N__45486\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__28667\,
            in1 => \N__28619\,
            in2 => \N__35795\,
            in3 => \N__31884\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45986\,
            ce => \N__29280\,
            sr => \N__45486\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31997\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33433\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45986\,
            ce => \N__29280\,
            sr => \N__45486\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27653\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29691\,
            in2 => \N__27531\,
            in3 => \N__29214\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32863\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32565\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_1_25_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29690\,
            in2 => \_gnd_net_\,
            in3 => \N__30614\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29211\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__29212\,
            in1 => \_gnd_net_\,
            in2 => \N__27663\,
            in3 => \N__30859\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32993\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45972\,
            ce => \N__32965\,
            sr => \N__45496\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33695\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45972\,
            ce => \N__32965\,
            sr => \N__45496\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27660\,
            in2 => \N__27654\,
            in3 => \N__27652\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30735\,
            in2 => \_gnd_net_\,
            in3 => \N__27612\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31689\,
            in2 => \_gnd_net_\,
            in3 => \N__27588\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28716\,
            in2 => \_gnd_net_\,
            in3 => \N__27585\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29433\,
            in2 => \_gnd_net_\,
            in3 => \N__27813\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28710\,
            in2 => \_gnd_net_\,
            in3 => \N__27810\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30741\,
            in2 => \_gnd_net_\,
            in3 => \N__27777\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29415\,
            in2 => \_gnd_net_\,
            in3 => \N__27774\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30789\,
            in2 => \_gnd_net_\,
            in3 => \N__27747\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30795\,
            in2 => \_gnd_net_\,
            in3 => \N__27744\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29427\,
            in2 => \_gnd_net_\,
            in3 => \N__27741\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29421\,
            in2 => \_gnd_net_\,
            in3 => \N__27714\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30765\,
            in2 => \_gnd_net_\,
            in3 => \N__27684\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30777\,
            in2 => \_gnd_net_\,
            in3 => \N__27924\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29409\,
            in2 => \_gnd_net_\,
            in3 => \N__27921\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27918\,
            in2 => \_gnd_net_\,
            in3 => \N__27909\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27906\,
            in2 => \_gnd_net_\,
            in3 => \N__27870\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30981\,
            in2 => \_gnd_net_\,
            in3 => \N__27849\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30993\,
            in2 => \_gnd_net_\,
            in3 => \N__27846\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30783\,
            in2 => \_gnd_net_\,
            in3 => \N__27843\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31005\,
            in3 => \N__27840\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30759\,
            in2 => \_gnd_net_\,
            in3 => \N__27816\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30771\,
            in2 => \_gnd_net_\,
            in3 => \N__28014\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28011\,
            in2 => \_gnd_net_\,
            in3 => \N__28002\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30753\,
            in2 => \_gnd_net_\,
            in3 => \N__27984\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30975\,
            in2 => \_gnd_net_\,
            in3 => \N__27981\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30987\,
            in2 => \_gnd_net_\,
            in3 => \N__27960\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30747\,
            in2 => \_gnd_net_\,
            in3 => \N__27957\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28164\,
            in2 => \_gnd_net_\,
            in3 => \N__27930\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27927\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28227\,
            in3 => \N__29782\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29783\,
            in1 => \N__32856\,
            in2 => \N__30693\,
            in3 => \N__28205\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__29813\,
            in1 => \N__28143\,
            in2 => \N__30605\,
            in3 => \N__32783\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32679\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__28142\,
            in1 => \N__29812\,
            in2 => \N__32784\,
            in3 => \N__30482\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__29810\,
            in1 => \N__28141\,
            in2 => \_gnd_net_\,
            in3 => \N__32779\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29842\,
            in1 => \N__32412\,
            in2 => \N__30606\,
            in3 => \N__28118\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29811\,
            in1 => \N__32447\,
            in2 => \N__30604\,
            in3 => \N__28082\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__29833\,
            in1 => \N__28046\,
            in2 => \N__30568\,
            in3 => \N__32907\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101111"
        )
    port map (
            in0 => \N__28481\,
            in1 => \N__30393\,
            in2 => \N__29846\,
            in3 => \N__32243\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__30830\,
            in1 => \N__29832\,
            in2 => \N__30567\,
            in3 => \N__32369\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29828\,
            in1 => \N__31607\,
            in2 => \N__30569\,
            in3 => \N__28433\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29843\,
            in1 => \N__32724\,
            in2 => \N__30566\,
            in3 => \N__28404\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29836\,
            in1 => \N__32168\,
            in2 => \N__30686\,
            in3 => \N__28370\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__30647\,
            in1 => \N__29837\,
            in2 => \N__32127\,
            in3 => \N__28337\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101111"
        )
    port map (
            in0 => \N__28304\,
            in1 => \N__30648\,
            in2 => \N__29847\,
            in3 => \N__32645\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__28268\,
            in1 => \N__29841\,
            in2 => \N__30687\,
            in3 => \N__32606\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__28584\,
            in1 => \N__29835\,
            in2 => \N__30691\,
            in3 => \N__32567\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29834\,
            in1 => \N__32566\,
            in2 => \N__30690\,
            in3 => \N__28583\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29845\,
            in2 => \_gnd_net_\,
            in3 => \N__28557\,
            lcout => \current_shift_inst.un4_control_input_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28501\,
            in2 => \_gnd_net_\,
            in3 => \N__37644\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_463_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__33062\,
            in1 => \N__31077\,
            in2 => \N__45623\,
            in3 => \N__31094\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__33068\,
            in1 => \N__31076\,
            in2 => \_gnd_net_\,
            in3 => \N__31093\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46022\,
            ce => 'H',
            sr => \N__45452\
        );

    \delay_measurement_inst.prev_tr_sig_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33069\,
            lcout => \delay_measurement_inst.prev_tr_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46022\,
            ce => 'H',
            sr => \N__45452\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__28505\,
            in1 => \N__28518\,
            in2 => \_gnd_net_\,
            in3 => \N__37649\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46022\,
            ce => 'H',
            sr => \N__45452\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31759\,
            in2 => \_gnd_net_\,
            in3 => \N__40793\,
            lcout => \phase_controller_inst2.start_timer_hc_RNO_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__28517\,
            in1 => \N__28506\,
            in2 => \_gnd_net_\,
            in3 => \N__37648\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_464_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__28699\,
            in1 => \N__35948\,
            in2 => \_gnd_net_\,
            in3 => \N__31882\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46005\,
            ce => \N__35369\,
            sr => \N__45459\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__28698\,
            in1 => \N__35997\,
            in2 => \_gnd_net_\,
            in3 => \N__31881\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46005\,
            ce => \N__35369\,
            sr => \N__45459\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43776\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46005\,
            ce => \N__35369\,
            sr => \N__45459\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__28605\,
            in1 => \N__36372\,
            in2 => \N__28703\,
            in3 => \N__31880\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46005\,
            ce => \N__35369\,
            sr => \N__45459\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__31879\,
            in1 => \N__28694\,
            in2 => \N__36489\,
            in3 => \N__28604\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46005\,
            ce => \N__35369\,
            sr => \N__45459\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__32000\,
            in1 => \N__33435\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45996\,
            ce => \N__35374\,
            sr => \N__45466\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__31875\,
            in1 => \N__28693\,
            in2 => \_gnd_net_\,
            in3 => \N__35733\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45996\,
            ce => \N__35374\,
            sr => \N__45466\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31462\,
            in2 => \_gnd_net_\,
            in3 => \N__33303\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45996\,
            ce => \N__35374\,
            sr => \N__45466\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31999\,
            in2 => \N__33441\,
            in3 => \N__31937\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45996\,
            ce => \N__35374\,
            sr => \N__45466\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__28692\,
            in1 => \N__28623\,
            in2 => \N__35799\,
            in3 => \N__31877\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45996\,
            ce => \N__35374\,
            sr => \N__45466\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31876\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35906\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45996\,
            ce => \N__35374\,
            sr => \N__45466\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35840\,
            in2 => \_gnd_net_\,
            in3 => \N__31878\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45996\,
            ce => \N__35374\,
            sr => \N__45466\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31461\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33257\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45996\,
            ce => \N__35374\,
            sr => \N__45466\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31465\,
            in2 => \_gnd_net_\,
            in3 => \N__33356\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45985\,
            ce => \N__35370\,
            sr => \N__45473\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31917\,
            in1 => \N__35941\,
            in2 => \N__35996\,
            in3 => \N__31966\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__28638\,
            in1 => \N__33127\,
            in2 => \_gnd_net_\,
            in3 => \N__31967\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__35833\,
            in1 => \N__35899\,
            in2 => \_gnd_net_\,
            in3 => \N__35728\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28632\,
            in1 => \N__33450\,
            in2 => \N__28626\,
            in3 => \N__33102\,
            lcout => \phase_controller_inst1.stoper_tr.N_257\,
            ltout => \phase_controller_inst1.stoper_tr.N_257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36367\,
            in2 => \N__28608\,
            in3 => \N__35788\,
            lcout => \phase_controller_inst1.stoper_tr.N_240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a3_1_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29373\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38217\,
            lcout => state_ns_i_a3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__29104\,
            in1 => \N__28769\,
            in2 => \_gnd_net_\,
            in3 => \N__28887\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29581\,
            in1 => \N__31672\,
            in2 => \N__30674\,
            in3 => \N__29252\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__29580\,
            in1 => \N__29220\,
            in2 => \_gnd_net_\,
            in3 => \N__29213\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__28866\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28751\,
            lcout => \phase_controller_inst2.stoper_tr.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_0_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__28767\,
            in1 => \N__28883\,
            in2 => \N__29115\,
            in3 => \N__29159\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45962\,
            ce => \N__42507\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_1_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__29160\,
            in1 => \N__29111\,
            in2 => \N__28927\,
            in3 => \N__28768\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45962\,
            ce => \N__42507\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31590\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32313\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32268\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31657\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29799\,
            in1 => \N__31550\,
            in2 => \N__30675\,
            in3 => \N__30722\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__30615\,
            in1 => \N__29800\,
            in2 => \N__32336\,
            in3 => \N__29466\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31549\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32101\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32067\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32227\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32587\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32148\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32187\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32394\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32626\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32889\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32022\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32923\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32803\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32707\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32356\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32428\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32740\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32464\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32771\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__30968\,
            in1 => \N__36149\,
            in2 => \N__36115\,
            in3 => \N__37623\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45947\,
            ce => 'H',
            sr => \N__45531\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30948\,
            in1 => \N__32357\,
            in2 => \_gnd_net_\,
            in3 => \N__30829\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__31159\,
            in1 => \N__31187\,
            in2 => \_gnd_net_\,
            in3 => \N__31137\,
            lcout => \current_shift_inst.timer_s1.N_186_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31158\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36095\,
            in2 => \_gnd_net_\,
            in3 => \N__36148\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__31186\,
            in1 => \N__31160\,
            in2 => \_gnd_net_\,
            in3 => \N__31136\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45940\,
            ce => 'H',
            sr => \N__45543\
        );

    \current_shift_inst.start_timer_s1_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__33007\,
            in1 => \N__31182\,
            in2 => \_gnd_net_\,
            in3 => \N__36110\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45937\,
            ce => 'H',
            sr => \N__45552\
        );

    \current_shift_inst.stop_timer_s1_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__36111\,
            in1 => \N__33008\,
            in2 => \N__31188\,
            in3 => \N__31135\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45937\,
            ce => 'H',
            sr => \N__45552\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31161\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31131\,
            lcout => \current_shift_inst.timer_s1.N_185_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__33061\,
            in1 => \N__31075\,
            in2 => \_gnd_net_\,
            in3 => \N__31095\,
            lcout => \delay_measurement_inst.tr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46034\,
            ce => \N__42508\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__31059\,
            in1 => \N__38231\,
            in2 => \N__44559\,
            in3 => \N__31044\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46024\,
            ce => 'H',
            sr => \N__45453\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31038\,
            in2 => \N__31032\,
            in3 => \N__35311\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31011\,
            in2 => \N__31023\,
            in3 => \N__35294\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31305\,
            in2 => \N__31314\,
            in3 => \N__35261\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31287\,
            in2 => \N__31299\,
            in3 => \N__35237\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31272\,
            in2 => \N__31281\,
            in3 => \N__35510\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31257\,
            in2 => \N__31266\,
            in3 => \N__35486\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31239\,
            in2 => \N__31251\,
            in3 => \N__42197\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31218\,
            in2 => \N__31233\,
            in3 => \N__42155\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31212\,
            in2 => \N__31506\,
            in3 => \N__42119\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35456\,
            in1 => \N__31194\,
            in2 => \N__31206\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35435\,
            in1 => \N__31416\,
            in2 => \N__31428\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31398\,
            in2 => \N__31410\,
            in3 => \N__35414\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31383\,
            in2 => \N__31392\,
            in3 => \N__35654\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31365\,
            in2 => \N__31377\,
            in3 => \N__35630\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31350\,
            in2 => \N__31359\,
            in3 => \N__35609\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31344\,
            in2 => \N__31494\,
            in3 => \N__38118\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31326\,
            in2 => \N__31338\,
            in3 => \N__35579\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31320\,
            in2 => \N__31524\,
            in3 => \N__35555\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31533\,
            in2 => \N__31515\,
            in3 => \N__35534\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31527\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43556\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45998\,
            ce => \N__35379\,
            sr => \N__45467\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38037\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45998\,
            ce => \N__35379\,
            sr => \N__45467\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000101"
        )
    port map (
            in0 => \N__31478\,
            in1 => \N__31979\,
            in2 => \N__33131\,
            in3 => \N__33377\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45987\,
            ce => \N__35378\,
            sr => \N__45474\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38075\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45987\,
            ce => \N__35378\,
            sr => \N__45474\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31479\,
            in2 => \_gnd_net_\,
            in3 => \N__33320\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45987\,
            ce => \N__35378\,
            sr => \N__45474\
        );

    \delay_measurement_inst.delay_tr_reg_esr_14_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__38511\,
            in1 => \N__43661\,
            in2 => \N__31809\,
            in3 => \N__43728\,
            lcout => measured_delay_tr_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45978\,
            ce => \N__43520\,
            sr => \N__45482\
        );

    \delay_measurement_inst.delay_tr_reg_esr_15_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__43729\,
            in1 => \N__37994\,
            in2 => \N__43676\,
            in3 => \N__38460\,
            lcout => measured_delay_tr_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45978\,
            ce => \N__43520\,
            sr => \N__45482\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110001"
        )
    port map (
            in0 => \N__31971\,
            in1 => \N__31918\,
            in2 => \N__33439\,
            in3 => \N__33101\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_RNO_0_14_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__43660\,
            in1 => \N__37993\,
            in2 => \_gnd_net_\,
            in3 => \N__38459\,
            lcout => \delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__43285\,
            in1 => \N__43083\,
            in2 => \_gnd_net_\,
            in3 => \N__43429\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_1_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__31800\,
            in1 => \N__31770\,
            in2 => \N__31726\,
            in3 => \N__40792\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45968\,
            ce => 'H',
            sr => \N__45490\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31624\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33696\,
            in2 => \N__33632\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__45963\,
            ce => \N__32964\,
            sr => \N__45497\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33605\,
            in2 => \N__33665\,
            in3 => \N__31611\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__45963\,
            ce => \N__32964\,
            sr => \N__45497\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33584\,
            in2 => \N__33633\,
            in3 => \N__31569\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__45963\,
            ce => \N__32964\,
            sr => \N__45497\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33606\,
            in2 => \N__33563\,
            in3 => \N__31536\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__45963\,
            ce => \N__32964\,
            sr => \N__45497\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33585\,
            in2 => \N__33537\,
            in3 => \N__32295\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__45963\,
            ce => \N__32964\,
            sr => \N__45497\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33503\,
            in2 => \N__33564\,
            in3 => \N__32250\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__45963\,
            ce => \N__32964\,
            sr => \N__45497\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33533\,
            in2 => \N__33476\,
            in3 => \N__32211\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__45963\,
            ce => \N__32964\,
            sr => \N__45497\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33504\,
            in2 => \N__33902\,
            in3 => \N__32172\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__45963\,
            ce => \N__32964\,
            sr => \N__45497\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33872\,
            in2 => \N__33480\,
            in3 => \N__32130\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__45957\,
            ce => \N__32963\,
            sr => \N__45506\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33845\,
            in2 => \N__33909\,
            in3 => \N__32088\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__45957\,
            ce => \N__32963\,
            sr => \N__45506\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33824\,
            in2 => \N__33876\,
            in3 => \N__32049\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__45957\,
            ce => \N__32963\,
            sr => \N__45506\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33846\,
            in2 => \N__33803\,
            in3 => \N__32004\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__45957\,
            ce => \N__32963\,
            sr => \N__45506\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33825\,
            in2 => \N__33776\,
            in3 => \N__32610\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__45957\,
            ce => \N__32963\,
            sr => \N__45506\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33746\,
            in2 => \N__33804\,
            in3 => \N__32571\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__45957\,
            ce => \N__32963\,
            sr => \N__45506\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33715\,
            in2 => \N__33777\,
            in3 => \N__32529\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__45957\,
            ce => \N__32963\,
            sr => \N__45506\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33747\,
            in2 => \N__34145\,
            in3 => \N__32487\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__45957\,
            ce => \N__32963\,
            sr => \N__45506\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34118\,
            in2 => \N__33723\,
            in3 => \N__32451\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__45953\,
            ce => \N__32962\,
            sr => \N__45514\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34094\,
            in2 => \N__34152\,
            in3 => \N__32415\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__45953\,
            ce => \N__32962\,
            sr => \N__45514\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34119\,
            in2 => \N__34073\,
            in3 => \N__32376\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__45953\,
            ce => \N__32962\,
            sr => \N__45514\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34095\,
            in2 => \N__34043\,
            in3 => \N__32340\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__45953\,
            ce => \N__32962\,
            sr => \N__45514\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34016\,
            in2 => \N__34074\,
            in3 => \N__32910\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__45953\,
            ce => \N__32962\,
            sr => \N__45514\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33995\,
            in2 => \N__34044\,
            in3 => \N__32871\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__45953\,
            ce => \N__32962\,
            sr => \N__45514\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34017\,
            in2 => \N__33962\,
            in3 => \N__32826\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__45953\,
            ce => \N__32962\,
            sr => \N__45514\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33925\,
            in2 => \N__33996\,
            in3 => \N__32787\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__45953\,
            ce => \N__32962\,
            sr => \N__45514\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34922\,
            in2 => \N__33966\,
            in3 => \N__32760\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__45950\,
            ce => \N__32961\,
            sr => \N__45523\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34895\,
            in2 => \N__33936\,
            in3 => \N__32727\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__45950\,
            ce => \N__32961\,
            sr => \N__45523\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34875\,
            in2 => \N__34926\,
            in3 => \N__32691\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__45950\,
            ce => \N__32961\,
            sr => \N__45523\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34896\,
            in2 => \N__34719\,
            in3 => \N__32652\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__45950\,
            ce => \N__32961\,
            sr => \N__45523\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32649\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32978\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45950\,
            ce => \N__32961\,
            sr => \N__45523\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43114\,
            in1 => \N__43470\,
            in2 => \N__43338\,
            in3 => \N__36504\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45948\,
            ce => 'H',
            sr => \N__45532\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43115\,
            in1 => \N__43471\,
            in2 => \N__43339\,
            in3 => \N__36294\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45948\,
            ce => 'H',
            sr => \N__45532\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43468\,
            in1 => \N__43316\,
            in2 => \N__43127\,
            in3 => \N__36246\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45948\,
            ce => 'H',
            sr => \N__45532\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__43116\,
            in1 => \N__36213\,
            in2 => \N__43340\,
            in3 => \N__43473\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45948\,
            ce => 'H',
            sr => \N__45532\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43469\,
            in1 => \N__43317\,
            in2 => \N__43128\,
            in3 => \N__36180\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45948\,
            ce => 'H',
            sr => \N__45532\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43117\,
            in1 => \N__43472\,
            in2 => \N__43341\,
            in3 => \N__36618\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45948\,
            ce => 'H',
            sr => \N__45532\
        );

    \phase_controller_inst1.stoper_hc.target_time_0_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__42078\,
            in1 => \N__41522\,
            in2 => \N__46941\,
            in3 => \N__41750\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45945\,
            ce => \N__38932\,
            sr => \N__45539\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__41747\,
            in1 => \N__46918\,
            in2 => \N__41538\,
            in3 => \N__40991\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45945\,
            ce => \N__38932\,
            sr => \N__45539\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__41123\,
            in1 => \N__41525\,
            in2 => \N__46944\,
            in3 => \N__41753\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45945\,
            ce => \N__38932\,
            sr => \N__45539\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__41521\,
            in1 => \N__46754\,
            in2 => \N__41376\,
            in3 => \N__46921\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45945\,
            ce => \N__38932\,
            sr => \N__45539\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__41071\,
            in1 => \N__41523\,
            in2 => \N__46942\,
            in3 => \N__41751\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45945\,
            ce => \N__38932\,
            sr => \N__45539\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__41749\,
            in1 => \N__46920\,
            in2 => \N__41540\,
            in3 => \N__40945\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45945\,
            ce => \N__38932\,
            sr => \N__45539\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__41034\,
            in1 => \N__41524\,
            in2 => \N__46943\,
            in3 => \N__41752\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45945\,
            ce => \N__38932\,
            sr => \N__45539\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__41748\,
            in1 => \N__46919\,
            in2 => \N__41539\,
            in3 => \N__41816\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45945\,
            ce => \N__38932\,
            sr => \N__45539\
        );

    \phase_controller_inst1.S1_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36116\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45941\,
            ce => 'H',
            sr => \N__45544\
        );

    \delay_measurement_inst.delay_hc_reg_3_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__46274\,
            in1 => \N__42401\,
            in2 => \N__46498\,
            in3 => \N__41622\,
            lcout => measured_delay_hc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45938\,
            ce => 'H',
            sr => \N__45553\
        );

    \delay_measurement_inst.delay_hc_reg_8_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__39530\,
            in1 => \N__46481\,
            in2 => \N__40937\,
            in3 => \N__46275\,
            lcout => measured_delay_hc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45938\,
            ce => 'H',
            sr => \N__45553\
        );

    \delay_measurement_inst.delay_hc_reg_13_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__39240\,
            in1 => \N__46473\,
            in2 => \N__41817\,
            in3 => \N__46271\,
            lcout => measured_delay_hc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45938\,
            ce => 'H',
            sr => \N__45553\
        );

    \delay_measurement_inst.delay_hc_reg_21_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__39554\,
            in1 => \N__46474\,
            in2 => \_gnd_net_\,
            in3 => \N__46272\,
            lcout => measured_delay_hc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45938\,
            ce => 'H',
            sr => \N__45553\
        );

    \delay_measurement_inst.delay_hc_reg_22_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__46273\,
            in1 => \_gnd_net_\,
            in2 => \N__46497\,
            in3 => \N__39173\,
            lcout => measured_delay_hc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45938\,
            ce => 'H',
            sr => \N__45553\
        );

    \SB_DFF_inst_DELAY_TR1_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33087\,
            lcout => delay_tr_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR2_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33075\,
            lcout => delay_tr_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__42630\,
            in1 => \N__42797\,
            in2 => \N__42960\,
            in3 => \N__42673\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46035\,
            ce => \N__42509\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__42621\,
            in1 => \N__42951\,
            in2 => \N__42805\,
            in3 => \N__35445\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46025\,
            ce => 'H',
            sr => \N__45454\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__38156\,
            in1 => \N__35315\,
            in2 => \_gnd_net_\,
            in3 => \N__42672\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42624\,
            in1 => \N__42950\,
            in2 => \N__33024\,
            in3 => \N__42780\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46025\,
            ce => 'H',
            sr => \N__45454\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__35424\,
            in1 => \N__42625\,
            in2 => \N__42808\,
            in3 => \N__42947\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46025\,
            ce => 'H',
            sr => \N__45454\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__42622\,
            in1 => \N__42952\,
            in2 => \N__42806\,
            in3 => \N__35403\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46025\,
            ce => 'H',
            sr => \N__45454\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42948\,
            in1 => \N__42626\,
            in2 => \N__35643\,
            in3 => \N__42775\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46025\,
            ce => 'H',
            sr => \N__45454\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__42623\,
            in1 => \N__42953\,
            in2 => \N__42807\,
            in3 => \N__35619\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46025\,
            ce => 'H',
            sr => \N__45454\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42949\,
            in1 => \N__42627\,
            in2 => \N__35598\,
            in3 => \N__42776\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46025\,
            ce => 'H',
            sr => \N__45454\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42603\,
            in1 => \N__42934\,
            in2 => \N__35568\,
            in3 => \N__42789\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => 'H',
            sr => \N__45456\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42785\,
            in1 => \N__42607\,
            in2 => \N__42955\,
            in3 => \N__35544\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => 'H',
            sr => \N__45456\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42604\,
            in1 => \N__42935\,
            in2 => \N__35520\,
            in3 => \N__42790\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => 'H',
            sr => \N__45456\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42786\,
            in1 => \N__42608\,
            in2 => \N__42956\,
            in3 => \N__35283\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => 'H',
            sr => \N__45456\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42605\,
            in1 => \N__42936\,
            in2 => \N__35250\,
            in3 => \N__42791\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => 'H',
            sr => \N__45456\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42787\,
            in1 => \N__42609\,
            in2 => \N__42957\,
            in3 => \N__35226\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => 'H',
            sr => \N__45456\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42606\,
            in1 => \N__42937\,
            in2 => \N__35499\,
            in3 => \N__42792\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => 'H',
            sr => \N__45456\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42788\,
            in1 => \N__42610\,
            in2 => \N__42958\,
            in3 => \N__35475\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46016\,
            ce => 'H',
            sr => \N__45456\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__33231\,
            in1 => \N__33204\,
            in2 => \_gnd_net_\,
            in3 => \N__33177\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38149\,
            in2 => \_gnd_net_\,
            in3 => \N__42659\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42581\,
            in2 => \_gnd_net_\,
            in3 => \N__42781\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed11\,
            ltout => \phase_controller_inst1.stoper_tr.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33135\,
            in3 => \N__42658\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_15_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45618\,
            in2 => \_gnd_net_\,
            in3 => \N__36415\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33289\,
            in1 => \N__33319\,
            in2 => \N__33250\,
            in3 => \N__33343\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33105\,
            in3 => \N__33376\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43542\,
            in1 => \N__43761\,
            in2 => \N__38041\,
            in3 => \N__38073\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__43543\,
            in1 => \N__43762\,
            in2 => \N__38042\,
            in3 => \N__38074\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__38627\,
            in1 => \N__43707\,
            in2 => \N__38469\,
            in3 => \N__35685\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.N_360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_9_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001110"
        )
    port map (
            in0 => \N__38628\,
            in1 => \N__33273\,
            in2 => \N__33387\,
            in3 => \N__43671\,
            lcout => measured_delay_tr_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45988\,
            ce => \N__43519\,
            sr => \N__45475\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001110"
        )
    port map (
            in0 => \N__38464\,
            in1 => \N__38510\,
            in2 => \N__37995\,
            in3 => \N__43706\,
            lcout => \delay_measurement_inst.N_354\,
            ltout => \delay_measurement_inst.N_354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_10_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43665\,
            in2 => \N__33360\,
            in3 => \N__38589\,
            lcout => measured_delay_tr_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45988\,
            ce => \N__43519\,
            sr => \N__45475\
        );

    \delay_measurement_inst.delay_tr_reg_esr_11_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__38568\,
            in1 => \N__43666\,
            in2 => \_gnd_net_\,
            in3 => \N__33270\,
            lcout => measured_delay_tr_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45988\,
            ce => \N__43519\,
            sr => \N__45475\
        );

    \delay_measurement_inst.delay_tr_reg_esr_12_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__33271\,
            in1 => \_gnd_net_\,
            in2 => \N__43677\,
            in3 => \N__38550\,
            lcout => measured_delay_tr_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45988\,
            ce => \N__43519\,
            sr => \N__45475\
        );

    \delay_measurement_inst.delay_tr_reg_esr_13_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__38532\,
            in1 => \N__33272\,
            in2 => \_gnd_net_\,
            in3 => \N__43670\,
            lcout => measured_delay_tr_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45988\,
            ce => \N__43519\,
            sr => \N__45475\
        );

    \current_shift_inst.timer_s1.counter_0_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34842\,
            in1 => \N__33688\,
            in2 => \_gnd_net_\,
            in3 => \N__33669\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__45979\,
            ce => \N__34700\,
            sr => \N__45483\
        );

    \current_shift_inst.timer_s1.counter_1_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34850\,
            in1 => \N__33652\,
            in2 => \_gnd_net_\,
            in3 => \N__33636\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__45979\,
            ce => \N__34700\,
            sr => \N__45483\
        );

    \current_shift_inst.timer_s1.counter_2_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34843\,
            in1 => \N__33625\,
            in2 => \_gnd_net_\,
            in3 => \N__33609\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__45979\,
            ce => \N__34700\,
            sr => \N__45483\
        );

    \current_shift_inst.timer_s1.counter_3_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34851\,
            in1 => \N__33604\,
            in2 => \_gnd_net_\,
            in3 => \N__33588\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__45979\,
            ce => \N__34700\,
            sr => \N__45483\
        );

    \current_shift_inst.timer_s1.counter_4_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34844\,
            in1 => \N__33583\,
            in2 => \_gnd_net_\,
            in3 => \N__33567\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__45979\,
            ce => \N__34700\,
            sr => \N__45483\
        );

    \current_shift_inst.timer_s1.counter_5_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34852\,
            in1 => \N__33556\,
            in2 => \_gnd_net_\,
            in3 => \N__33540\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__45979\,
            ce => \N__34700\,
            sr => \N__45483\
        );

    \current_shift_inst.timer_s1.counter_6_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34845\,
            in1 => \N__33529\,
            in2 => \_gnd_net_\,
            in3 => \N__33507\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__45979\,
            ce => \N__34700\,
            sr => \N__45483\
        );

    \current_shift_inst.timer_s1.counter_7_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34853\,
            in1 => \N__33497\,
            in2 => \_gnd_net_\,
            in3 => \N__33483\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__45979\,
            ce => \N__34700\,
            sr => \N__45483\
        );

    \current_shift_inst.timer_s1.counter_8_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34841\,
            in1 => \N__33475\,
            in2 => \_gnd_net_\,
            in3 => \N__33453\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__45973\,
            ce => \N__34701\,
            sr => \N__45487\
        );

    \current_shift_inst.timer_s1.counter_9_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34837\,
            in1 => \N__33901\,
            in2 => \_gnd_net_\,
            in3 => \N__33879\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__45973\,
            ce => \N__34701\,
            sr => \N__45487\
        );

    \current_shift_inst.timer_s1.counter_10_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34838\,
            in1 => \N__33865\,
            in2 => \_gnd_net_\,
            in3 => \N__33849\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__45973\,
            ce => \N__34701\,
            sr => \N__45487\
        );

    \current_shift_inst.timer_s1.counter_11_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34834\,
            in1 => \N__33844\,
            in2 => \_gnd_net_\,
            in3 => \N__33828\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__45973\,
            ce => \N__34701\,
            sr => \N__45487\
        );

    \current_shift_inst.timer_s1.counter_12_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34839\,
            in1 => \N__33823\,
            in2 => \_gnd_net_\,
            in3 => \N__33807\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__45973\,
            ce => \N__34701\,
            sr => \N__45487\
        );

    \current_shift_inst.timer_s1.counter_13_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34835\,
            in1 => \N__33796\,
            in2 => \_gnd_net_\,
            in3 => \N__33780\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__45973\,
            ce => \N__34701\,
            sr => \N__45487\
        );

    \current_shift_inst.timer_s1.counter_14_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34840\,
            in1 => \N__33764\,
            in2 => \_gnd_net_\,
            in3 => \N__33750\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__45973\,
            ce => \N__34701\,
            sr => \N__45487\
        );

    \current_shift_inst.timer_s1.counter_15_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34836\,
            in1 => \N__33740\,
            in2 => \_gnd_net_\,
            in3 => \N__33726\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__45973\,
            ce => \N__34701\,
            sr => \N__45487\
        );

    \current_shift_inst.timer_s1.counter_16_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34846\,
            in1 => \N__33719\,
            in2 => \_gnd_net_\,
            in3 => \N__33699\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__45969\,
            ce => \N__34696\,
            sr => \N__45491\
        );

    \current_shift_inst.timer_s1.counter_17_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34854\,
            in1 => \N__34144\,
            in2 => \_gnd_net_\,
            in3 => \N__34122\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__45969\,
            ce => \N__34696\,
            sr => \N__45491\
        );

    \current_shift_inst.timer_s1.counter_18_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34847\,
            in1 => \N__34112\,
            in2 => \_gnd_net_\,
            in3 => \N__34098\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__45969\,
            ce => \N__34696\,
            sr => \N__45491\
        );

    \current_shift_inst.timer_s1.counter_19_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34855\,
            in1 => \N__34093\,
            in2 => \_gnd_net_\,
            in3 => \N__34077\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__45969\,
            ce => \N__34696\,
            sr => \N__45491\
        );

    \current_shift_inst.timer_s1.counter_20_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34848\,
            in1 => \N__34061\,
            in2 => \_gnd_net_\,
            in3 => \N__34047\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__45969\,
            ce => \N__34696\,
            sr => \N__45491\
        );

    \current_shift_inst.timer_s1.counter_21_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34856\,
            in1 => \N__34036\,
            in2 => \_gnd_net_\,
            in3 => \N__34020\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__45969\,
            ce => \N__34696\,
            sr => \N__45491\
        );

    \current_shift_inst.timer_s1.counter_22_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34849\,
            in1 => \N__34015\,
            in2 => \_gnd_net_\,
            in3 => \N__33999\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__45969\,
            ce => \N__34696\,
            sr => \N__45491\
        );

    \current_shift_inst.timer_s1.counter_23_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34857\,
            in1 => \N__33988\,
            in2 => \_gnd_net_\,
            in3 => \N__33969\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__45969\,
            ce => \N__34696\,
            sr => \N__45491\
        );

    \current_shift_inst.timer_s1.counter_24_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34830\,
            in1 => \N__33961\,
            in2 => \_gnd_net_\,
            in3 => \N__33939\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__45964\,
            ce => \N__34695\,
            sr => \N__45498\
        );

    \current_shift_inst.timer_s1.counter_25_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34774\,
            in1 => \N__33929\,
            in2 => \_gnd_net_\,
            in3 => \N__34929\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__45964\,
            ce => \N__34695\,
            sr => \N__45498\
        );

    \current_shift_inst.timer_s1.counter_26_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34831\,
            in1 => \N__34915\,
            in2 => \_gnd_net_\,
            in3 => \N__34899\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__45964\,
            ce => \N__34695\,
            sr => \N__45498\
        );

    \current_shift_inst.timer_s1.counter_27_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34775\,
            in1 => \N__34894\,
            in2 => \_gnd_net_\,
            in3 => \N__34878\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__45964\,
            ce => \N__34695\,
            sr => \N__45498\
        );

    \current_shift_inst.timer_s1.counter_28_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34832\,
            in1 => \N__34874\,
            in2 => \_gnd_net_\,
            in3 => \N__34860\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__45964\,
            ce => \N__34695\,
            sr => \N__45498\
        );

    \current_shift_inst.timer_s1.counter_29_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__34715\,
            in1 => \N__34833\,
            in2 => \_gnd_net_\,
            in3 => \N__34722\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45964\,
            ce => \N__34695\,
            sr => \N__45498\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__41940\,
            in1 => \N__40902\,
            in2 => \N__41541\,
            in3 => \N__46934\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45958\,
            ce => \N__38925\,
            sr => \N__45507\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__34653\,
            in1 => \N__34574\,
            in2 => \_gnd_net_\,
            in3 => \N__34629\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__34575\,
            in1 => \_gnd_net_\,
            in2 => \N__34209\,
            in3 => \N__34205\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43098\,
            in1 => \N__43446\,
            in2 => \N__43331\,
            in3 => \N__36579\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45954\,
            ce => 'H',
            sr => \N__45515\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__43156\,
            in1 => \N__39098\,
            in2 => \_gnd_net_\,
            in3 => \N__36332\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__43290\,
            in1 => \N__43101\,
            in2 => \N__34962\,
            in3 => \N__43449\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45954\,
            ce => 'H',
            sr => \N__45515\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43444\,
            in1 => \N__43291\,
            in2 => \N__43124\,
            in3 => \N__36555\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45954\,
            ce => 'H',
            sr => \N__45515\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43099\,
            in1 => \N__43447\,
            in2 => \N__43332\,
            in3 => \N__36531\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45954\,
            ce => 'H',
            sr => \N__45515\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43100\,
            in1 => \N__43448\,
            in2 => \N__43333\,
            in3 => \N__36735\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45954\,
            ce => 'H',
            sr => \N__45515\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43445\,
            in1 => \N__43292\,
            in2 => \N__43125\,
            in3 => \N__36711\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45954\,
            ce => 'H',
            sr => \N__45515\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34959\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34941\,
            in2 => \N__34953\,
            in3 => \N__36328\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34935\,
            in2 => \N__39039\,
            in3 => \N__36305\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35046\,
            in2 => \N__38952\,
            in3 => \N__36272\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35031\,
            in2 => \N__35040\,
            in3 => \N__36224\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35025\,
            in2 => \N__38979\,
            in3 => \N__36191\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35019\,
            in2 => \N__38967\,
            in3 => \N__36629\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35013\,
            in2 => \N__39027\,
            in3 => \N__38871\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35007\,
            in2 => \N__35001\,
            in3 => \N__38847\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34983\,
            in2 => \N__34992\,
            in3 => \N__36860\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34968\,
            in2 => \N__34977\,
            in3 => \N__36594\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35112\,
            in2 => \N__35124\,
            in3 => \N__36570\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36546\,
            in1 => \N__35097\,
            in2 => \N__35106\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36515\,
            in1 => \N__35082\,
            in2 => \N__35091\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35076\,
            in2 => \N__38994\,
            in3 => \N__36750\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35070\,
            in2 => \N__39012\,
            in3 => \N__36726\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35064\,
            in2 => \N__36822\,
            in3 => \N__36702\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35058\,
            in2 => \N__36813\,
            in3 => \N__36884\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35052\,
            in2 => \N__36804\,
            in3 => \N__36842\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36647\,
            in1 => \N__35136\,
            in2 => \N__36831\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35130\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35127\,
            in3 => \N__39097\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_9_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__46270\,
            in1 => \N__41360\,
            in2 => \N__46496\,
            in3 => \N__39138\,
            lcout => measured_delay_hc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45942\,
            ce => 'H',
            sr => \N__45545\
        );

    \delay_measurement_inst.delay_hc_reg_14_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011101110"
        )
    port map (
            in0 => \N__39156\,
            in1 => \N__46465\,
            in2 => \N__41592\,
            in3 => \N__46267\,
            lcout => measured_delay_hc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45942\,
            ce => 'H',
            sr => \N__45545\
        );

    \delay_measurement_inst.delay_hc_reg_23_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__46268\,
            in1 => \_gnd_net_\,
            in2 => \N__46495\,
            in3 => \N__39188\,
            lcout => measured_delay_hc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45942\,
            ce => 'H',
            sr => \N__45545\
        );

    \delay_measurement_inst.delay_hc_reg_24_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__39203\,
            in1 => \N__46469\,
            in2 => \_gnd_net_\,
            in3 => \N__46269\,
            lcout => measured_delay_hc_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45942\,
            ce => 'H',
            sr => \N__45545\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBOIH1_14_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__46292\,
            in1 => \N__39154\,
            in2 => \N__42400\,
            in3 => \N__39136\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36794\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45934\,
            ce => \N__37856\,
            sr => \N__45558\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36773\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45934\,
            ce => \N__37856\,
            sr => \N__45558\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37772\,
            in1 => \N__36790\,
            in2 => \_gnd_net_\,
            in3 => \N__35163\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__45933\,
            ce => \N__37818\,
            sr => \N__45564\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37768\,
            in1 => \N__36769\,
            in2 => \_gnd_net_\,
            in3 => \N__35160\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__45933\,
            ce => \N__37818\,
            sr => \N__45564\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37773\,
            in1 => \N__37111\,
            in2 => \_gnd_net_\,
            in3 => \N__35157\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__45933\,
            ce => \N__37818\,
            sr => \N__45564\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37769\,
            in1 => \N__37079\,
            in2 => \_gnd_net_\,
            in3 => \N__35154\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__45933\,
            ce => \N__37818\,
            sr => \N__45564\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37774\,
            in1 => \N__37055\,
            in2 => \_gnd_net_\,
            in3 => \N__35151\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__45933\,
            ce => \N__37818\,
            sr => \N__45564\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37770\,
            in1 => \N__37031\,
            in2 => \_gnd_net_\,
            in3 => \N__35148\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__45933\,
            ce => \N__37818\,
            sr => \N__45564\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37775\,
            in1 => \N__37001\,
            in2 => \_gnd_net_\,
            in3 => \N__35145\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__45933\,
            ce => \N__37818\,
            sr => \N__45564\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37771\,
            in1 => \N__36971\,
            in2 => \_gnd_net_\,
            in3 => \N__35142\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__45933\,
            ce => \N__37818\,
            sr => \N__45564\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37736\,
            in1 => \N__36943\,
            in2 => \_gnd_net_\,
            in3 => \N__35139\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__45931\,
            ce => \N__37810\,
            sr => \N__45568\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37726\,
            in1 => \N__36913\,
            in2 => \_gnd_net_\,
            in3 => \N__35190\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__45931\,
            ce => \N__37810\,
            sr => \N__45568\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37733\,
            in1 => \N__37357\,
            in2 => \_gnd_net_\,
            in3 => \N__35187\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__45931\,
            ce => \N__37810\,
            sr => \N__45568\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37723\,
            in1 => \N__37325\,
            in2 => \_gnd_net_\,
            in3 => \N__35184\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__45931\,
            ce => \N__37810\,
            sr => \N__45568\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37734\,
            in1 => \N__37306\,
            in2 => \_gnd_net_\,
            in3 => \N__35181\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__45931\,
            ce => \N__37810\,
            sr => \N__45568\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37724\,
            in1 => \N__37280\,
            in2 => \_gnd_net_\,
            in3 => \N__35178\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__45931\,
            ce => \N__37810\,
            sr => \N__45568\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37735\,
            in1 => \N__37250\,
            in2 => \_gnd_net_\,
            in3 => \N__35175\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__45931\,
            ce => \N__37810\,
            sr => \N__45568\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37725\,
            in1 => \N__37220\,
            in2 => \_gnd_net_\,
            in3 => \N__35172\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__45931\,
            ce => \N__37810\,
            sr => \N__45568\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37776\,
            in1 => \N__37195\,
            in2 => \_gnd_net_\,
            in3 => \N__35169\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_27_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__45929\,
            ce => \N__37811\,
            sr => \N__45571\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37764\,
            in1 => \N__37165\,
            in2 => \_gnd_net_\,
            in3 => \N__35166\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__45929\,
            ce => \N__37811\,
            sr => \N__45571\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37777\,
            in1 => \N__37135\,
            in2 => \_gnd_net_\,
            in3 => \N__35217\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__45929\,
            ce => \N__37811\,
            sr => \N__45571\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37765\,
            in1 => \N__37595\,
            in2 => \_gnd_net_\,
            in3 => \N__35214\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__45929\,
            ce => \N__37811\,
            sr => \N__45571\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37778\,
            in1 => \N__37571\,
            in2 => \_gnd_net_\,
            in3 => \N__35211\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__45929\,
            ce => \N__37811\,
            sr => \N__45571\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37766\,
            in1 => \N__37547\,
            in2 => \_gnd_net_\,
            in3 => \N__35208\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__45929\,
            ce => \N__37811\,
            sr => \N__45571\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37779\,
            in1 => \N__37517\,
            in2 => \_gnd_net_\,
            in3 => \N__35205\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__45929\,
            ce => \N__37811\,
            sr => \N__45571\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37767\,
            in1 => \N__37487\,
            in2 => \_gnd_net_\,
            in3 => \N__35202\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__45929\,
            ce => \N__37811\,
            sr => \N__45571\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37727\,
            in1 => \N__37462\,
            in2 => \_gnd_net_\,
            in3 => \N__35199\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_28_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__45928\,
            ce => \N__37809\,
            sr => \N__45574\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37731\,
            in1 => \N__37432\,
            in2 => \_gnd_net_\,
            in3 => \N__35196\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__45928\,
            ce => \N__37809\,
            sr => \N__45574\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37728\,
            in1 => \N__37384\,
            in2 => \_gnd_net_\,
            in3 => \N__35193\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__45928\,
            ce => \N__37809\,
            sr => \N__45574\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37732\,
            in1 => \N__37882\,
            in2 => \_gnd_net_\,
            in3 => \N__35394\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__45928\,
            ce => \N__37809\,
            sr => \N__45574\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37729\,
            in1 => \N__37406\,
            in2 => \_gnd_net_\,
            in3 => \N__35391\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__45928\,
            ce => \N__37809\,
            sr => \N__45574\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__37904\,
            in1 => \N__37730\,
            in2 => \_gnd_net_\,
            in3 => \N__35388\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45928\,
            ce => \N__37809\,
            sr => \N__45574\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35385\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__42848\,
            in1 => \N__42620\,
            in2 => \_gnd_net_\,
            in3 => \N__42753\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35325\,
            in2 => \N__35316\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35295\,
            in2 => \_gnd_net_\,
            in3 => \N__35277\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35274\,
            in2 => \N__35265\,
            in3 => \N__35241\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35238\,
            in2 => \_gnd_net_\,
            in3 => \N__35220\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35511\,
            in2 => \_gnd_net_\,
            in3 => \N__35490\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35487\,
            in2 => \_gnd_net_\,
            in3 => \N__35469\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42198\,
            in2 => \_gnd_net_\,
            in3 => \N__35466\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42156\,
            in2 => \_gnd_net_\,
            in3 => \N__35463\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42120\,
            in2 => \_gnd_net_\,
            in3 => \N__35460\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35457\,
            in2 => \_gnd_net_\,
            in3 => \N__35439\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35436\,
            in2 => \_gnd_net_\,
            in3 => \N__35418\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35415\,
            in2 => \_gnd_net_\,
            in3 => \N__35397\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35655\,
            in2 => \_gnd_net_\,
            in3 => \N__35634\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35631\,
            in2 => \_gnd_net_\,
            in3 => \N__35613\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35610\,
            in2 => \_gnd_net_\,
            in3 => \N__35586\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38114\,
            in2 => \_gnd_net_\,
            in3 => \N__35583\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35580\,
            in2 => \_gnd_net_\,
            in3 => \N__35559\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35556\,
            in2 => \_gnd_net_\,
            in3 => \N__35538\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35535\,
            in2 => \_gnd_net_\,
            in3 => \N__35523\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_6_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38508\,
            in1 => \N__38614\,
            in2 => \N__38468\,
            in3 => \N__38259\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__35742\,
            in1 => \N__38337\,
            in2 => \N__43674\,
            in3 => \N__35673\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111110"
        )
    port map (
            in0 => \N__37976\,
            in1 => \N__35697\,
            in2 => \N__43675\,
            in3 => \N__43705\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31\,
            ltout => \delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_6_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001101"
        )
    port map (
            in0 => \N__35672\,
            in1 => \N__38442\,
            in2 => \N__35736\,
            in3 => \N__38262\,
            lcout => measured_delay_tr_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46007\,
            ce => \N__43511\,
            sr => \N__45460\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_15_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__37953\,
            in1 => \N__35671\,
            in2 => \N__38458\,
            in3 => \N__35706\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38546\,
            in1 => \N__38564\,
            in2 => \N__38531\,
            in3 => \N__38582\,
            lcout => \delay_measurement_inst.N_381\,
            ltout => \delay_measurement_inst.N_381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010001"
        )
    port map (
            in0 => \N__38451\,
            in1 => \N__38501\,
            in2 => \N__35700\,
            in3 => \N__38615\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIE5AP1_23_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38817\,
            in1 => \N__38826\,
            in2 => \N__38808\,
            in3 => \N__38679\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38694\,
            in1 => \N__35751\,
            in2 => \N__35691\,
            in3 => \N__40335\,
            lcout => \delay_measurement_inst.N_498\,
            ltout => \delay_measurement_inst.N_498_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__38642\,
            in1 => \N__38663\,
            in2 => \N__35688\,
            in3 => \N__35684\,
            lcout => \delay_measurement_inst.N_384\,
            ltout => \delay_measurement_inst.N_384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3UDFH_6_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__38452\,
            in1 => \N__35852\,
            in2 => \N__36000\,
            in3 => \N__38261\,
            lcout => \delay_measurement_inst.delay_tr_reg_5_tz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_4_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38298\,
            in1 => \N__36388\,
            in2 => \N__35982\,
            in3 => \N__36431\,
            lcout => measured_delay_tr_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45989\,
            ce => 'H',
            sr => \N__45476\
        );

    \delay_measurement_inst.delay_tr_reg_5_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__36432\,
            in1 => \N__35926\,
            in2 => \N__36397\,
            in3 => \N__38280\,
            lcout => measured_delay_tr_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45989\,
            ce => 'H',
            sr => \N__45476\
        );

    \delay_measurement_inst.delay_tr_reg_7_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38670\,
            in1 => \N__35858\,
            in2 => \N__35898\,
            in3 => \N__36433\,
            lcout => measured_delay_tr_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45989\,
            ce => 'H',
            sr => \N__45476\
        );

    \delay_measurement_inst.delay_tr_reg_8_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__36434\,
            in1 => \N__35823\,
            in2 => \N__35862\,
            in3 => \N__38649\,
            lcout => measured_delay_tr_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45989\,
            ce => 'H',
            sr => \N__45476\
        );

    \delay_measurement_inst.start_timer_hc_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__40719\,
            in1 => \N__40865\,
            in2 => \_gnd_net_\,
            in3 => \N__40759\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45989\,
            ce => 'H',
            sr => \N__45476\
        );

    \delay_measurement_inst.delay_tr_reg_3_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38316\,
            in1 => \N__36387\,
            in2 => \N__35787\,
            in3 => \N__36430\,
            lcout => measured_delay_tr_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45989\,
            ce => 'H',
            sr => \N__45476\
        );

    \phase_controller_inst1.state_1_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__38402\,
            in1 => \N__36069\,
            in2 => \N__36048\,
            in3 => \N__37932\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45989\,
            ce => 'H',
            sr => \N__45476\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38778\,
            in1 => \N__38787\,
            in2 => \N__38769\,
            in3 => \N__38796\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36064\,
            in2 => \_gnd_net_\,
            in3 => \N__36036\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.start_timer_hc_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__43227\,
            in1 => \N__36165\,
            in2 => \N__36153\,
            in3 => \N__38230\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45974\,
            ce => 'H',
            sr => \N__45488\
        );

    \phase_controller_inst1.state_2_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__36150\,
            in1 => \N__36065\,
            in2 => \N__36044\,
            in3 => \N__36117\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45974\,
            ce => 'H',
            sr => \N__45488\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__36040\,
            in1 => \N__39099\,
            in2 => \N__40881\,
            in3 => \N__43165\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45974\,
            ce => 'H',
            sr => \N__45488\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43396\,
            in1 => \N__43069\,
            in2 => \N__43283\,
            in3 => \N__36684\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45974\,
            ce => 'H',
            sr => \N__45488\
        );

    \delay_measurement_inst.delay_hc_reg_7_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__39408\,
            in1 => \N__46491\,
            in2 => \N__41238\,
            in3 => \N__46281\,
            lcout => measured_delay_hc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45970\,
            ce => 'H',
            sr => \N__45492\
        );

    \delay_measurement_inst.delay_hc_reg_4_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__46279\,
            in1 => \N__41118\,
            in2 => \N__46499\,
            in3 => \N__39429\,
            lcout => measured_delay_hc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45970\,
            ce => 'H',
            sr => \N__45492\
        );

    \delay_measurement_inst.delay_hc_reg_30_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41321\,
            in1 => \N__46484\,
            in2 => \_gnd_net_\,
            in3 => \N__46278\,
            lcout => measured_delay_hc_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45970\,
            ce => 'H',
            sr => \N__45492\
        );

    \delay_measurement_inst.delay_hc_reg_5_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__46280\,
            in1 => \N__41186\,
            in2 => \N__46500\,
            in3 => \N__42372\,
            lcout => measured_delay_hc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45970\,
            ce => 'H',
            sr => \N__45492\
        );

    \phase_controller_inst1.S2_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37945\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45970\,
            ce => 'H',
            sr => \N__45492\
        );

    \delay_measurement_inst.delay_tr_reg_1_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__43854\,
            in1 => \N__36398\,
            in2 => \N__36475\,
            in3 => \N__36440\,
            lcout => measured_delay_tr_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45970\,
            ce => 'H',
            sr => \N__45492\
        );

    \delay_measurement_inst.delay_tr_reg_2_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__36441\,
            in1 => \N__36349\,
            in2 => \N__36402\,
            in3 => \N__38367\,
            lcout => measured_delay_tr_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45970\,
            ce => 'H',
            sr => \N__45492\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__37838\,
            in1 => \N__40837\,
            in2 => \_gnd_net_\,
            in3 => \N__39847\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45970\,
            ce => 'H',
            sr => \N__45492\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36663\,
            in2 => \N__36333\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36312\,
            in2 => \_gnd_net_\,
            in3 => \N__36282\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36279\,
            in2 => \N__36261\,
            in3 => \N__36234\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36231\,
            in2 => \_gnd_net_\,
            in3 => \N__36201\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36198\,
            in2 => \_gnd_net_\,
            in3 => \N__36168\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36636\,
            in2 => \_gnd_net_\,
            in3 => \N__36606\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38870\,
            in2 => \_gnd_net_\,
            in3 => \N__36603\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38843\,
            in2 => \_gnd_net_\,
            in3 => \N__36600\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36864\,
            in2 => \_gnd_net_\,
            in3 => \N__36597\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36593\,
            in2 => \_gnd_net_\,
            in3 => \N__36573\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36569\,
            in2 => \_gnd_net_\,
            in3 => \N__36549\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36545\,
            in2 => \_gnd_net_\,
            in3 => \N__36525\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36522\,
            in2 => \_gnd_net_\,
            in3 => \N__36492\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36749\,
            in2 => \_gnd_net_\,
            in3 => \N__36729\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36725\,
            in2 => \_gnd_net_\,
            in3 => \N__36705\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36701\,
            in2 => \_gnd_net_\,
            in3 => \N__36675\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36885\,
            in2 => \_gnd_net_\,
            in3 => \N__36672\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36843\,
            in2 => \_gnd_net_\,
            in3 => \N__36669\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36648\,
            in2 => \_gnd_net_\,
            in3 => \N__36666\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39078\,
            in2 => \_gnd_net_\,
            in3 => \N__43155\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43110\,
            in1 => \N__43453\,
            in2 => \N__43336\,
            in3 => \N__36654\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45951\,
            ce => 'H',
            sr => \N__45524\
        );

    \delay_measurement_inst.delay_hc_reg_10_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__46439\,
            in1 => \N__39219\,
            in2 => \N__41075\,
            in3 => \N__46255\,
            lcout => measured_delay_hc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45951\,
            ce => 'H',
            sr => \N__45524\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43108\,
            in1 => \N__43452\,
            in2 => \N__43334\,
            in3 => \N__36891\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45951\,
            ce => 'H',
            sr => \N__45524\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100010001100"
        )
    port map (
            in0 => \N__43451\,
            in1 => \N__36873\,
            in2 => \N__43126\,
            in3 => \N__43311\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45951\,
            ce => 'H',
            sr => \N__45524\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__43109\,
            in1 => \N__36849\,
            in2 => \N__43335\,
            in3 => \N__43454\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45951\,
            ce => 'H',
            sr => \N__45524\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46730\,
            in2 => \_gnd_net_\,
            in3 => \N__47021\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45949\,
            ce => \N__38937\,
            sr => \N__45533\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__46731\,
            in1 => \N__46995\,
            in2 => \_gnd_net_\,
            in3 => \N__46830\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45949\,
            ce => \N__38937\,
            sr => \N__45533\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__46828\,
            in1 => \N__46732\,
            in2 => \_gnd_net_\,
            in3 => \N__46643\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45949\,
            ce => \N__38937\,
            sr => \N__45533\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__46829\,
            in1 => \N__46733\,
            in2 => \_gnd_net_\,
            in3 => \N__41868\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45949\,
            ce => \N__38937\,
            sr => \N__45533\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36795\,
            in2 => \N__37118\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__45946\,
            ce => \N__37860\,
            sr => \N__45540\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36774\,
            in2 => \N__37091\,
            in3 => \N__36753\,
            lcout => \delay_measurement_inst.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__45946\,
            ce => \N__37860\,
            sr => \N__45540\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37061\,
            in2 => \N__37119\,
            in3 => \N__37095\,
            lcout => \delay_measurement_inst.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__45946\,
            ce => \N__37860\,
            sr => \N__45540\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37037\,
            in2 => \N__37092\,
            in3 => \N__37065\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__45946\,
            ce => \N__37860\,
            sr => \N__45540\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37062\,
            in2 => \N__37013\,
            in3 => \N__37041\,
            lcout => \delay_measurement_inst.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__45946\,
            ce => \N__37860\,
            sr => \N__45540\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37038\,
            in2 => \N__36983\,
            in3 => \N__37017\,
            lcout => \delay_measurement_inst.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__45946\,
            ce => \N__37860\,
            sr => \N__45540\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36953\,
            in2 => \N__37014\,
            in3 => \N__36987\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__45946\,
            ce => \N__37860\,
            sr => \N__45540\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36921\,
            in2 => \N__36984\,
            in3 => \N__36957\,
            lcout => \delay_measurement_inst.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__45946\,
            ce => \N__37860\,
            sr => \N__45540\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36954\,
            in2 => \N__37364\,
            in3 => \N__36924\,
            lcout => \delay_measurement_inst.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__45943\,
            ce => \N__37859\,
            sr => \N__45546\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36920\,
            in2 => \N__37337\,
            in3 => \N__36894\,
            lcout => \delay_measurement_inst.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__45943\,
            ce => \N__37859\,
            sr => \N__45546\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37307\,
            in2 => \N__37365\,
            in3 => \N__37341\,
            lcout => \delay_measurement_inst.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__45943\,
            ce => \N__37859\,
            sr => \N__45546\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37286\,
            in2 => \N__37338\,
            in3 => \N__37311\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__45943\,
            ce => \N__37859\,
            sr => \N__45546\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37308\,
            in2 => \N__37262\,
            in3 => \N__37290\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__45943\,
            ce => \N__37859\,
            sr => \N__45546\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37287\,
            in2 => \N__37232\,
            in3 => \N__37266\,
            lcout => \delay_measurement_inst.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__45943\,
            ce => \N__37859\,
            sr => \N__45546\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37203\,
            in2 => \N__37263\,
            in3 => \N__37236\,
            lcout => \delay_measurement_inst.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__45943\,
            ce => \N__37859\,
            sr => \N__45546\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37173\,
            in2 => \N__37233\,
            in3 => \N__37206\,
            lcout => \delay_measurement_inst.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__45943\,
            ce => \N__37859\,
            sr => \N__45546\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37202\,
            in2 => \N__37142\,
            in3 => \N__37176\,
            lcout => \delay_measurement_inst.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__45939\,
            ce => \N__37858\,
            sr => \N__45554\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37172\,
            in2 => \N__37607\,
            in3 => \N__37146\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__45939\,
            ce => \N__37858\,
            sr => \N__45554\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37577\,
            in2 => \N__37143\,
            in3 => \N__37611\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__45939\,
            ce => \N__37858\,
            sr => \N__45554\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37553\,
            in2 => \N__37608\,
            in3 => \N__37581\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__45939\,
            ce => \N__37858\,
            sr => \N__45554\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37578\,
            in2 => \N__37529\,
            in3 => \N__37557\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__45939\,
            ce => \N__37858\,
            sr => \N__45554\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37554\,
            in2 => \N__37499\,
            in3 => \N__37533\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__45939\,
            ce => \N__37858\,
            sr => \N__45554\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37470\,
            in2 => \N__37530\,
            in3 => \N__37503\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__45939\,
            ce => \N__37858\,
            sr => \N__45554\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37440\,
            in2 => \N__37500\,
            in3 => \N__37473\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__45939\,
            ce => \N__37858\,
            sr => \N__45554\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37469\,
            in2 => \N__37391\,
            in3 => \N__37443\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_15_25_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__45935\,
            ce => \N__37857\,
            sr => \N__45559\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37439\,
            in2 => \N__37889\,
            in3 => \N__37413\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__45935\,
            ce => \N__37857\,
            sr => \N__45559\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37410\,
            in2 => \N__37392\,
            in3 => \N__37368\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__45935\,
            ce => \N__37857\,
            sr => \N__45559\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37908\,
            in2 => \N__37890\,
            in3 => \N__37866\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__45935\,
            ce => \N__37857\,
            sr => \N__45559\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37863\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45935\,
            ce => \N__37857\,
            sr => \N__45559\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__37839\,
            in1 => \N__40842\,
            in2 => \_gnd_net_\,
            in3 => \N__39864\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_462_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39863\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39788\,
            lcout => \delay_measurement_inst.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46060\,
            ce => \N__43825\,
            sr => \N__45440\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI104I_2_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38509\,
            in2 => \_gnd_net_\,
            in3 => \N__38356\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__42849\,
            in1 => \N__42629\,
            in2 => \_gnd_net_\,
            in3 => \N__42793\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37653\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38095\,
            in2 => \_gnd_net_\,
            in3 => \N__38084\,
            lcout => \phase_controller_inst1.state_RNI7NN7Z0Z_0\,
            ltout => \phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__38376\,
            in1 => \N__42918\,
            in2 => \N__38235\,
            in3 => \N__38232\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46044\,
            ce => 'H',
            sr => \N__45443\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__38099\,
            in1 => \N__38160\,
            in2 => \N__38133\,
            in3 => \N__42681\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46044\,
            ce => 'H',
            sr => \N__45443\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__42628\,
            in1 => \N__42812\,
            in2 => \N__42954\,
            in3 => \N__38124\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46044\,
            ce => 'H',
            sr => \N__45443\
        );

    \phase_controller_inst1.state_0_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__38085\,
            in1 => \N__37947\,
            in2 => \N__38100\,
            in3 => \N__38401\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46044\,
            ce => 'H',
            sr => \N__45443\
        );

    \delay_measurement_inst.delay_tr_reg_esr_16_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__43721\,
            in1 => \N__43647\,
            in2 => \_gnd_net_\,
            in3 => \N__38751\,
            lcout => measured_delay_tr_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46036\,
            ce => \N__43521\,
            sr => \N__45446\
        );

    \delay_measurement_inst.delay_tr_reg_esr_19_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__43722\,
            in1 => \N__43648\,
            in2 => \_gnd_net_\,
            in3 => \N__38720\,
            lcout => measured_delay_tr_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46036\,
            ce => \N__43521\,
            sr => \N__45446\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__38750\,
            in1 => \N__38719\,
            in2 => \N__43806\,
            in3 => \N__43577\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16\,
            ltout => \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH1A23_1_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__38331\,
            in1 => \N__38322\,
            in2 => \N__37965\,
            in3 => \N__37962\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37946\,
            in2 => \_gnd_net_\,
            in3 => \N__38403\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__43576\,
            in1 => \N__38311\,
            in2 => \N__38721\,
            in3 => \N__38363\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__43801\,
            in1 => \N__38749\,
            in2 => \N__38340\,
            in3 => \N__38330\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38276\,
            in2 => \_gnd_net_\,
            in3 => \N__38294\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_373_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__38613\,
            in1 => \N__38312\,
            in2 => \N__43850\,
            in3 => \N__38260\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43881\,
            in2 => \N__39758\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__46017\,
            ce => \N__43826\,
            sr => \N__45457\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39731\,
            in2 => \N__39795\,
            in3 => \N__38283\,
            lcout => \delay_measurement_inst.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__46017\,
            ce => \N__43826\,
            sr => \N__45457\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39710\,
            in2 => \N__39759\,
            in3 => \N__38265\,
            lcout => \delay_measurement_inst.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__46017\,
            ce => \N__43826\,
            sr => \N__45457\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39732\,
            in2 => \N__39681\,
            in3 => \N__38238\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__46017\,
            ce => \N__43826\,
            sr => \N__45457\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40079\,
            in2 => \N__39711\,
            in3 => \N__38652\,
            lcout => \delay_measurement_inst.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__46017\,
            ce => \N__43826\,
            sr => \N__45457\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39677\,
            in2 => \N__40058\,
            in3 => \N__38631\,
            lcout => \delay_measurement_inst.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__46017\,
            ce => \N__43826\,
            sr => \N__45457\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40080\,
            in2 => \N__40028\,
            in3 => \N__38592\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__46017\,
            ce => \N__43826\,
            sr => \N__45457\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39991\,
            in2 => \N__40059\,
            in3 => \N__38571\,
            lcout => \delay_measurement_inst.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__46017\,
            ce => \N__43826\,
            sr => \N__45457\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40029\,
            in2 => \N__39965\,
            in3 => \N__38553\,
            lcout => \delay_measurement_inst.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_16_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__46008\,
            ce => \N__43827\,
            sr => \N__45461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39938\,
            in2 => \N__39999\,
            in3 => \N__38535\,
            lcout => \delay_measurement_inst.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__46008\,
            ce => \N__43827\,
            sr => \N__45461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39917\,
            in2 => \N__39966\,
            in3 => \N__38514\,
            lcout => \delay_measurement_inst.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__46008\,
            ce => \N__43827\,
            sr => \N__45461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39939\,
            in2 => \N__39894\,
            in3 => \N__38472\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__46008\,
            ce => \N__43827\,
            sr => \N__45461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39918\,
            in2 => \N__40325\,
            in3 => \N__38754\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__46008\,
            ce => \N__43827\,
            sr => \N__45461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39890\,
            in2 => \N__40295\,
            in3 => \N__38730\,
            lcout => \delay_measurement_inst.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__46008\,
            ce => \N__43827\,
            sr => \N__45461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40268\,
            in2 => \N__40326\,
            in3 => \N__38727\,
            lcout => \delay_measurement_inst.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__46008\,
            ce => \N__43827\,
            sr => \N__45461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40232\,
            in2 => \N__40296\,
            in3 => \N__38724\,
            lcout => \delay_measurement_inst.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__46008\,
            ce => \N__43827\,
            sr => \N__45461\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40269\,
            in2 => \N__40208\,
            in3 => \N__38697\,
            lcout => \delay_measurement_inst.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__45999\,
            ce => \N__43829\,
            sr => \N__45468\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40236\,
            in2 => \N__40181\,
            in3 => \N__38688\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__45999\,
            ce => \N__43829\,
            sr => \N__45468\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40151\,
            in2 => \N__40209\,
            in3 => \N__38685\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__45999\,
            ce => \N__43829\,
            sr => \N__45468\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40121\,
            in2 => \N__40182\,
            in3 => \N__38682\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__45999\,
            ce => \N__43829\,
            sr => \N__45468\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40100\,
            in2 => \N__40152\,
            in3 => \N__38673\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__45999\,
            ce => \N__43829\,
            sr => \N__45468\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40122\,
            in2 => \N__40691\,
            in3 => \N__38820\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__45999\,
            ce => \N__43829\,
            sr => \N__45468\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40101\,
            in2 => \N__40664\,
            in3 => \N__38811\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__45999\,
            ce => \N__43829\,
            sr => \N__45468\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40628\,
            in2 => \N__40692\,
            in3 => \N__38799\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__45999\,
            ce => \N__43829\,
            sr => \N__45468\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40665\,
            in2 => \N__40601\,
            in3 => \N__38790\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_16_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__45990\,
            ce => \N__43830\,
            sr => \N__45477\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40574\,
            in2 => \N__40635\,
            in3 => \N__38781\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__45990\,
            ce => \N__43830\,
            sr => \N__45477\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40554\,
            in2 => \N__40602\,
            in3 => \N__38772\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__45990\,
            ce => \N__43830\,
            sr => \N__45477\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40575\,
            in2 => \N__40407\,
            in3 => \N__38760\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__45990\,
            ce => \N__43830\,
            sr => \N__45477\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38757\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45990\,
            ce => \N__43830\,
            sr => \N__45477\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__43046\,
            in1 => \N__43428\,
            in2 => \N__43284\,
            in3 => \N__43172\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45980\,
            ce => \N__42502\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_state_0_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__40708\,
            in1 => \N__40858\,
            in2 => \_gnd_net_\,
            in3 => \N__40760\,
            lcout => \delay_measurement_inst.hc_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45980\,
            ce => \N__42502\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0_3_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41644\,
            in1 => \N__46131\,
            in2 => \N__41187\,
            in3 => \N__41934\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__41224\,
            in1 => \N__41097\,
            in2 => \N__38889\,
            in3 => \N__42076\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.N_316_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto8_i_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101110"
        )
    port map (
            in0 => \N__40946\,
            in1 => \N__41293\,
            in2 => \N__38886\,
            in3 => \N__41225\,
            lcout => \phase_controller_inst1.stoper_hc.N_388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__43071\,
            in1 => \N__43315\,
            in2 => \N__38883\,
            in3 => \N__43443\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45965\,
            ce => 'H',
            sr => \N__45499\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43442\,
            in1 => \N__43072\,
            in2 => \N__43337\,
            in3 => \N__38853\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45965\,
            ce => 'H',
            sr => \N__45499\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto13_2_0_a2_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40970\,
            in2 => \_gnd_net_\,
            in3 => \N__41018\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlt31_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3_2_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__41070\,
            in1 => \N__41828\,
            in2 => \N__38829\,
            in3 => \N__42259\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_11_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__39258\,
            in1 => \N__46461\,
            in2 => \N__41029\,
            in3 => \N__46265\,
            lcout => measured_delay_hc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45965\,
            ce => 'H',
            sr => \N__45499\
        );

    \delay_measurement_inst.delay_hc_reg_12_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__46266\,
            in1 => \N__40971\,
            in2 => \N__46494\,
            in3 => \N__39276\,
            lcout => measured_delay_hc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45965\,
            ce => 'H',
            sr => \N__45499\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__41456\,
            in1 => \N__46130\,
            in2 => \N__41769\,
            in3 => \N__46914\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45959\,
            ce => \N__38933\,
            sr => \N__45508\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__46912\,
            in1 => \N__41746\,
            in2 => \N__41500\,
            in3 => \N__41241\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45959\,
            ce => \N__38933\,
            sr => \N__45508\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__41455\,
            in1 => \N__42261\,
            in2 => \N__41768\,
            in3 => \N__46913\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45959\,
            ce => \N__38933\,
            sr => \N__45508\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__46909\,
            in1 => \N__46746\,
            in2 => \N__41595\,
            in3 => \N__41458\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45959\,
            ce => \N__38933\,
            sr => \N__45508\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__41457\,
            in1 => \N__41191\,
            in2 => \N__41770\,
            in3 => \N__46915\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45959\,
            ce => \N__38933\,
            sr => \N__45508\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__46911\,
            in1 => \N__46747\,
            in2 => \N__41295\,
            in3 => \N__41460\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45959\,
            ce => \N__38933\,
            sr => \N__45508\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__46910\,
            in1 => \N__41646\,
            in2 => \N__41655\,
            in3 => \N__41459\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45959\,
            ce => \N__38933\,
            sr => \N__45508\
        );

    \phase_controller_inst1.stoper_hc.un3_start_i_0_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__41669\,
            in1 => \N__39108\,
            in2 => \N__42005\,
            in3 => \N__46702\,
            lcout => \phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_0_o2_1_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__41935\,
            in1 => \N__41637\,
            in2 => \_gnd_net_\,
            in3 => \N__46129\,
            lcout => \phase_controller_inst1.stoper_hc.N_406\,
            ltout => \phase_controller_inst1.stoper_hc.N_406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0_1_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__46701\,
            in1 => \N__41668\,
            in2 => \N__39102\,
            in3 => \N__47020\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43070\,
            in2 => \_gnd_net_\,
            in3 => \N__43397\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_8_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41282\,
            in1 => \N__41028\,
            in2 => \N__40990\,
            in3 => \N__41239\,
            lcout => \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_7_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41867\,
            in1 => \N__41373\,
            in2 => \N__41593\,
            in3 => \N__41119\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39060\,
            in1 => \N__39051\,
            in2 => \N__39054\,
            in3 => \N__39045\,
            lcout => \phase_controller_inst1.stoper_hc.N_459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_5_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__42257\,
            in1 => \N__46637\,
            in2 => \_gnd_net_\,
            in3 => \N__46983\,
            lcout => \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3_18_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__41582\,
            in1 => \N__39282\,
            in2 => \_gnd_net_\,
            in3 => \N__42258\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_6_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41069\,
            in1 => \N__40938\,
            in2 => \N__41827\,
            in3 => \N__41195\,
            lcout => \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_19_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41990\,
            in2 => \_gnd_net_\,
            in3 => \N__46791\,
            lcout => \phase_controller_inst1.stoper_hc.N_453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2_18_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__41859\,
            in1 => \N__46642\,
            in2 => \N__41998\,
            in3 => \N__46982\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TRB1_16_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41953\,
            in1 => \N__39424\,
            in2 => \N__39464\,
            in3 => \N__42358\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39269\,
            in1 => \N__39251\,
            in2 => \N__39236\,
            in3 => \N__39215\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7_19_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39204\,
            in1 => \N__46515\,
            in2 => \N__39486\,
            in3 => \N__39189\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7Z0Z_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_19_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__41304\,
            in1 => \N__39174\,
            in2 => \N__39159\,
            in3 => \N__39540\,
            lcout => \phase_controller_inst1.stoper_hc.N_449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__41954\,
            in1 => \N__41884\,
            in2 => \N__42044\,
            in3 => \N__39460\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_14_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__39155\,
            in1 => \N__39137\,
            in2 => \_gnd_net_\,
            in3 => \N__39307\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.N_299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGMFO5_15_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000000"
        )
    port map (
            in0 => \N__42278\,
            in1 => \N__39294\,
            in2 => \N__39120\,
            in3 => \N__39117\,
            lcout => \delay_measurement_inst.N_332\,
            ltout => \delay_measurement_inst.N_332_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICFUBH_31_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__39651\,
            in1 => \N__39363\,
            in2 => \N__39111\,
            in3 => \N__42306\,
            lcout => \delay_measurement_inst.N_298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42277\,
            in1 => \N__39523\,
            in2 => \N__39404\,
            in3 => \N__39425\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHVTL_7_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39397\,
            in2 => \_gnd_net_\,
            in3 => \N__42276\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_318_1\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_318_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO11I2_18_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__42040\,
            in1 => \N__41885\,
            in2 => \N__39384\,
            in3 => \N__39381\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_14_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__39375\,
            in1 => \N__39503\,
            in2 => \N__39366\,
            in3 => \N__39308\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__39357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39351\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__39345\,
            in1 => \N__39564\,
            in2 => \N__39336\,
            in3 => \N__39597\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_328\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOFS27_1_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39315\,
            in1 => \N__42345\,
            in2 => \N__39333\,
            in3 => \N__39330\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI71JB5_6_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__39321\,
            in1 => \N__39314\,
            in2 => \N__39504\,
            in3 => \N__39293\,
            lcout => \delay_measurement_inst.N_318\,
            ltout => \delay_measurement_inst.N_318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDM4FI_31_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39647\,
            in1 => \N__39633\,
            in2 => \N__39627\,
            in3 => \N__42318\,
            lcout => \delay_measurement_inst.N_312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39624\,
            in1 => \N__39618\,
            in2 => \N__39612\,
            in3 => \N__39603\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39591\,
            in1 => \N__39585\,
            in2 => \N__39579\,
            in3 => \N__39570\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0_19_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39558\,
            in2 => \_gnd_net_\,
            in3 => \N__39440\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI21LR_6_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39531\,
            in2 => \_gnd_net_\,
            in3 => \N__42335\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_26_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__39479\,
            in1 => \N__46380\,
            in2 => \_gnd_net_\,
            in3 => \N__46222\,
            lcout => measured_delay_hc_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45936\,
            ce => 'H',
            sr => \N__45560\
        );

    \delay_measurement_inst.delay_hc_reg_17_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011101110"
        )
    port map (
            in0 => \N__39465\,
            in1 => \N__46378\,
            in2 => \N__46641\,
            in3 => \N__46220\,
            lcout => measured_delay_hc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45936\,
            ce => 'H',
            sr => \N__45560\
        );

    \delay_measurement_inst.delay_hc_reg_20_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__39441\,
            in1 => \N__46379\,
            in2 => \_gnd_net_\,
            in3 => \N__46221\,
            lcout => measured_delay_hc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45936\,
            ce => 'H',
            sr => \N__45560\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40838\,
            in2 => \_gnd_net_\,
            in3 => \N__39856\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_461_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC1_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39813\,
            lcout => delay_hc_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC2_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39804\,
            lcout => delay_hc_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40461\,
            in1 => \N__43870\,
            in2 => \_gnd_net_\,
            in3 => \N__39798\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__46053\,
            ce => \N__40385\,
            sr => \N__45441\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40456\,
            in1 => \N__39781\,
            in2 => \_gnd_net_\,
            in3 => \N__39762\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__46053\,
            ce => \N__40385\,
            sr => \N__45441\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40462\,
            in1 => \N__39751\,
            in2 => \_gnd_net_\,
            in3 => \N__39735\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__46053\,
            ce => \N__40385\,
            sr => \N__45441\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40457\,
            in1 => \N__39730\,
            in2 => \_gnd_net_\,
            in3 => \N__39714\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__46053\,
            ce => \N__40385\,
            sr => \N__45441\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40463\,
            in1 => \N__39703\,
            in2 => \_gnd_net_\,
            in3 => \N__39684\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__46053\,
            ce => \N__40385\,
            sr => \N__45441\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40458\,
            in1 => \N__39673\,
            in2 => \_gnd_net_\,
            in3 => \N__39654\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__46053\,
            ce => \N__40385\,
            sr => \N__45441\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40460\,
            in1 => \N__40078\,
            in2 => \_gnd_net_\,
            in3 => \N__40062\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__46053\,
            ce => \N__40385\,
            sr => \N__45441\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40459\,
            in1 => \N__40046\,
            in2 => \_gnd_net_\,
            in3 => \N__40032\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__46053\,
            ce => \N__40385\,
            sr => \N__45441\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40525\,
            in1 => \N__40021\,
            in2 => \_gnd_net_\,
            in3 => \N__40002\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__46045\,
            ce => \N__40377\,
            sr => \N__45444\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40529\,
            in1 => \N__39995\,
            in2 => \_gnd_net_\,
            in3 => \N__39969\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__46045\,
            ce => \N__40377\,
            sr => \N__45444\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40522\,
            in1 => \N__39958\,
            in2 => \_gnd_net_\,
            in3 => \N__39942\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__46045\,
            ce => \N__40377\,
            sr => \N__45444\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40526\,
            in1 => \N__39937\,
            in2 => \_gnd_net_\,
            in3 => \N__39921\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__46045\,
            ce => \N__40377\,
            sr => \N__45444\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40523\,
            in1 => \N__39911\,
            in2 => \_gnd_net_\,
            in3 => \N__39897\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__46045\,
            ce => \N__40377\,
            sr => \N__45444\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40527\,
            in1 => \N__39886\,
            in2 => \_gnd_net_\,
            in3 => \N__39867\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__46045\,
            ce => \N__40377\,
            sr => \N__45444\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40524\,
            in1 => \N__40313\,
            in2 => \_gnd_net_\,
            in3 => \N__40299\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__46045\,
            ce => \N__40377\,
            sr => \N__45444\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40528\,
            in1 => \N__40288\,
            in2 => \_gnd_net_\,
            in3 => \N__40272\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__46045\,
            ce => \N__40377\,
            sr => \N__45444\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40530\,
            in1 => \N__40258\,
            in2 => \_gnd_net_\,
            in3 => \N__40239\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__46037\,
            ce => \N__40386\,
            sr => \N__45447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40485\,
            in1 => \N__40231\,
            in2 => \_gnd_net_\,
            in3 => \N__40212\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__46037\,
            ce => \N__40386\,
            sr => \N__45447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40531\,
            in1 => \N__40201\,
            in2 => \_gnd_net_\,
            in3 => \N__40185\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__46037\,
            ce => \N__40386\,
            sr => \N__45447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40486\,
            in1 => \N__40169\,
            in2 => \_gnd_net_\,
            in3 => \N__40155\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__46037\,
            ce => \N__40386\,
            sr => \N__45447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40532\,
            in1 => \N__40144\,
            in2 => \_gnd_net_\,
            in3 => \N__40125\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__46037\,
            ce => \N__40386\,
            sr => \N__45447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40487\,
            in1 => \N__40120\,
            in2 => \_gnd_net_\,
            in3 => \N__40104\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__46037\,
            ce => \N__40386\,
            sr => \N__45447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40533\,
            in1 => \N__40099\,
            in2 => \_gnd_net_\,
            in3 => \N__40083\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__46037\,
            ce => \N__40386\,
            sr => \N__45447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40488\,
            in1 => \N__40684\,
            in2 => \_gnd_net_\,
            in3 => \N__40668\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__46037\,
            ce => \N__40386\,
            sr => \N__45447\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40489\,
            in1 => \N__40657\,
            in2 => \_gnd_net_\,
            in3 => \N__40638\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__46026\,
            ce => \N__40378\,
            sr => \N__45455\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40493\,
            in1 => \N__40627\,
            in2 => \_gnd_net_\,
            in3 => \N__40605\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__46026\,
            ce => \N__40378\,
            sr => \N__45455\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40490\,
            in1 => \N__40594\,
            in2 => \_gnd_net_\,
            in3 => \N__40578\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__46026\,
            ce => \N__40378\,
            sr => \N__45455\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40494\,
            in1 => \N__40573\,
            in2 => \_gnd_net_\,
            in3 => \N__40557\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__46026\,
            ce => \N__40378\,
            sr => \N__45455\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40491\,
            in1 => \N__40550\,
            in2 => \_gnd_net_\,
            in3 => \N__40536\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__46026\,
            ce => \N__40378\,
            sr => \N__45455\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__40400\,
            in1 => \N__40492\,
            in2 => \_gnd_net_\,
            in3 => \N__40410\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46026\,
            ce => \N__40378\,
            sr => \N__45455\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40347\,
            in2 => \_gnd_net_\,
            in3 => \N__40341\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__43286\,
            in1 => \N__42996\,
            in2 => \_gnd_net_\,
            in3 => \N__43401\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__40715\,
            in1 => \N__40866\,
            in2 => \N__45624\,
            in3 => \N__40749\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__44584\,
            in1 => \N__44429\,
            in2 => \_gnd_net_\,
            in3 => \N__44300\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__40782\,
            in1 => \N__43944\,
            in2 => \N__40797\,
            in3 => \N__47070\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46000\,
            ce => 'H',
            sr => \N__45469\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44428\,
            in2 => \_gnd_net_\,
            in3 => \N__44299\,
            lcout => \phase_controller_inst2.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__44301\,
            in1 => \N__44585\,
            in2 => \N__44474\,
            in3 => \N__43998\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46000\,
            ce => 'H',
            sr => \N__45469\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__44476\,
            in1 => \N__44338\,
            in2 => \N__44641\,
            in3 => \N__43962\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45991\,
            ce => 'H',
            sr => \N__45478\
        );

    \delay_measurement_inst.prev_hc_sig_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40761\,
            lcout => \delay_measurement_inst.prev_hc_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45991\,
            ce => 'H',
            sr => \N__45478\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__44477\,
            in1 => \N__44019\,
            in2 => \N__44642\,
            in3 => \N__44339\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45991\,
            ce => 'H',
            sr => \N__45478\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__44475\,
            in1 => \N__44337\,
            in2 => \N__44640\,
            in3 => \N__43971\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45991\,
            ce => 'H',
            sr => \N__45478\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010000010"
        )
    port map (
            in0 => \N__43896\,
            in1 => \N__44482\,
            in2 => \N__44663\,
            in3 => \N__44345\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45981\,
            ce => 'H',
            sr => \N__45484\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100010001100"
        )
    port map (
            in0 => \N__44342\,
            in1 => \N__44085\,
            in2 => \N__44507\,
            in3 => \N__44639\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45981\,
            ce => 'H',
            sr => \N__45484\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__44341\,
            in1 => \N__44632\,
            in2 => \N__44506\,
            in3 => \N__44094\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45981\,
            ce => 'H',
            sr => \N__45484\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010000010"
        )
    port map (
            in0 => \N__43986\,
            in1 => \N__44481\,
            in2 => \N__44662\,
            in3 => \N__44344\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45981\,
            ce => 'H',
            sr => \N__45484\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__44631\,
            in1 => \N__44343\,
            in2 => \N__44505\,
            in3 => \N__44073\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45981\,
            ce => 'H',
            sr => \N__45484\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__41294\,
            in1 => \N__41464\,
            in2 => \N__46755\,
            in3 => \N__46939\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45975\,
            ce => \N__46561\,
            sr => \N__45489\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__46937\,
            in1 => \N__41778\,
            in2 => \N__41497\,
            in3 => \N__40950\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45975\,
            ce => \N__46561\,
            sr => \N__45489\
        );

    \phase_controller_inst2.stoper_hc.target_time_0_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__42077\,
            in1 => \N__41463\,
            in2 => \N__41780\,
            in3 => \N__46938\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45975\,
            ce => \N__46561\,
            sr => \N__45489\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__46935\,
            in1 => \N__41936\,
            in2 => \N__41495\,
            in3 => \N__40898\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45975\,
            ce => \N__46561\,
            sr => \N__45489\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__41240\,
            in1 => \N__41465\,
            in2 => \N__41781\,
            in3 => \N__46940\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45975\,
            ce => \N__46561\,
            sr => \N__45489\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__46936\,
            in1 => \N__41771\,
            in2 => \N__41496\,
            in3 => \N__41196\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45975\,
            ce => \N__46561\,
            sr => \N__45489\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_18_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011111100"
        )
    port map (
            in0 => \N__41375\,
            in1 => \N__41151\,
            in2 => \N__41142\,
            in3 => \N__41133\,
            lcout => \phase_controller_inst1.stoper_hc.N_405\,
            ltout => \phase_controller_inst1.stoper_hc.N_405_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__46890\,
            in1 => \N__41764\,
            in2 => \N__41127\,
            in3 => \N__46128\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45971\,
            ce => \N__46579\,
            sr => \N__45493\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__41124\,
            in1 => \N__41462\,
            in2 => \N__41779\,
            in3 => \N__46892\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45971\,
            ce => \N__46579\,
            sr => \N__45493\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__41763\,
            in1 => \N__41461\,
            in2 => \N__41079\,
            in3 => \N__46891\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45971\,
            ce => \N__46579\,
            sr => \N__45493\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__41733\,
            in1 => \N__41475\,
            in2 => \N__41030\,
            in3 => \N__46835\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45966\,
            ce => \N__46577\,
            sr => \N__45500\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__46833\,
            in1 => \N__42260\,
            in2 => \N__41499\,
            in3 => \N__41736\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45966\,
            ce => \N__46577\,
            sr => \N__45500\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__41734\,
            in1 => \N__41476\,
            in2 => \N__40992\,
            in3 => \N__46836\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45966\,
            ce => \N__46577\,
            sr => \N__45500\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__46832\,
            in1 => \N__41829\,
            in2 => \N__41498\,
            in3 => \N__41735\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45966\,
            ce => \N__46577\,
            sr => \N__45500\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0_3_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__41670\,
            in1 => \N__46729\,
            in2 => \N__42006\,
            in3 => \N__46831\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__46834\,
            in1 => \N__41645\,
            in2 => \N__41598\,
            in3 => \N__41494\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45966\,
            ce => \N__46577\,
            sr => \N__45500\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__46844\,
            in1 => \N__46717\,
            in2 => \N__41594\,
            in3 => \N__41493\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45960\,
            ce => \N__46581\,
            sr => \N__45509\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__41492\,
            in1 => \N__41374\,
            in2 => \N__46734\,
            in3 => \N__46846\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45960\,
            ce => \N__46581\,
            sr => \N__45509\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6_19_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41252\,
            in1 => \N__42089\,
            in2 => \N__41328\,
            in3 => \N__42101\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__46716\,
            in1 => \N__41866\,
            in2 => \_gnd_net_\,
            in3 => \N__46845\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45960\,
            ce => \N__46581\,
            sr => \N__45509\
        );

    \delay_measurement_inst.delay_hc_reg_6_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011111011"
        )
    port map (
            in0 => \N__46460\,
            in1 => \N__46253\,
            in2 => \N__41292\,
            in3 => \N__42294\,
            lcout => measured_delay_hc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45955\,
            ce => 'H',
            sr => \N__45516\
        );

    \delay_measurement_inst.delay_hc_reg_29_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__46251\,
            in1 => \_gnd_net_\,
            in2 => \N__46493\,
            in3 => \N__41253\,
            lcout => measured_delay_hc_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45955\,
            ce => 'H',
            sr => \N__45516\
        );

    \delay_measurement_inst.delay_hc_reg_27_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__42102\,
            in1 => \N__46452\,
            in2 => \_gnd_net_\,
            in3 => \N__46249\,
            lcout => measured_delay_hc_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45955\,
            ce => 'H',
            sr => \N__45516\
        );

    \delay_measurement_inst.delay_hc_reg_28_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__46250\,
            in1 => \_gnd_net_\,
            in2 => \N__46492\,
            in3 => \N__42090\,
            lcout => measured_delay_hc_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45955\,
            ce => 'H',
            sr => \N__45516\
        );

    \delay_measurement_inst.delay_hc_reg_31_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__46713\,
            in1 => \N__46459\,
            in2 => \_gnd_net_\,
            in3 => \N__46252\,
            lcout => measured_delay_hc_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45955\,
            ce => 'H',
            sr => \N__45516\
        );

    \delay_measurement_inst.delay_hc_reg_0_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__42066\,
            in1 => \N__46451\,
            in2 => \_gnd_net_\,
            in3 => \N__46248\,
            lcout => measured_delay_hc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45955\,
            ce => 'H',
            sr => \N__45516\
        );

    \delay_measurement_inst.delay_hc_reg_19_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__46176\,
            in1 => \N__42045\,
            in2 => \N__46449\,
            in3 => \N__41997\,
            lcout => measured_delay_hc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45952\,
            ce => 'H',
            sr => \N__45525\
        );

    \delay_measurement_inst.delay_hc_reg_16_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011101110"
        )
    port map (
            in0 => \N__41961\,
            in1 => \N__46387\,
            in2 => \N__46994\,
            in3 => \N__46174\,
            lcout => measured_delay_hc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45952\,
            ce => 'H',
            sr => \N__45525\
        );

    \delay_measurement_inst.delay_hc_reg_1_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__46177\,
            in1 => \N__42423\,
            in2 => \N__46450\,
            in3 => \N__41921\,
            lcout => measured_delay_hc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45952\,
            ce => 'H',
            sr => \N__45525\
        );

    \delay_measurement_inst.delay_hc_reg_18_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__41858\,
            in1 => \N__46388\,
            in2 => \N__41895\,
            in3 => \N__46175\,
            lcout => measured_delay_hc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45952\,
            ce => 'H',
            sr => \N__45525\
        );

    \reset_ibuf_gb_io_RNI79U7_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45619\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => red_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42422\,
            in1 => \N__46304\,
            in2 => \N__42405\,
            in3 => \N__42371\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_6_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__42339\,
            in1 => \N__42317\,
            in2 => \_gnd_net_\,
            in3 => \N__42305\,
            lcout => \delay_measurement_inst.N_295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_15_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__42285\,
            in1 => \N__46352\,
            in2 => \N__42256\,
            in3 => \N__46254\,
            lcout => measured_delay_hc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45944\,
            ce => 'H',
            sr => \N__45547\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42617\,
            in1 => \N__42938\,
            in2 => \N__42213\,
            in3 => \N__42814\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45442\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42813\,
            in1 => \N__42619\,
            in2 => \N__42959\,
            in3 => \N__42168\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45442\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42618\,
            in1 => \N__42939\,
            in2 => \N__42132\,
            in3 => \N__42815\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45442\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__43953\,
            in1 => \N__44221\,
            in2 => \_gnd_net_\,
            in3 => \N__47069\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__44473\,
            in1 => \N__44666\,
            in2 => \N__42105\,
            in3 => \N__44357\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45442\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__44472\,
            in1 => \N__44667\,
            in2 => \N__44358\,
            in3 => \N__44010\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46054\,
            ce => 'H',
            sr => \N__45442\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43880\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46046\,
            ce => \N__43828\,
            sr => \N__45445\
        );

    \delay_measurement_inst.delay_tr_reg_esr_17_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__43672\,
            in1 => \N__43805\,
            in2 => \_gnd_net_\,
            in3 => \N__43730\,
            lcout => measured_delay_tr_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46038\,
            ce => \N__43515\,
            sr => \N__45448\
        );

    \delay_measurement_inst.delay_tr_reg_esr_18_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__43731\,
            in1 => \N__43673\,
            in2 => \_gnd_net_\,
            in3 => \N__43581\,
            lcout => measured_delay_tr_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46038\,
            ce => \N__43515\,
            sr => \N__45448\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001001010"
        )
    port map (
            in0 => \N__43450\,
            in1 => \N__43330\,
            in2 => \N__43031\,
            in3 => \N__43176\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46027\,
            ce => \N__42510\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100001011000"
        )
    port map (
            in0 => \N__42540\,
            in1 => \N__42943\,
            in2 => \N__42819\,
            in3 => \N__42680\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46027\,
            ce => \N__42510\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_0_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__44444\,
            in1 => \N__44653\,
            in2 => \N__44340\,
            in3 => \N__47061\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46027\,
            ce => \N__42510\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_1_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111000000"
        )
    port map (
            in0 => \N__47062\,
            in1 => \N__44445\,
            in2 => \N__44665\,
            in3 => \N__44298\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__46027\,
            ce => \N__42510\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43945\,
            in2 => \_gnd_net_\,
            in3 => \N__47059\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__47060\,
            in1 => \_gnd_net_\,
            in2 => \N__43952\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43923\,
            in2 => \N__44229\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44184\,
            in2 => \_gnd_net_\,
            in3 => \N__43917\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43914\,
            in2 => \N__44163\,
            in3 => \N__43908\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44115\,
            in2 => \_gnd_net_\,
            in3 => \N__43905\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44904\,
            in2 => \_gnd_net_\,
            in3 => \N__43902\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44883\,
            in2 => \_gnd_net_\,
            in3 => \N__43899\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44853\,
            in2 => \_gnd_net_\,
            in3 => \N__43887\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44814\,
            in2 => \_gnd_net_\,
            in3 => \N__43884\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44774\,
            in2 => \_gnd_net_\,
            in3 => \N__44013\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44744\,
            in2 => \_gnd_net_\,
            in3 => \N__44001\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44708\,
            in2 => \_gnd_net_\,
            in3 => \N__43992\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45150\,
            in2 => \_gnd_net_\,
            in3 => \N__43989\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45126\,
            in2 => \_gnd_net_\,
            in3 => \N__43977\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45077\,
            in2 => \_gnd_net_\,
            in3 => \N__43974\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45032\,
            in2 => \_gnd_net_\,
            in3 => \N__43965\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45008\,
            in2 => \_gnd_net_\,
            in3 => \N__43956\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44987\,
            in2 => \_gnd_net_\,
            in3 => \N__44088\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44957\,
            in2 => \_gnd_net_\,
            in3 => \N__44079\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44936\,
            in2 => \_gnd_net_\,
            in3 => \N__44076\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__44560\,
            in1 => \N__44433\,
            in2 => \_gnd_net_\,
            in3 => \N__44302\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__44346\,
            in1 => \N__44646\,
            in2 => \N__44508\,
            in3 => \N__44067\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45992\,
            ce => 'H',
            sr => \N__45479\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__44645\,
            in1 => \N__44492\,
            in2 => \N__44058\,
            in3 => \N__44352\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45992\,
            ce => 'H',
            sr => \N__45479\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__44348\,
            in1 => \N__44648\,
            in2 => \N__44510\,
            in3 => \N__44046\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45992\,
            ce => 'H',
            sr => \N__45479\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010000010"
        )
    port map (
            in0 => \N__44037\,
            in1 => \N__44489\,
            in2 => \N__44664\,
            in3 => \N__44353\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45992\,
            ce => 'H',
            sr => \N__45479\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__44347\,
            in1 => \N__44647\,
            in2 => \N__44509\,
            in3 => \N__44028\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45992\,
            ce => 'H',
            sr => \N__45479\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__44643\,
            in1 => \N__44490\,
            in2 => \N__44688\,
            in3 => \N__44350\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45992\,
            ce => 'H',
            sr => \N__45479\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__44349\,
            in1 => \N__44649\,
            in2 => \N__44511\,
            in3 => \N__44676\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45992\,
            ce => 'H',
            sr => \N__45479\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__44644\,
            in1 => \N__44491\,
            in2 => \N__44373\,
            in3 => \N__44351\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45992\,
            ce => 'H',
            sr => \N__45479\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44247\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44202\,
            in2 => \N__44238\,
            in3 => \N__44228\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44169\,
            in2 => \N__44196\,
            in3 => \N__44180\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44156\,
            in1 => \N__44130\,
            in2 => \N__44145\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44100\,
            in2 => \N__44124\,
            in3 => \N__44111\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44889\,
            in2 => \N__44916\,
            in3 => \N__44900\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44879\,
            in1 => \N__44859\,
            in2 => \N__44868\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44849\,
            in1 => \N__44826\,
            in2 => \N__44838\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44820\,
            in2 => \N__44796\,
            in3 => \N__44813\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44760\,
            in2 => \N__44787\,
            in3 => \N__44775\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44727\,
            in2 => \N__44754\,
            in3 => \N__44745\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44694\,
            in2 => \N__44721\,
            in3 => \N__44712\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45132\,
            in2 => \N__45159\,
            in3 => \N__45149\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45122\,
            in1 => \N__45096\,
            in2 => \N__45108\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45090\,
            in2 => \N__45057\,
            in3 => \N__45078\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45018\,
            in2 => \N__45048\,
            in3 => \N__45036\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44994\,
            in2 => \N__46956\,
            in3 => \N__45012\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44973\,
            in2 => \N__46593\,
            in3 => \N__44988\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44943\,
            in2 => \N__44967\,
            in3 => \N__44958\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44922\,
            in2 => \N__47004\,
            in3 => \N__44937\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47073\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46712\,
            in2 => \_gnd_net_\,
            in3 => \N__47028\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45967\,
            ce => \N__46580\,
            sr => \N__45501\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__46714\,
            in1 => \N__46984\,
            in2 => \_gnd_net_\,
            in3 => \N__46917\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45961\,
            ce => \N__46578\,
            sr => \N__45510\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__46916\,
            in1 => \N__46715\,
            in2 => \_gnd_net_\,
            in3 => \N__46647\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45961\,
            ce => \N__46578\,
            sr => \N__45510\
        );

    \delay_measurement_inst.delay_hc_reg_25_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__46514\,
            in1 => \N__46482\,
            in2 => \_gnd_net_\,
            in3 => \N__46276\,
            lcout => measured_delay_hc_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45956\,
            ce => 'H',
            sr => \N__45517\
        );

    \delay_measurement_inst.delay_hc_reg_2_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__46112\,
            in1 => \N__46483\,
            in2 => \N__46311\,
            in3 => \N__46277\,
            lcout => measured_delay_hc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45956\,
            ce => 'H',
            sr => \N__45517\
        );
end \INTERFACE\;
